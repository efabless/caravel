magic
tech sky130A
magscale 1 2
timestamp 1665682149
<< viali >>
rect 1869 3553 1903 3587
rect 6745 3485 6779 3519
rect 1133 3417 1167 3451
rect 6009 3417 6043 3451
rect 1869 3077 1903 3111
rect 3249 3077 3283 3111
rect 5825 3077 5859 3111
rect 2605 2941 2639 2975
rect 3985 2941 4019 2975
rect 6561 2941 6595 2975
rect 2697 2397 2731 2431
rect 4169 2397 4203 2431
rect 5549 2397 5583 2431
rect 1961 2329 1995 2363
rect 4905 2329 4939 2363
rect 6285 2329 6319 2363
rect 1133 1989 1167 2023
rect 3249 1989 3283 2023
rect 3709 1989 3743 2023
rect 5825 1989 5859 2023
rect 1869 1921 1903 1955
rect 2513 1853 2547 1887
rect 4445 1853 4479 1887
rect 6561 1853 6595 1887
rect 1869 1309 1903 1343
rect 5273 1309 5307 1343
rect 6745 1309 6779 1343
rect 1133 1241 1167 1275
rect 4537 1241 4571 1275
rect 6009 1241 6043 1275
<< metal1 >>
rect 368 3834 7544 3856
rect 368 3782 1110 3834
rect 1162 3782 1174 3834
rect 1226 3782 1238 3834
rect 1290 3782 1302 3834
rect 1354 3782 1366 3834
rect 1418 3782 2903 3834
rect 2955 3782 2967 3834
rect 3019 3782 3031 3834
rect 3083 3782 3095 3834
rect 3147 3782 3159 3834
rect 3211 3782 4696 3834
rect 4748 3782 4760 3834
rect 4812 3782 4824 3834
rect 4876 3782 4888 3834
rect 4940 3782 4952 3834
rect 5004 3782 6489 3834
rect 6541 3782 6553 3834
rect 6605 3782 6617 3834
rect 6669 3782 6681 3834
rect 6733 3782 6745 3834
rect 6797 3782 7544 3834
rect 368 3760 7544 3782
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1544 3556 1869 3584
rect 1544 3544 1550 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3516 6791 3519
rect 6822 3516 6828 3528
rect 6779 3488 6828 3516
rect 6779 3485 6791 3488
rect 6733 3479 6791 3485
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 1121 3451 1179 3457
rect 1121 3448 1133 3451
rect 1084 3420 1133 3448
rect 1084 3408 1090 3420
rect 1121 3417 1133 3420
rect 1167 3417 1179 3451
rect 1121 3411 1179 3417
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3448 6055 3451
rect 6043 3420 6868 3448
rect 6043 3417 6055 3420
rect 5997 3411 6055 3417
rect 6840 3392 6868 3420
rect 6822 3340 6828 3392
rect 6880 3340 6886 3392
rect 368 3290 7699 3312
rect 368 3238 2006 3290
rect 2058 3238 2070 3290
rect 2122 3238 2134 3290
rect 2186 3238 2198 3290
rect 2250 3238 2262 3290
rect 2314 3238 3799 3290
rect 3851 3238 3863 3290
rect 3915 3238 3927 3290
rect 3979 3238 3991 3290
rect 4043 3238 4055 3290
rect 4107 3238 5592 3290
rect 5644 3238 5656 3290
rect 5708 3238 5720 3290
rect 5772 3238 5784 3290
rect 5836 3238 5848 3290
rect 5900 3238 7385 3290
rect 7437 3238 7449 3290
rect 7501 3238 7513 3290
rect 7565 3238 7577 3290
rect 7629 3238 7641 3290
rect 7693 3238 7699 3290
rect 368 3216 7699 3238
rect 1854 3108 1860 3120
rect 1815 3080 1860 3108
rect 1854 3068 1860 3080
rect 1912 3068 1918 3120
rect 3234 3108 3240 3120
rect 3195 3080 3240 3108
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 5994 3108 6000 3120
rect 5859 3080 6000 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 2406 2932 2412 2984
rect 2464 2972 2470 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2464 2944 2605 2972
rect 2464 2932 2470 2944
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 2593 2935 2651 2941
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3568 2944 3985 2972
rect 3568 2932 3574 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6052 2944 6561 2972
rect 6052 2932 6058 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 368 2746 7544 2768
rect 368 2694 1110 2746
rect 1162 2694 1174 2746
rect 1226 2694 1238 2746
rect 1290 2694 1302 2746
rect 1354 2694 1366 2746
rect 1418 2694 2903 2746
rect 2955 2694 2967 2746
rect 3019 2694 3031 2746
rect 3083 2694 3095 2746
rect 3147 2694 3159 2746
rect 3211 2694 4696 2746
rect 4748 2694 4760 2746
rect 4812 2694 4824 2746
rect 4876 2694 4888 2746
rect 4940 2694 4952 2746
rect 5004 2694 6489 2746
rect 6541 2694 6553 2746
rect 6605 2694 6617 2746
rect 6669 2694 6681 2746
rect 6733 2694 6745 2746
rect 6797 2694 7544 2746
rect 368 2672 7544 2694
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 4154 2428 4160 2440
rect 4115 2400 4160 2428
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5316 2400 5549 2428
rect 5316 2388 5322 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 2590 2360 2596 2372
rect 1995 2332 2596 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2590 2320 2596 2332
rect 2648 2320 2654 2372
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 4893 2363 4951 2369
rect 4893 2360 4905 2363
rect 4488 2332 4905 2360
rect 4488 2320 4494 2332
rect 4893 2329 4905 2332
rect 4939 2329 4951 2363
rect 4893 2323 4951 2329
rect 5074 2320 5080 2372
rect 5132 2360 5138 2372
rect 6273 2363 6331 2369
rect 6273 2360 6285 2363
rect 5132 2332 6285 2360
rect 5132 2320 5138 2332
rect 6273 2329 6285 2332
rect 6319 2329 6331 2363
rect 6273 2323 6331 2329
rect 368 2202 7699 2224
rect 368 2150 2006 2202
rect 2058 2150 2070 2202
rect 2122 2150 2134 2202
rect 2186 2150 2198 2202
rect 2250 2150 2262 2202
rect 2314 2150 3799 2202
rect 3851 2150 3863 2202
rect 3915 2150 3927 2202
rect 3979 2150 3991 2202
rect 4043 2150 4055 2202
rect 4107 2150 5592 2202
rect 5644 2150 5656 2202
rect 5708 2150 5720 2202
rect 5772 2150 5784 2202
rect 5836 2150 5848 2202
rect 5900 2150 7385 2202
rect 7437 2150 7449 2202
rect 7501 2150 7513 2202
rect 7565 2150 7577 2202
rect 7629 2150 7641 2202
rect 7693 2150 7699 2202
rect 368 2128 7699 2150
rect 1121 2023 1179 2029
rect 1121 1989 1133 2023
rect 1167 2020 1179 2023
rect 1578 2020 1584 2032
rect 1167 1992 1584 2020
rect 1167 1989 1179 1992
rect 1121 1983 1179 1989
rect 1578 1980 1584 1992
rect 1636 1980 1642 2032
rect 2774 1980 2780 2032
rect 2832 2020 2838 2032
rect 3237 2023 3295 2029
rect 3237 2020 3249 2023
rect 2832 1992 3249 2020
rect 2832 1980 2838 1992
rect 3237 1989 3249 1992
rect 3283 1989 3295 2023
rect 3694 2020 3700 2032
rect 3655 1992 3700 2020
rect 3237 1983 3295 1989
rect 3694 1980 3700 1992
rect 3752 1980 3758 2032
rect 5350 1980 5356 2032
rect 5408 2020 5414 2032
rect 5813 2023 5871 2029
rect 5813 2020 5825 2023
rect 5408 1992 5825 2020
rect 5408 1980 5414 1992
rect 5813 1989 5825 1992
rect 5859 1989 5871 2023
rect 5813 1983 5871 1989
rect 1670 1912 1676 1964
rect 1728 1952 1734 1964
rect 1857 1955 1915 1961
rect 1857 1952 1869 1955
rect 1728 1924 1869 1952
rect 1728 1912 1734 1924
rect 1857 1921 1869 1924
rect 1903 1921 1915 1955
rect 1857 1915 1915 1921
rect 2501 1887 2559 1893
rect 2501 1853 2513 1887
rect 2547 1884 2559 1887
rect 2774 1884 2780 1896
rect 2547 1856 2780 1884
rect 2547 1853 2559 1856
rect 2501 1847 2559 1853
rect 2774 1844 2780 1856
rect 2832 1844 2838 1896
rect 4154 1844 4160 1896
rect 4212 1884 4218 1896
rect 4433 1887 4491 1893
rect 4433 1884 4445 1887
rect 4212 1856 4445 1884
rect 4212 1844 4218 1856
rect 4433 1853 4445 1856
rect 4479 1853 4491 1887
rect 4433 1847 4491 1853
rect 5350 1844 5356 1896
rect 5408 1884 5414 1896
rect 6549 1887 6607 1893
rect 6549 1884 6561 1887
rect 5408 1856 6561 1884
rect 5408 1844 5414 1856
rect 6549 1853 6561 1856
rect 6595 1853 6607 1887
rect 6549 1847 6607 1853
rect 368 1658 7544 1680
rect 368 1606 1110 1658
rect 1162 1606 1174 1658
rect 1226 1606 1238 1658
rect 1290 1606 1302 1658
rect 1354 1606 1366 1658
rect 1418 1606 2903 1658
rect 2955 1606 2967 1658
rect 3019 1606 3031 1658
rect 3083 1606 3095 1658
rect 3147 1606 3159 1658
rect 3211 1606 4696 1658
rect 4748 1606 4760 1658
rect 4812 1606 4824 1658
rect 4876 1606 4888 1658
rect 4940 1606 4952 1658
rect 5004 1606 6489 1658
rect 6541 1606 6553 1658
rect 6605 1606 6617 1658
rect 6669 1606 6681 1658
rect 6733 1606 6745 1658
rect 6797 1606 7544 1658
rect 368 1584 7544 1606
rect 6288 1380 6868 1408
rect 934 1300 940 1352
rect 992 1340 998 1352
rect 1857 1343 1915 1349
rect 1857 1340 1869 1343
rect 992 1312 1869 1340
rect 992 1300 998 1312
rect 1857 1309 1869 1312
rect 1903 1309 1915 1343
rect 1857 1303 1915 1309
rect 5261 1343 5319 1349
rect 5261 1309 5273 1343
rect 5307 1340 5319 1343
rect 6288 1340 6316 1380
rect 5307 1312 6316 1340
rect 5307 1309 5319 1312
rect 5261 1303 5319 1309
rect 6362 1300 6368 1352
rect 6420 1340 6426 1352
rect 6733 1343 6791 1349
rect 6733 1340 6745 1343
rect 6420 1312 6745 1340
rect 6420 1300 6426 1312
rect 6733 1309 6745 1312
rect 6779 1309 6791 1343
rect 6840 1340 6868 1380
rect 7190 1340 7196 1352
rect 6840 1312 7196 1340
rect 6733 1303 6791 1309
rect 7190 1300 7196 1312
rect 7248 1300 7254 1352
rect 750 1232 756 1284
rect 808 1272 814 1284
rect 1121 1275 1179 1281
rect 1121 1272 1133 1275
rect 808 1244 1133 1272
rect 808 1232 814 1244
rect 1121 1241 1133 1244
rect 1167 1241 1179 1275
rect 1121 1235 1179 1241
rect 4525 1275 4583 1281
rect 4525 1241 4537 1275
rect 4571 1241 4583 1275
rect 4525 1235 4583 1241
rect 5997 1275 6055 1281
rect 5997 1241 6009 1275
rect 6043 1272 6055 1275
rect 6270 1272 6276 1284
rect 6043 1244 6276 1272
rect 6043 1241 6055 1244
rect 5997 1235 6055 1241
rect 4540 1204 4568 1235
rect 6270 1232 6276 1244
rect 6328 1232 6334 1284
rect 7190 1204 7196 1216
rect 4540 1176 7196 1204
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
rect 368 1114 7699 1136
rect 368 1062 2006 1114
rect 2058 1062 2070 1114
rect 2122 1062 2134 1114
rect 2186 1062 2198 1114
rect 2250 1062 2262 1114
rect 2314 1062 3799 1114
rect 3851 1062 3863 1114
rect 3915 1062 3927 1114
rect 3979 1062 3991 1114
rect 4043 1062 4055 1114
rect 4107 1062 5592 1114
rect 5644 1062 5656 1114
rect 5708 1062 5720 1114
rect 5772 1062 5784 1114
rect 5836 1062 5848 1114
rect 5900 1062 7385 1114
rect 7437 1062 7449 1114
rect 7501 1062 7513 1114
rect 7565 1062 7577 1114
rect 7629 1062 7641 1114
rect 7693 1062 7699 1114
rect 368 1040 7699 1062
<< via1 >>
rect 1110 3782 1162 3834
rect 1174 3782 1226 3834
rect 1238 3782 1290 3834
rect 1302 3782 1354 3834
rect 1366 3782 1418 3834
rect 2903 3782 2955 3834
rect 2967 3782 3019 3834
rect 3031 3782 3083 3834
rect 3095 3782 3147 3834
rect 3159 3782 3211 3834
rect 4696 3782 4748 3834
rect 4760 3782 4812 3834
rect 4824 3782 4876 3834
rect 4888 3782 4940 3834
rect 4952 3782 5004 3834
rect 6489 3782 6541 3834
rect 6553 3782 6605 3834
rect 6617 3782 6669 3834
rect 6681 3782 6733 3834
rect 6745 3782 6797 3834
rect 1492 3544 1544 3596
rect 6828 3476 6880 3528
rect 1032 3408 1084 3460
rect 6828 3340 6880 3392
rect 2006 3238 2058 3290
rect 2070 3238 2122 3290
rect 2134 3238 2186 3290
rect 2198 3238 2250 3290
rect 2262 3238 2314 3290
rect 3799 3238 3851 3290
rect 3863 3238 3915 3290
rect 3927 3238 3979 3290
rect 3991 3238 4043 3290
rect 4055 3238 4107 3290
rect 5592 3238 5644 3290
rect 5656 3238 5708 3290
rect 5720 3238 5772 3290
rect 5784 3238 5836 3290
rect 5848 3238 5900 3290
rect 7385 3238 7437 3290
rect 7449 3238 7501 3290
rect 7513 3238 7565 3290
rect 7577 3238 7629 3290
rect 7641 3238 7693 3290
rect 1860 3111 1912 3120
rect 1860 3077 1869 3111
rect 1869 3077 1903 3111
rect 1903 3077 1912 3111
rect 1860 3068 1912 3077
rect 3240 3111 3292 3120
rect 3240 3077 3249 3111
rect 3249 3077 3283 3111
rect 3283 3077 3292 3111
rect 3240 3068 3292 3077
rect 6000 3068 6052 3120
rect 2412 2932 2464 2984
rect 3516 2932 3568 2984
rect 6000 2932 6052 2984
rect 1110 2694 1162 2746
rect 1174 2694 1226 2746
rect 1238 2694 1290 2746
rect 1302 2694 1354 2746
rect 1366 2694 1418 2746
rect 2903 2694 2955 2746
rect 2967 2694 3019 2746
rect 3031 2694 3083 2746
rect 3095 2694 3147 2746
rect 3159 2694 3211 2746
rect 4696 2694 4748 2746
rect 4760 2694 4812 2746
rect 4824 2694 4876 2746
rect 4888 2694 4940 2746
rect 4952 2694 5004 2746
rect 6489 2694 6541 2746
rect 6553 2694 6605 2746
rect 6617 2694 6669 2746
rect 6681 2694 6733 2746
rect 6745 2694 6797 2746
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 5264 2388 5316 2440
rect 2596 2320 2648 2372
rect 4436 2320 4488 2372
rect 5080 2320 5132 2372
rect 2006 2150 2058 2202
rect 2070 2150 2122 2202
rect 2134 2150 2186 2202
rect 2198 2150 2250 2202
rect 2262 2150 2314 2202
rect 3799 2150 3851 2202
rect 3863 2150 3915 2202
rect 3927 2150 3979 2202
rect 3991 2150 4043 2202
rect 4055 2150 4107 2202
rect 5592 2150 5644 2202
rect 5656 2150 5708 2202
rect 5720 2150 5772 2202
rect 5784 2150 5836 2202
rect 5848 2150 5900 2202
rect 7385 2150 7437 2202
rect 7449 2150 7501 2202
rect 7513 2150 7565 2202
rect 7577 2150 7629 2202
rect 7641 2150 7693 2202
rect 1584 1980 1636 2032
rect 2780 1980 2832 2032
rect 3700 2023 3752 2032
rect 3700 1989 3709 2023
rect 3709 1989 3743 2023
rect 3743 1989 3752 2023
rect 3700 1980 3752 1989
rect 5356 1980 5408 2032
rect 1676 1912 1728 1964
rect 2780 1844 2832 1896
rect 4160 1844 4212 1896
rect 5356 1844 5408 1896
rect 1110 1606 1162 1658
rect 1174 1606 1226 1658
rect 1238 1606 1290 1658
rect 1302 1606 1354 1658
rect 1366 1606 1418 1658
rect 2903 1606 2955 1658
rect 2967 1606 3019 1658
rect 3031 1606 3083 1658
rect 3095 1606 3147 1658
rect 3159 1606 3211 1658
rect 4696 1606 4748 1658
rect 4760 1606 4812 1658
rect 4824 1606 4876 1658
rect 4888 1606 4940 1658
rect 4952 1606 5004 1658
rect 6489 1606 6541 1658
rect 6553 1606 6605 1658
rect 6617 1606 6669 1658
rect 6681 1606 6733 1658
rect 6745 1606 6797 1658
rect 940 1300 992 1352
rect 6368 1300 6420 1352
rect 7196 1300 7248 1352
rect 756 1232 808 1284
rect 6276 1232 6328 1284
rect 7196 1164 7248 1216
rect 2006 1062 2058 1114
rect 2070 1062 2122 1114
rect 2134 1062 2186 1114
rect 2198 1062 2250 1114
rect 2262 1062 2314 1114
rect 3799 1062 3851 1114
rect 3863 1062 3915 1114
rect 3927 1062 3979 1114
rect 3991 1062 4043 1114
rect 4055 1062 4107 1114
rect 5592 1062 5644 1114
rect 5656 1062 5708 1114
rect 5720 1062 5772 1114
rect 5784 1062 5836 1114
rect 5848 1062 5900 1114
rect 7385 1062 7437 1114
rect 7449 1062 7501 1114
rect 7513 1062 7565 1114
rect 7577 1062 7629 1114
rect 7641 1062 7693 1114
<< metal2 >>
rect 754 4298 810 5000
rect 1214 4298 1270 5000
rect 1674 4298 1730 5000
rect 2134 4298 2190 5000
rect 754 4270 980 4298
rect 754 4200 810 4270
rect 952 1358 980 4270
rect 1214 4270 1532 4298
rect 1214 4200 1270 4270
rect 1110 3836 1418 3845
rect 1110 3834 1116 3836
rect 1172 3834 1196 3836
rect 1252 3834 1276 3836
rect 1332 3834 1356 3836
rect 1412 3834 1418 3836
rect 1172 3782 1174 3834
rect 1354 3782 1356 3834
rect 1110 3780 1116 3782
rect 1172 3780 1196 3782
rect 1252 3780 1276 3782
rect 1332 3780 1356 3782
rect 1412 3780 1418 3782
rect 1110 3771 1418 3780
rect 1504 3602 1532 4270
rect 1596 4270 1730 4298
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 1044 1442 1072 3402
rect 1110 2748 1418 2757
rect 1110 2746 1116 2748
rect 1172 2746 1196 2748
rect 1252 2746 1276 2748
rect 1332 2746 1356 2748
rect 1412 2746 1418 2748
rect 1172 2694 1174 2746
rect 1354 2694 1356 2746
rect 1110 2692 1116 2694
rect 1172 2692 1196 2694
rect 1252 2692 1276 2694
rect 1332 2692 1356 2694
rect 1412 2692 1418 2694
rect 1110 2683 1418 2692
rect 1596 2038 1624 4270
rect 1674 4200 1730 4270
rect 1872 4270 2190 4298
rect 1872 3126 1900 4270
rect 2134 4200 2190 4270
rect 2594 4298 2650 5000
rect 3054 4298 3110 5000
rect 3514 4298 3570 5000
rect 3974 4298 4030 5000
rect 4434 4298 4490 5000
rect 2594 4270 2728 4298
rect 2594 4200 2650 4270
rect 2006 3292 2314 3301
rect 2006 3290 2012 3292
rect 2068 3290 2092 3292
rect 2148 3290 2172 3292
rect 2228 3290 2252 3292
rect 2308 3290 2314 3292
rect 2068 3238 2070 3290
rect 2250 3238 2252 3290
rect 2006 3236 2012 3238
rect 2068 3236 2092 3238
rect 2148 3236 2172 3238
rect 2228 3236 2252 3238
rect 2308 3236 2314 3238
rect 2006 3227 2314 3236
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2006 2204 2314 2213
rect 2006 2202 2012 2204
rect 2068 2202 2092 2204
rect 2148 2202 2172 2204
rect 2228 2202 2252 2204
rect 2308 2202 2314 2204
rect 2068 2150 2070 2202
rect 2250 2150 2252 2202
rect 2006 2148 2012 2150
rect 2068 2148 2092 2150
rect 2148 2148 2172 2150
rect 2228 2148 2252 2150
rect 2308 2148 2314 2150
rect 2006 2139 2314 2148
rect 1584 2032 1636 2038
rect 1584 1974 1636 1980
rect 1676 1964 1728 1970
rect 1676 1906 1728 1912
rect 1110 1660 1418 1669
rect 1110 1658 1116 1660
rect 1172 1658 1196 1660
rect 1252 1658 1276 1660
rect 1332 1658 1356 1660
rect 1412 1658 1418 1660
rect 1172 1606 1174 1658
rect 1354 1606 1356 1658
rect 1110 1604 1116 1606
rect 1172 1604 1196 1606
rect 1252 1604 1276 1606
rect 1332 1604 1356 1606
rect 1412 1604 1418 1606
rect 1110 1595 1418 1604
rect 1044 1414 1256 1442
rect 940 1352 992 1358
rect 940 1294 992 1300
rect 756 1284 808 1290
rect 756 1226 808 1232
rect 768 800 796 1226
rect 1228 800 1256 1414
rect 1688 800 1716 1906
rect 2006 1116 2314 1125
rect 2006 1114 2012 1116
rect 2068 1114 2092 1116
rect 2148 1114 2172 1116
rect 2228 1114 2252 1116
rect 2308 1114 2314 1116
rect 2068 1062 2070 1114
rect 2250 1062 2252 1114
rect 2006 1060 2012 1062
rect 2068 1060 2092 1062
rect 2148 1060 2172 1062
rect 2228 1060 2252 1062
rect 2308 1060 2314 1062
rect 2006 1051 2314 1060
rect 2148 870 2268 898
rect 2148 800 2176 870
rect 754 0 810 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2240 762 2268 870
rect 2424 762 2452 2926
rect 2700 2446 2728 4270
rect 2792 4270 3110 4298
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2608 800 2636 2314
rect 2792 2038 2820 4270
rect 3054 4200 3110 4270
rect 3252 4270 3570 4298
rect 2903 3836 3211 3845
rect 2903 3834 2909 3836
rect 2965 3834 2989 3836
rect 3045 3834 3069 3836
rect 3125 3834 3149 3836
rect 3205 3834 3211 3836
rect 2965 3782 2967 3834
rect 3147 3782 3149 3834
rect 2903 3780 2909 3782
rect 2965 3780 2989 3782
rect 3045 3780 3069 3782
rect 3125 3780 3149 3782
rect 3205 3780 3211 3782
rect 2903 3771 3211 3780
rect 3252 3126 3280 4270
rect 3514 4200 3570 4270
rect 3712 4270 4030 4298
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 2903 2748 3211 2757
rect 2903 2746 2909 2748
rect 2965 2746 2989 2748
rect 3045 2746 3069 2748
rect 3125 2746 3149 2748
rect 3205 2746 3211 2748
rect 2965 2694 2967 2746
rect 3147 2694 3149 2746
rect 2903 2692 2909 2694
rect 2965 2692 2989 2694
rect 3045 2692 3069 2694
rect 3125 2692 3149 2694
rect 3205 2692 3211 2694
rect 2903 2683 3211 2692
rect 2780 2032 2832 2038
rect 2780 1974 2832 1980
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2240 734 2452 762
rect 2594 0 2650 800
rect 2792 762 2820 1838
rect 2903 1660 3211 1669
rect 2903 1658 2909 1660
rect 2965 1658 2989 1660
rect 3045 1658 3069 1660
rect 3125 1658 3149 1660
rect 3205 1658 3211 1660
rect 2965 1606 2967 1658
rect 3147 1606 3149 1658
rect 2903 1604 2909 1606
rect 2965 1604 2989 1606
rect 3045 1604 3069 1606
rect 3125 1604 3149 1606
rect 3205 1604 3211 1606
rect 2903 1595 3211 1604
rect 2976 870 3096 898
rect 2976 762 3004 870
rect 3068 800 3096 870
rect 3528 800 3556 2926
rect 3712 2038 3740 4270
rect 3974 4200 4030 4270
rect 4172 4270 4490 4298
rect 3799 3292 4107 3301
rect 3799 3290 3805 3292
rect 3861 3290 3885 3292
rect 3941 3290 3965 3292
rect 4021 3290 4045 3292
rect 4101 3290 4107 3292
rect 3861 3238 3863 3290
rect 4043 3238 4045 3290
rect 3799 3236 3805 3238
rect 3861 3236 3885 3238
rect 3941 3236 3965 3238
rect 4021 3236 4045 3238
rect 4101 3236 4107 3238
rect 3799 3227 4107 3236
rect 4172 2446 4200 4270
rect 4434 4200 4490 4270
rect 4894 4298 4950 5000
rect 4894 4270 5304 4298
rect 4894 4200 4950 4270
rect 4696 3836 5004 3845
rect 4696 3834 4702 3836
rect 4758 3834 4782 3836
rect 4838 3834 4862 3836
rect 4918 3834 4942 3836
rect 4998 3834 5004 3836
rect 4758 3782 4760 3834
rect 4940 3782 4942 3834
rect 4696 3780 4702 3782
rect 4758 3780 4782 3782
rect 4838 3780 4862 3782
rect 4918 3780 4942 3782
rect 4998 3780 5004 3782
rect 4696 3771 5004 3780
rect 4696 2748 5004 2757
rect 4696 2746 4702 2748
rect 4758 2746 4782 2748
rect 4838 2746 4862 2748
rect 4918 2746 4942 2748
rect 4998 2746 5004 2748
rect 4758 2694 4760 2746
rect 4940 2694 4942 2746
rect 4696 2692 4702 2694
rect 4758 2692 4782 2694
rect 4838 2692 4862 2694
rect 4918 2692 4942 2694
rect 4998 2692 5004 2694
rect 4696 2683 5004 2692
rect 5276 2446 5304 4270
rect 5354 4200 5410 5000
rect 5814 4200 5870 5000
rect 6274 4298 6330 5000
rect 6274 4270 6408 4298
rect 6274 4200 6330 4270
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 5080 2372 5132 2378
rect 5080 2314 5132 2320
rect 3799 2204 4107 2213
rect 3799 2202 3805 2204
rect 3861 2202 3885 2204
rect 3941 2202 3965 2204
rect 4021 2202 4045 2204
rect 4101 2202 4107 2204
rect 3861 2150 3863 2202
rect 4043 2150 4045 2202
rect 3799 2148 3805 2150
rect 3861 2148 3885 2150
rect 3941 2148 3965 2150
rect 4021 2148 4045 2150
rect 4101 2148 4107 2150
rect 3799 2139 4107 2148
rect 3700 2032 3752 2038
rect 3700 1974 3752 1980
rect 4160 1896 4212 1902
rect 4160 1838 4212 1844
rect 3799 1116 4107 1125
rect 3799 1114 3805 1116
rect 3861 1114 3885 1116
rect 3941 1114 3965 1116
rect 4021 1114 4045 1116
rect 4101 1114 4107 1116
rect 3861 1062 3863 1114
rect 4043 1062 4045 1114
rect 3799 1060 3805 1062
rect 3861 1060 3885 1062
rect 3941 1060 3965 1062
rect 4021 1060 4045 1062
rect 4101 1060 4107 1062
rect 3799 1051 4107 1060
rect 4172 898 4200 1838
rect 3988 870 4200 898
rect 3988 800 4016 870
rect 4448 800 4476 2314
rect 4696 1660 5004 1669
rect 4696 1658 4702 1660
rect 4758 1658 4782 1660
rect 4838 1658 4862 1660
rect 4918 1658 4942 1660
rect 4998 1658 5004 1660
rect 4758 1606 4760 1658
rect 4940 1606 4942 1658
rect 4696 1604 4702 1606
rect 4758 1604 4782 1606
rect 4838 1604 4862 1606
rect 4918 1604 4942 1606
rect 4998 1604 5004 1606
rect 4696 1595 5004 1604
rect 5092 1170 5120 2314
rect 5368 2038 5396 4200
rect 5828 3618 5856 4200
rect 5828 3590 6040 3618
rect 5592 3292 5900 3301
rect 5592 3290 5598 3292
rect 5654 3290 5678 3292
rect 5734 3290 5758 3292
rect 5814 3290 5838 3292
rect 5894 3290 5900 3292
rect 5654 3238 5656 3290
rect 5836 3238 5838 3290
rect 5592 3236 5598 3238
rect 5654 3236 5678 3238
rect 5734 3236 5758 3238
rect 5814 3236 5838 3238
rect 5894 3236 5900 3238
rect 5592 3227 5900 3236
rect 6012 3126 6040 3590
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5592 2204 5900 2213
rect 5592 2202 5598 2204
rect 5654 2202 5678 2204
rect 5734 2202 5758 2204
rect 5814 2202 5838 2204
rect 5894 2202 5900 2204
rect 5654 2150 5656 2202
rect 5836 2150 5838 2202
rect 5592 2148 5598 2150
rect 5654 2148 5678 2150
rect 5734 2148 5758 2150
rect 5814 2148 5838 2150
rect 5894 2148 5900 2150
rect 5592 2139 5900 2148
rect 5356 2032 5408 2038
rect 5356 1974 5408 1980
rect 5356 1896 5408 1902
rect 5356 1838 5408 1844
rect 4908 1142 5120 1170
rect 4908 800 4936 1142
rect 5368 800 5396 1838
rect 5592 1116 5900 1125
rect 5592 1114 5598 1116
rect 5654 1114 5678 1116
rect 5734 1114 5758 1116
rect 5814 1114 5838 1116
rect 5894 1114 5900 1116
rect 5654 1062 5656 1114
rect 5836 1062 5838 1114
rect 5592 1060 5598 1062
rect 5654 1060 5678 1062
rect 5734 1060 5758 1062
rect 5814 1060 5838 1062
rect 5894 1060 5900 1062
rect 5592 1051 5900 1060
rect 6012 898 6040 2926
rect 6380 1358 6408 4270
rect 6734 4200 6790 5000
rect 7194 4200 7250 5000
rect 6748 4026 6776 4200
rect 6748 3998 6868 4026
rect 6489 3836 6797 3845
rect 6489 3834 6495 3836
rect 6551 3834 6575 3836
rect 6631 3834 6655 3836
rect 6711 3834 6735 3836
rect 6791 3834 6797 3836
rect 6551 3782 6553 3834
rect 6733 3782 6735 3834
rect 6489 3780 6495 3782
rect 6551 3780 6575 3782
rect 6631 3780 6655 3782
rect 6711 3780 6735 3782
rect 6791 3780 6797 3782
rect 6489 3771 6797 3780
rect 6840 3534 6868 3998
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6489 2748 6797 2757
rect 6489 2746 6495 2748
rect 6551 2746 6575 2748
rect 6631 2746 6655 2748
rect 6711 2746 6735 2748
rect 6791 2746 6797 2748
rect 6551 2694 6553 2746
rect 6733 2694 6735 2746
rect 6489 2692 6495 2694
rect 6551 2692 6575 2694
rect 6631 2692 6655 2694
rect 6711 2692 6735 2694
rect 6791 2692 6797 2694
rect 6489 2683 6797 2692
rect 6489 1660 6797 1669
rect 6489 1658 6495 1660
rect 6551 1658 6575 1660
rect 6631 1658 6655 1660
rect 6711 1658 6735 1660
rect 6791 1658 6797 1660
rect 6551 1606 6553 1658
rect 6733 1606 6735 1658
rect 6489 1604 6495 1606
rect 6551 1604 6575 1606
rect 6631 1604 6655 1606
rect 6711 1604 6735 1606
rect 6791 1604 6797 1606
rect 6489 1595 6797 1604
rect 6840 1442 6868 3334
rect 6748 1414 6868 1442
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6276 1284 6328 1290
rect 6276 1226 6328 1232
rect 5828 870 6040 898
rect 5828 800 5856 870
rect 6288 800 6316 1226
rect 6748 800 6776 1414
rect 7208 1358 7236 4200
rect 7385 3292 7693 3301
rect 7385 3290 7391 3292
rect 7447 3290 7471 3292
rect 7527 3290 7551 3292
rect 7607 3290 7631 3292
rect 7687 3290 7693 3292
rect 7447 3238 7449 3290
rect 7629 3238 7631 3290
rect 7385 3236 7391 3238
rect 7447 3236 7471 3238
rect 7527 3236 7551 3238
rect 7607 3236 7631 3238
rect 7687 3236 7693 3238
rect 7385 3227 7693 3236
rect 7385 2204 7693 2213
rect 7385 2202 7391 2204
rect 7447 2202 7471 2204
rect 7527 2202 7551 2204
rect 7607 2202 7631 2204
rect 7687 2202 7693 2204
rect 7447 2150 7449 2202
rect 7629 2150 7631 2202
rect 7385 2148 7391 2150
rect 7447 2148 7471 2150
rect 7527 2148 7551 2150
rect 7607 2148 7631 2150
rect 7687 2148 7693 2150
rect 7385 2139 7693 2148
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 7208 800 7236 1158
rect 7385 1116 7693 1125
rect 7385 1114 7391 1116
rect 7447 1114 7471 1116
rect 7527 1114 7551 1116
rect 7607 1114 7631 1116
rect 7687 1114 7693 1116
rect 7447 1062 7449 1114
rect 7629 1062 7631 1114
rect 7385 1060 7391 1062
rect 7447 1060 7471 1062
rect 7527 1060 7551 1062
rect 7607 1060 7631 1062
rect 7687 1060 7693 1062
rect 7385 1051 7693 1060
rect 2792 734 3004 762
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
<< via2 >>
rect 1116 3834 1172 3836
rect 1196 3834 1252 3836
rect 1276 3834 1332 3836
rect 1356 3834 1412 3836
rect 1116 3782 1162 3834
rect 1162 3782 1172 3834
rect 1196 3782 1226 3834
rect 1226 3782 1238 3834
rect 1238 3782 1252 3834
rect 1276 3782 1290 3834
rect 1290 3782 1302 3834
rect 1302 3782 1332 3834
rect 1356 3782 1366 3834
rect 1366 3782 1412 3834
rect 1116 3780 1172 3782
rect 1196 3780 1252 3782
rect 1276 3780 1332 3782
rect 1356 3780 1412 3782
rect 1116 2746 1172 2748
rect 1196 2746 1252 2748
rect 1276 2746 1332 2748
rect 1356 2746 1412 2748
rect 1116 2694 1162 2746
rect 1162 2694 1172 2746
rect 1196 2694 1226 2746
rect 1226 2694 1238 2746
rect 1238 2694 1252 2746
rect 1276 2694 1290 2746
rect 1290 2694 1302 2746
rect 1302 2694 1332 2746
rect 1356 2694 1366 2746
rect 1366 2694 1412 2746
rect 1116 2692 1172 2694
rect 1196 2692 1252 2694
rect 1276 2692 1332 2694
rect 1356 2692 1412 2694
rect 2012 3290 2068 3292
rect 2092 3290 2148 3292
rect 2172 3290 2228 3292
rect 2252 3290 2308 3292
rect 2012 3238 2058 3290
rect 2058 3238 2068 3290
rect 2092 3238 2122 3290
rect 2122 3238 2134 3290
rect 2134 3238 2148 3290
rect 2172 3238 2186 3290
rect 2186 3238 2198 3290
rect 2198 3238 2228 3290
rect 2252 3238 2262 3290
rect 2262 3238 2308 3290
rect 2012 3236 2068 3238
rect 2092 3236 2148 3238
rect 2172 3236 2228 3238
rect 2252 3236 2308 3238
rect 2012 2202 2068 2204
rect 2092 2202 2148 2204
rect 2172 2202 2228 2204
rect 2252 2202 2308 2204
rect 2012 2150 2058 2202
rect 2058 2150 2068 2202
rect 2092 2150 2122 2202
rect 2122 2150 2134 2202
rect 2134 2150 2148 2202
rect 2172 2150 2186 2202
rect 2186 2150 2198 2202
rect 2198 2150 2228 2202
rect 2252 2150 2262 2202
rect 2262 2150 2308 2202
rect 2012 2148 2068 2150
rect 2092 2148 2148 2150
rect 2172 2148 2228 2150
rect 2252 2148 2308 2150
rect 1116 1658 1172 1660
rect 1196 1658 1252 1660
rect 1276 1658 1332 1660
rect 1356 1658 1412 1660
rect 1116 1606 1162 1658
rect 1162 1606 1172 1658
rect 1196 1606 1226 1658
rect 1226 1606 1238 1658
rect 1238 1606 1252 1658
rect 1276 1606 1290 1658
rect 1290 1606 1302 1658
rect 1302 1606 1332 1658
rect 1356 1606 1366 1658
rect 1366 1606 1412 1658
rect 1116 1604 1172 1606
rect 1196 1604 1252 1606
rect 1276 1604 1332 1606
rect 1356 1604 1412 1606
rect 2012 1114 2068 1116
rect 2092 1114 2148 1116
rect 2172 1114 2228 1116
rect 2252 1114 2308 1116
rect 2012 1062 2058 1114
rect 2058 1062 2068 1114
rect 2092 1062 2122 1114
rect 2122 1062 2134 1114
rect 2134 1062 2148 1114
rect 2172 1062 2186 1114
rect 2186 1062 2198 1114
rect 2198 1062 2228 1114
rect 2252 1062 2262 1114
rect 2262 1062 2308 1114
rect 2012 1060 2068 1062
rect 2092 1060 2148 1062
rect 2172 1060 2228 1062
rect 2252 1060 2308 1062
rect 2909 3834 2965 3836
rect 2989 3834 3045 3836
rect 3069 3834 3125 3836
rect 3149 3834 3205 3836
rect 2909 3782 2955 3834
rect 2955 3782 2965 3834
rect 2989 3782 3019 3834
rect 3019 3782 3031 3834
rect 3031 3782 3045 3834
rect 3069 3782 3083 3834
rect 3083 3782 3095 3834
rect 3095 3782 3125 3834
rect 3149 3782 3159 3834
rect 3159 3782 3205 3834
rect 2909 3780 2965 3782
rect 2989 3780 3045 3782
rect 3069 3780 3125 3782
rect 3149 3780 3205 3782
rect 2909 2746 2965 2748
rect 2989 2746 3045 2748
rect 3069 2746 3125 2748
rect 3149 2746 3205 2748
rect 2909 2694 2955 2746
rect 2955 2694 2965 2746
rect 2989 2694 3019 2746
rect 3019 2694 3031 2746
rect 3031 2694 3045 2746
rect 3069 2694 3083 2746
rect 3083 2694 3095 2746
rect 3095 2694 3125 2746
rect 3149 2694 3159 2746
rect 3159 2694 3205 2746
rect 2909 2692 2965 2694
rect 2989 2692 3045 2694
rect 3069 2692 3125 2694
rect 3149 2692 3205 2694
rect 2909 1658 2965 1660
rect 2989 1658 3045 1660
rect 3069 1658 3125 1660
rect 3149 1658 3205 1660
rect 2909 1606 2955 1658
rect 2955 1606 2965 1658
rect 2989 1606 3019 1658
rect 3019 1606 3031 1658
rect 3031 1606 3045 1658
rect 3069 1606 3083 1658
rect 3083 1606 3095 1658
rect 3095 1606 3125 1658
rect 3149 1606 3159 1658
rect 3159 1606 3205 1658
rect 2909 1604 2965 1606
rect 2989 1604 3045 1606
rect 3069 1604 3125 1606
rect 3149 1604 3205 1606
rect 3805 3290 3861 3292
rect 3885 3290 3941 3292
rect 3965 3290 4021 3292
rect 4045 3290 4101 3292
rect 3805 3238 3851 3290
rect 3851 3238 3861 3290
rect 3885 3238 3915 3290
rect 3915 3238 3927 3290
rect 3927 3238 3941 3290
rect 3965 3238 3979 3290
rect 3979 3238 3991 3290
rect 3991 3238 4021 3290
rect 4045 3238 4055 3290
rect 4055 3238 4101 3290
rect 3805 3236 3861 3238
rect 3885 3236 3941 3238
rect 3965 3236 4021 3238
rect 4045 3236 4101 3238
rect 4702 3834 4758 3836
rect 4782 3834 4838 3836
rect 4862 3834 4918 3836
rect 4942 3834 4998 3836
rect 4702 3782 4748 3834
rect 4748 3782 4758 3834
rect 4782 3782 4812 3834
rect 4812 3782 4824 3834
rect 4824 3782 4838 3834
rect 4862 3782 4876 3834
rect 4876 3782 4888 3834
rect 4888 3782 4918 3834
rect 4942 3782 4952 3834
rect 4952 3782 4998 3834
rect 4702 3780 4758 3782
rect 4782 3780 4838 3782
rect 4862 3780 4918 3782
rect 4942 3780 4998 3782
rect 4702 2746 4758 2748
rect 4782 2746 4838 2748
rect 4862 2746 4918 2748
rect 4942 2746 4998 2748
rect 4702 2694 4748 2746
rect 4748 2694 4758 2746
rect 4782 2694 4812 2746
rect 4812 2694 4824 2746
rect 4824 2694 4838 2746
rect 4862 2694 4876 2746
rect 4876 2694 4888 2746
rect 4888 2694 4918 2746
rect 4942 2694 4952 2746
rect 4952 2694 4998 2746
rect 4702 2692 4758 2694
rect 4782 2692 4838 2694
rect 4862 2692 4918 2694
rect 4942 2692 4998 2694
rect 3805 2202 3861 2204
rect 3885 2202 3941 2204
rect 3965 2202 4021 2204
rect 4045 2202 4101 2204
rect 3805 2150 3851 2202
rect 3851 2150 3861 2202
rect 3885 2150 3915 2202
rect 3915 2150 3927 2202
rect 3927 2150 3941 2202
rect 3965 2150 3979 2202
rect 3979 2150 3991 2202
rect 3991 2150 4021 2202
rect 4045 2150 4055 2202
rect 4055 2150 4101 2202
rect 3805 2148 3861 2150
rect 3885 2148 3941 2150
rect 3965 2148 4021 2150
rect 4045 2148 4101 2150
rect 3805 1114 3861 1116
rect 3885 1114 3941 1116
rect 3965 1114 4021 1116
rect 4045 1114 4101 1116
rect 3805 1062 3851 1114
rect 3851 1062 3861 1114
rect 3885 1062 3915 1114
rect 3915 1062 3927 1114
rect 3927 1062 3941 1114
rect 3965 1062 3979 1114
rect 3979 1062 3991 1114
rect 3991 1062 4021 1114
rect 4045 1062 4055 1114
rect 4055 1062 4101 1114
rect 3805 1060 3861 1062
rect 3885 1060 3941 1062
rect 3965 1060 4021 1062
rect 4045 1060 4101 1062
rect 4702 1658 4758 1660
rect 4782 1658 4838 1660
rect 4862 1658 4918 1660
rect 4942 1658 4998 1660
rect 4702 1606 4748 1658
rect 4748 1606 4758 1658
rect 4782 1606 4812 1658
rect 4812 1606 4824 1658
rect 4824 1606 4838 1658
rect 4862 1606 4876 1658
rect 4876 1606 4888 1658
rect 4888 1606 4918 1658
rect 4942 1606 4952 1658
rect 4952 1606 4998 1658
rect 4702 1604 4758 1606
rect 4782 1604 4838 1606
rect 4862 1604 4918 1606
rect 4942 1604 4998 1606
rect 5598 3290 5654 3292
rect 5678 3290 5734 3292
rect 5758 3290 5814 3292
rect 5838 3290 5894 3292
rect 5598 3238 5644 3290
rect 5644 3238 5654 3290
rect 5678 3238 5708 3290
rect 5708 3238 5720 3290
rect 5720 3238 5734 3290
rect 5758 3238 5772 3290
rect 5772 3238 5784 3290
rect 5784 3238 5814 3290
rect 5838 3238 5848 3290
rect 5848 3238 5894 3290
rect 5598 3236 5654 3238
rect 5678 3236 5734 3238
rect 5758 3236 5814 3238
rect 5838 3236 5894 3238
rect 5598 2202 5654 2204
rect 5678 2202 5734 2204
rect 5758 2202 5814 2204
rect 5838 2202 5894 2204
rect 5598 2150 5644 2202
rect 5644 2150 5654 2202
rect 5678 2150 5708 2202
rect 5708 2150 5720 2202
rect 5720 2150 5734 2202
rect 5758 2150 5772 2202
rect 5772 2150 5784 2202
rect 5784 2150 5814 2202
rect 5838 2150 5848 2202
rect 5848 2150 5894 2202
rect 5598 2148 5654 2150
rect 5678 2148 5734 2150
rect 5758 2148 5814 2150
rect 5838 2148 5894 2150
rect 5598 1114 5654 1116
rect 5678 1114 5734 1116
rect 5758 1114 5814 1116
rect 5838 1114 5894 1116
rect 5598 1062 5644 1114
rect 5644 1062 5654 1114
rect 5678 1062 5708 1114
rect 5708 1062 5720 1114
rect 5720 1062 5734 1114
rect 5758 1062 5772 1114
rect 5772 1062 5784 1114
rect 5784 1062 5814 1114
rect 5838 1062 5848 1114
rect 5848 1062 5894 1114
rect 5598 1060 5654 1062
rect 5678 1060 5734 1062
rect 5758 1060 5814 1062
rect 5838 1060 5894 1062
rect 6495 3834 6551 3836
rect 6575 3834 6631 3836
rect 6655 3834 6711 3836
rect 6735 3834 6791 3836
rect 6495 3782 6541 3834
rect 6541 3782 6551 3834
rect 6575 3782 6605 3834
rect 6605 3782 6617 3834
rect 6617 3782 6631 3834
rect 6655 3782 6669 3834
rect 6669 3782 6681 3834
rect 6681 3782 6711 3834
rect 6735 3782 6745 3834
rect 6745 3782 6791 3834
rect 6495 3780 6551 3782
rect 6575 3780 6631 3782
rect 6655 3780 6711 3782
rect 6735 3780 6791 3782
rect 6495 2746 6551 2748
rect 6575 2746 6631 2748
rect 6655 2746 6711 2748
rect 6735 2746 6791 2748
rect 6495 2694 6541 2746
rect 6541 2694 6551 2746
rect 6575 2694 6605 2746
rect 6605 2694 6617 2746
rect 6617 2694 6631 2746
rect 6655 2694 6669 2746
rect 6669 2694 6681 2746
rect 6681 2694 6711 2746
rect 6735 2694 6745 2746
rect 6745 2694 6791 2746
rect 6495 2692 6551 2694
rect 6575 2692 6631 2694
rect 6655 2692 6711 2694
rect 6735 2692 6791 2694
rect 6495 1658 6551 1660
rect 6575 1658 6631 1660
rect 6655 1658 6711 1660
rect 6735 1658 6791 1660
rect 6495 1606 6541 1658
rect 6541 1606 6551 1658
rect 6575 1606 6605 1658
rect 6605 1606 6617 1658
rect 6617 1606 6631 1658
rect 6655 1606 6669 1658
rect 6669 1606 6681 1658
rect 6681 1606 6711 1658
rect 6735 1606 6745 1658
rect 6745 1606 6791 1658
rect 6495 1604 6551 1606
rect 6575 1604 6631 1606
rect 6655 1604 6711 1606
rect 6735 1604 6791 1606
rect 7391 3290 7447 3292
rect 7471 3290 7527 3292
rect 7551 3290 7607 3292
rect 7631 3290 7687 3292
rect 7391 3238 7437 3290
rect 7437 3238 7447 3290
rect 7471 3238 7501 3290
rect 7501 3238 7513 3290
rect 7513 3238 7527 3290
rect 7551 3238 7565 3290
rect 7565 3238 7577 3290
rect 7577 3238 7607 3290
rect 7631 3238 7641 3290
rect 7641 3238 7687 3290
rect 7391 3236 7447 3238
rect 7471 3236 7527 3238
rect 7551 3236 7607 3238
rect 7631 3236 7687 3238
rect 7391 2202 7447 2204
rect 7471 2202 7527 2204
rect 7551 2202 7607 2204
rect 7631 2202 7687 2204
rect 7391 2150 7437 2202
rect 7437 2150 7447 2202
rect 7471 2150 7501 2202
rect 7501 2150 7513 2202
rect 7513 2150 7527 2202
rect 7551 2150 7565 2202
rect 7565 2150 7577 2202
rect 7577 2150 7607 2202
rect 7631 2150 7641 2202
rect 7641 2150 7687 2202
rect 7391 2148 7447 2150
rect 7471 2148 7527 2150
rect 7551 2148 7607 2150
rect 7631 2148 7687 2150
rect 7391 1114 7447 1116
rect 7471 1114 7527 1116
rect 7551 1114 7607 1116
rect 7631 1114 7687 1116
rect 7391 1062 7437 1114
rect 7437 1062 7447 1114
rect 7471 1062 7501 1114
rect 7501 1062 7513 1114
rect 7513 1062 7527 1114
rect 7551 1062 7565 1114
rect 7565 1062 7577 1114
rect 7577 1062 7607 1114
rect 7631 1062 7641 1114
rect 7641 1062 7687 1114
rect 7391 1060 7447 1062
rect 7471 1060 7527 1062
rect 7551 1060 7607 1062
rect 7631 1060 7687 1062
<< metal3 >>
rect 1106 3840 1422 3841
rect 1106 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1272 3840
rect 1336 3776 1352 3840
rect 1416 3776 1422 3840
rect 1106 3775 1422 3776
rect 2899 3840 3215 3841
rect 2899 3776 2905 3840
rect 2969 3776 2985 3840
rect 3049 3776 3065 3840
rect 3129 3776 3145 3840
rect 3209 3776 3215 3840
rect 2899 3775 3215 3776
rect 4692 3840 5008 3841
rect 4692 3776 4698 3840
rect 4762 3776 4778 3840
rect 4842 3776 4858 3840
rect 4922 3776 4938 3840
rect 5002 3776 5008 3840
rect 4692 3775 5008 3776
rect 6485 3840 6801 3841
rect 6485 3776 6491 3840
rect 6555 3776 6571 3840
rect 6635 3776 6651 3840
rect 6715 3776 6731 3840
rect 6795 3776 6801 3840
rect 6485 3775 6801 3776
rect 2002 3296 2318 3297
rect 2002 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2168 3296
rect 2232 3232 2248 3296
rect 2312 3232 2318 3296
rect 2002 3231 2318 3232
rect 3795 3296 4111 3297
rect 3795 3232 3801 3296
rect 3865 3232 3881 3296
rect 3945 3232 3961 3296
rect 4025 3232 4041 3296
rect 4105 3232 4111 3296
rect 3795 3231 4111 3232
rect 5588 3296 5904 3297
rect 5588 3232 5594 3296
rect 5658 3232 5674 3296
rect 5738 3232 5754 3296
rect 5818 3232 5834 3296
rect 5898 3232 5904 3296
rect 5588 3231 5904 3232
rect 7381 3296 7697 3297
rect 7381 3232 7387 3296
rect 7451 3232 7467 3296
rect 7531 3232 7547 3296
rect 7611 3232 7627 3296
rect 7691 3232 7697 3296
rect 7381 3231 7697 3232
rect 1106 2752 1422 2753
rect 1106 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1272 2752
rect 1336 2688 1352 2752
rect 1416 2688 1422 2752
rect 1106 2687 1422 2688
rect 2899 2752 3215 2753
rect 2899 2688 2905 2752
rect 2969 2688 2985 2752
rect 3049 2688 3065 2752
rect 3129 2688 3145 2752
rect 3209 2688 3215 2752
rect 2899 2687 3215 2688
rect 4692 2752 5008 2753
rect 4692 2688 4698 2752
rect 4762 2688 4778 2752
rect 4842 2688 4858 2752
rect 4922 2688 4938 2752
rect 5002 2688 5008 2752
rect 4692 2687 5008 2688
rect 6485 2752 6801 2753
rect 6485 2688 6491 2752
rect 6555 2688 6571 2752
rect 6635 2688 6651 2752
rect 6715 2688 6731 2752
rect 6795 2688 6801 2752
rect 6485 2687 6801 2688
rect 2002 2208 2318 2209
rect 2002 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2168 2208
rect 2232 2144 2248 2208
rect 2312 2144 2318 2208
rect 2002 2143 2318 2144
rect 3795 2208 4111 2209
rect 3795 2144 3801 2208
rect 3865 2144 3881 2208
rect 3945 2144 3961 2208
rect 4025 2144 4041 2208
rect 4105 2144 4111 2208
rect 3795 2143 4111 2144
rect 5588 2208 5904 2209
rect 5588 2144 5594 2208
rect 5658 2144 5674 2208
rect 5738 2144 5754 2208
rect 5818 2144 5834 2208
rect 5898 2144 5904 2208
rect 5588 2143 5904 2144
rect 7381 2208 7697 2209
rect 7381 2144 7387 2208
rect 7451 2144 7467 2208
rect 7531 2144 7547 2208
rect 7611 2144 7627 2208
rect 7691 2144 7697 2208
rect 7381 2143 7697 2144
rect 1106 1664 1422 1665
rect 1106 1600 1112 1664
rect 1176 1600 1192 1664
rect 1256 1600 1272 1664
rect 1336 1600 1352 1664
rect 1416 1600 1422 1664
rect 1106 1599 1422 1600
rect 2899 1664 3215 1665
rect 2899 1600 2905 1664
rect 2969 1600 2985 1664
rect 3049 1600 3065 1664
rect 3129 1600 3145 1664
rect 3209 1600 3215 1664
rect 2899 1599 3215 1600
rect 4692 1664 5008 1665
rect 4692 1600 4698 1664
rect 4762 1600 4778 1664
rect 4842 1600 4858 1664
rect 4922 1600 4938 1664
rect 5002 1600 5008 1664
rect 4692 1599 5008 1600
rect 6485 1664 6801 1665
rect 6485 1600 6491 1664
rect 6555 1600 6571 1664
rect 6635 1600 6651 1664
rect 6715 1600 6731 1664
rect 6795 1600 6801 1664
rect 6485 1599 6801 1600
rect 2002 1120 2318 1121
rect 2002 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2168 1120
rect 2232 1056 2248 1120
rect 2312 1056 2318 1120
rect 2002 1055 2318 1056
rect 3795 1120 4111 1121
rect 3795 1056 3801 1120
rect 3865 1056 3881 1120
rect 3945 1056 3961 1120
rect 4025 1056 4041 1120
rect 4105 1056 4111 1120
rect 3795 1055 4111 1056
rect 5588 1120 5904 1121
rect 5588 1056 5594 1120
rect 5658 1056 5674 1120
rect 5738 1056 5754 1120
rect 5818 1056 5834 1120
rect 5898 1056 5904 1120
rect 5588 1055 5904 1056
rect 7381 1120 7697 1121
rect 7381 1056 7387 1120
rect 7451 1056 7467 1120
rect 7531 1056 7547 1120
rect 7611 1056 7627 1120
rect 7691 1056 7697 1120
rect 7381 1055 7697 1056
<< via3 >>
rect 1112 3836 1176 3840
rect 1112 3780 1116 3836
rect 1116 3780 1172 3836
rect 1172 3780 1176 3836
rect 1112 3776 1176 3780
rect 1192 3836 1256 3840
rect 1192 3780 1196 3836
rect 1196 3780 1252 3836
rect 1252 3780 1256 3836
rect 1192 3776 1256 3780
rect 1272 3836 1336 3840
rect 1272 3780 1276 3836
rect 1276 3780 1332 3836
rect 1332 3780 1336 3836
rect 1272 3776 1336 3780
rect 1352 3836 1416 3840
rect 1352 3780 1356 3836
rect 1356 3780 1412 3836
rect 1412 3780 1416 3836
rect 1352 3776 1416 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 2985 3836 3049 3840
rect 2985 3780 2989 3836
rect 2989 3780 3045 3836
rect 3045 3780 3049 3836
rect 2985 3776 3049 3780
rect 3065 3836 3129 3840
rect 3065 3780 3069 3836
rect 3069 3780 3125 3836
rect 3125 3780 3129 3836
rect 3065 3776 3129 3780
rect 3145 3836 3209 3840
rect 3145 3780 3149 3836
rect 3149 3780 3205 3836
rect 3205 3780 3209 3836
rect 3145 3776 3209 3780
rect 4698 3836 4762 3840
rect 4698 3780 4702 3836
rect 4702 3780 4758 3836
rect 4758 3780 4762 3836
rect 4698 3776 4762 3780
rect 4778 3836 4842 3840
rect 4778 3780 4782 3836
rect 4782 3780 4838 3836
rect 4838 3780 4842 3836
rect 4778 3776 4842 3780
rect 4858 3836 4922 3840
rect 4858 3780 4862 3836
rect 4862 3780 4918 3836
rect 4918 3780 4922 3836
rect 4858 3776 4922 3780
rect 4938 3836 5002 3840
rect 4938 3780 4942 3836
rect 4942 3780 4998 3836
rect 4998 3780 5002 3836
rect 4938 3776 5002 3780
rect 6491 3836 6555 3840
rect 6491 3780 6495 3836
rect 6495 3780 6551 3836
rect 6551 3780 6555 3836
rect 6491 3776 6555 3780
rect 6571 3836 6635 3840
rect 6571 3780 6575 3836
rect 6575 3780 6631 3836
rect 6631 3780 6635 3836
rect 6571 3776 6635 3780
rect 6651 3836 6715 3840
rect 6651 3780 6655 3836
rect 6655 3780 6711 3836
rect 6711 3780 6715 3836
rect 6651 3776 6715 3780
rect 6731 3836 6795 3840
rect 6731 3780 6735 3836
rect 6735 3780 6791 3836
rect 6791 3780 6795 3836
rect 6731 3776 6795 3780
rect 2008 3292 2072 3296
rect 2008 3236 2012 3292
rect 2012 3236 2068 3292
rect 2068 3236 2072 3292
rect 2008 3232 2072 3236
rect 2088 3292 2152 3296
rect 2088 3236 2092 3292
rect 2092 3236 2148 3292
rect 2148 3236 2152 3292
rect 2088 3232 2152 3236
rect 2168 3292 2232 3296
rect 2168 3236 2172 3292
rect 2172 3236 2228 3292
rect 2228 3236 2232 3292
rect 2168 3232 2232 3236
rect 2248 3292 2312 3296
rect 2248 3236 2252 3292
rect 2252 3236 2308 3292
rect 2308 3236 2312 3292
rect 2248 3232 2312 3236
rect 3801 3292 3865 3296
rect 3801 3236 3805 3292
rect 3805 3236 3861 3292
rect 3861 3236 3865 3292
rect 3801 3232 3865 3236
rect 3881 3292 3945 3296
rect 3881 3236 3885 3292
rect 3885 3236 3941 3292
rect 3941 3236 3945 3292
rect 3881 3232 3945 3236
rect 3961 3292 4025 3296
rect 3961 3236 3965 3292
rect 3965 3236 4021 3292
rect 4021 3236 4025 3292
rect 3961 3232 4025 3236
rect 4041 3292 4105 3296
rect 4041 3236 4045 3292
rect 4045 3236 4101 3292
rect 4101 3236 4105 3292
rect 4041 3232 4105 3236
rect 5594 3292 5658 3296
rect 5594 3236 5598 3292
rect 5598 3236 5654 3292
rect 5654 3236 5658 3292
rect 5594 3232 5658 3236
rect 5674 3292 5738 3296
rect 5674 3236 5678 3292
rect 5678 3236 5734 3292
rect 5734 3236 5738 3292
rect 5674 3232 5738 3236
rect 5754 3292 5818 3296
rect 5754 3236 5758 3292
rect 5758 3236 5814 3292
rect 5814 3236 5818 3292
rect 5754 3232 5818 3236
rect 5834 3292 5898 3296
rect 5834 3236 5838 3292
rect 5838 3236 5894 3292
rect 5894 3236 5898 3292
rect 5834 3232 5898 3236
rect 7387 3292 7451 3296
rect 7387 3236 7391 3292
rect 7391 3236 7447 3292
rect 7447 3236 7451 3292
rect 7387 3232 7451 3236
rect 7467 3292 7531 3296
rect 7467 3236 7471 3292
rect 7471 3236 7527 3292
rect 7527 3236 7531 3292
rect 7467 3232 7531 3236
rect 7547 3292 7611 3296
rect 7547 3236 7551 3292
rect 7551 3236 7607 3292
rect 7607 3236 7611 3292
rect 7547 3232 7611 3236
rect 7627 3292 7691 3296
rect 7627 3236 7631 3292
rect 7631 3236 7687 3292
rect 7687 3236 7691 3292
rect 7627 3232 7691 3236
rect 1112 2748 1176 2752
rect 1112 2692 1116 2748
rect 1116 2692 1172 2748
rect 1172 2692 1176 2748
rect 1112 2688 1176 2692
rect 1192 2748 1256 2752
rect 1192 2692 1196 2748
rect 1196 2692 1252 2748
rect 1252 2692 1256 2748
rect 1192 2688 1256 2692
rect 1272 2748 1336 2752
rect 1272 2692 1276 2748
rect 1276 2692 1332 2748
rect 1332 2692 1336 2748
rect 1272 2688 1336 2692
rect 1352 2748 1416 2752
rect 1352 2692 1356 2748
rect 1356 2692 1412 2748
rect 1412 2692 1416 2748
rect 1352 2688 1416 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 2985 2748 3049 2752
rect 2985 2692 2989 2748
rect 2989 2692 3045 2748
rect 3045 2692 3049 2748
rect 2985 2688 3049 2692
rect 3065 2748 3129 2752
rect 3065 2692 3069 2748
rect 3069 2692 3125 2748
rect 3125 2692 3129 2748
rect 3065 2688 3129 2692
rect 3145 2748 3209 2752
rect 3145 2692 3149 2748
rect 3149 2692 3205 2748
rect 3205 2692 3209 2748
rect 3145 2688 3209 2692
rect 4698 2748 4762 2752
rect 4698 2692 4702 2748
rect 4702 2692 4758 2748
rect 4758 2692 4762 2748
rect 4698 2688 4762 2692
rect 4778 2748 4842 2752
rect 4778 2692 4782 2748
rect 4782 2692 4838 2748
rect 4838 2692 4842 2748
rect 4778 2688 4842 2692
rect 4858 2748 4922 2752
rect 4858 2692 4862 2748
rect 4862 2692 4918 2748
rect 4918 2692 4922 2748
rect 4858 2688 4922 2692
rect 4938 2748 5002 2752
rect 4938 2692 4942 2748
rect 4942 2692 4998 2748
rect 4998 2692 5002 2748
rect 4938 2688 5002 2692
rect 6491 2748 6555 2752
rect 6491 2692 6495 2748
rect 6495 2692 6551 2748
rect 6551 2692 6555 2748
rect 6491 2688 6555 2692
rect 6571 2748 6635 2752
rect 6571 2692 6575 2748
rect 6575 2692 6631 2748
rect 6631 2692 6635 2748
rect 6571 2688 6635 2692
rect 6651 2748 6715 2752
rect 6651 2692 6655 2748
rect 6655 2692 6711 2748
rect 6711 2692 6715 2748
rect 6651 2688 6715 2692
rect 6731 2748 6795 2752
rect 6731 2692 6735 2748
rect 6735 2692 6791 2748
rect 6791 2692 6795 2748
rect 6731 2688 6795 2692
rect 2008 2204 2072 2208
rect 2008 2148 2012 2204
rect 2012 2148 2068 2204
rect 2068 2148 2072 2204
rect 2008 2144 2072 2148
rect 2088 2204 2152 2208
rect 2088 2148 2092 2204
rect 2092 2148 2148 2204
rect 2148 2148 2152 2204
rect 2088 2144 2152 2148
rect 2168 2204 2232 2208
rect 2168 2148 2172 2204
rect 2172 2148 2228 2204
rect 2228 2148 2232 2204
rect 2168 2144 2232 2148
rect 2248 2204 2312 2208
rect 2248 2148 2252 2204
rect 2252 2148 2308 2204
rect 2308 2148 2312 2204
rect 2248 2144 2312 2148
rect 3801 2204 3865 2208
rect 3801 2148 3805 2204
rect 3805 2148 3861 2204
rect 3861 2148 3865 2204
rect 3801 2144 3865 2148
rect 3881 2204 3945 2208
rect 3881 2148 3885 2204
rect 3885 2148 3941 2204
rect 3941 2148 3945 2204
rect 3881 2144 3945 2148
rect 3961 2204 4025 2208
rect 3961 2148 3965 2204
rect 3965 2148 4021 2204
rect 4021 2148 4025 2204
rect 3961 2144 4025 2148
rect 4041 2204 4105 2208
rect 4041 2148 4045 2204
rect 4045 2148 4101 2204
rect 4101 2148 4105 2204
rect 4041 2144 4105 2148
rect 5594 2204 5658 2208
rect 5594 2148 5598 2204
rect 5598 2148 5654 2204
rect 5654 2148 5658 2204
rect 5594 2144 5658 2148
rect 5674 2204 5738 2208
rect 5674 2148 5678 2204
rect 5678 2148 5734 2204
rect 5734 2148 5738 2204
rect 5674 2144 5738 2148
rect 5754 2204 5818 2208
rect 5754 2148 5758 2204
rect 5758 2148 5814 2204
rect 5814 2148 5818 2204
rect 5754 2144 5818 2148
rect 5834 2204 5898 2208
rect 5834 2148 5838 2204
rect 5838 2148 5894 2204
rect 5894 2148 5898 2204
rect 5834 2144 5898 2148
rect 7387 2204 7451 2208
rect 7387 2148 7391 2204
rect 7391 2148 7447 2204
rect 7447 2148 7451 2204
rect 7387 2144 7451 2148
rect 7467 2204 7531 2208
rect 7467 2148 7471 2204
rect 7471 2148 7527 2204
rect 7527 2148 7531 2204
rect 7467 2144 7531 2148
rect 7547 2204 7611 2208
rect 7547 2148 7551 2204
rect 7551 2148 7607 2204
rect 7607 2148 7611 2204
rect 7547 2144 7611 2148
rect 7627 2204 7691 2208
rect 7627 2148 7631 2204
rect 7631 2148 7687 2204
rect 7687 2148 7691 2204
rect 7627 2144 7691 2148
rect 1112 1660 1176 1664
rect 1112 1604 1116 1660
rect 1116 1604 1172 1660
rect 1172 1604 1176 1660
rect 1112 1600 1176 1604
rect 1192 1660 1256 1664
rect 1192 1604 1196 1660
rect 1196 1604 1252 1660
rect 1252 1604 1256 1660
rect 1192 1600 1256 1604
rect 1272 1660 1336 1664
rect 1272 1604 1276 1660
rect 1276 1604 1332 1660
rect 1332 1604 1336 1660
rect 1272 1600 1336 1604
rect 1352 1660 1416 1664
rect 1352 1604 1356 1660
rect 1356 1604 1412 1660
rect 1412 1604 1416 1660
rect 1352 1600 1416 1604
rect 2905 1660 2969 1664
rect 2905 1604 2909 1660
rect 2909 1604 2965 1660
rect 2965 1604 2969 1660
rect 2905 1600 2969 1604
rect 2985 1660 3049 1664
rect 2985 1604 2989 1660
rect 2989 1604 3045 1660
rect 3045 1604 3049 1660
rect 2985 1600 3049 1604
rect 3065 1660 3129 1664
rect 3065 1604 3069 1660
rect 3069 1604 3125 1660
rect 3125 1604 3129 1660
rect 3065 1600 3129 1604
rect 3145 1660 3209 1664
rect 3145 1604 3149 1660
rect 3149 1604 3205 1660
rect 3205 1604 3209 1660
rect 3145 1600 3209 1604
rect 4698 1660 4762 1664
rect 4698 1604 4702 1660
rect 4702 1604 4758 1660
rect 4758 1604 4762 1660
rect 4698 1600 4762 1604
rect 4778 1660 4842 1664
rect 4778 1604 4782 1660
rect 4782 1604 4838 1660
rect 4838 1604 4842 1660
rect 4778 1600 4842 1604
rect 4858 1660 4922 1664
rect 4858 1604 4862 1660
rect 4862 1604 4918 1660
rect 4918 1604 4922 1660
rect 4858 1600 4922 1604
rect 4938 1660 5002 1664
rect 4938 1604 4942 1660
rect 4942 1604 4998 1660
rect 4998 1604 5002 1660
rect 4938 1600 5002 1604
rect 6491 1660 6555 1664
rect 6491 1604 6495 1660
rect 6495 1604 6551 1660
rect 6551 1604 6555 1660
rect 6491 1600 6555 1604
rect 6571 1660 6635 1664
rect 6571 1604 6575 1660
rect 6575 1604 6631 1660
rect 6631 1604 6635 1660
rect 6571 1600 6635 1604
rect 6651 1660 6715 1664
rect 6651 1604 6655 1660
rect 6655 1604 6711 1660
rect 6711 1604 6715 1660
rect 6651 1600 6715 1604
rect 6731 1660 6795 1664
rect 6731 1604 6735 1660
rect 6735 1604 6791 1660
rect 6791 1604 6795 1660
rect 6731 1600 6795 1604
rect 2008 1116 2072 1120
rect 2008 1060 2012 1116
rect 2012 1060 2068 1116
rect 2068 1060 2072 1116
rect 2008 1056 2072 1060
rect 2088 1116 2152 1120
rect 2088 1060 2092 1116
rect 2092 1060 2148 1116
rect 2148 1060 2152 1116
rect 2088 1056 2152 1060
rect 2168 1116 2232 1120
rect 2168 1060 2172 1116
rect 2172 1060 2228 1116
rect 2228 1060 2232 1116
rect 2168 1056 2232 1060
rect 2248 1116 2312 1120
rect 2248 1060 2252 1116
rect 2252 1060 2308 1116
rect 2308 1060 2312 1116
rect 2248 1056 2312 1060
rect 3801 1116 3865 1120
rect 3801 1060 3805 1116
rect 3805 1060 3861 1116
rect 3861 1060 3865 1116
rect 3801 1056 3865 1060
rect 3881 1116 3945 1120
rect 3881 1060 3885 1116
rect 3885 1060 3941 1116
rect 3941 1060 3945 1116
rect 3881 1056 3945 1060
rect 3961 1116 4025 1120
rect 3961 1060 3965 1116
rect 3965 1060 4021 1116
rect 4021 1060 4025 1116
rect 3961 1056 4025 1060
rect 4041 1116 4105 1120
rect 4041 1060 4045 1116
rect 4045 1060 4101 1116
rect 4101 1060 4105 1116
rect 4041 1056 4105 1060
rect 5594 1116 5658 1120
rect 5594 1060 5598 1116
rect 5598 1060 5654 1116
rect 5654 1060 5658 1116
rect 5594 1056 5658 1060
rect 5674 1116 5738 1120
rect 5674 1060 5678 1116
rect 5678 1060 5734 1116
rect 5734 1060 5738 1116
rect 5674 1056 5738 1060
rect 5754 1116 5818 1120
rect 5754 1060 5758 1116
rect 5758 1060 5814 1116
rect 5814 1060 5818 1116
rect 5754 1056 5818 1060
rect 5834 1116 5898 1120
rect 5834 1060 5838 1116
rect 5838 1060 5894 1116
rect 5894 1060 5898 1116
rect 5834 1056 5898 1060
rect 7387 1116 7451 1120
rect 7387 1060 7391 1116
rect 7391 1060 7447 1116
rect 7447 1060 7451 1116
rect 7387 1056 7451 1060
rect 7467 1116 7531 1120
rect 7467 1060 7471 1116
rect 7471 1060 7527 1116
rect 7527 1060 7531 1116
rect 7467 1056 7531 1060
rect 7547 1116 7611 1120
rect 7547 1060 7551 1116
rect 7551 1060 7607 1116
rect 7607 1060 7611 1116
rect 7547 1056 7611 1060
rect 7627 1116 7691 1120
rect 7627 1060 7631 1116
rect 7631 1060 7687 1116
rect 7687 1060 7691 1116
rect 7627 1056 7691 1060
<< metal4 >>
rect 1104 3840 1424 3856
rect 1104 3776 1112 3840
rect 1176 3776 1192 3840
rect 1256 3776 1272 3840
rect 1336 3776 1352 3840
rect 1416 3776 1424 3840
rect 1104 2752 1424 3776
rect 1104 2688 1112 2752
rect 1176 2688 1192 2752
rect 1256 2688 1272 2752
rect 1336 2688 1352 2752
rect 1416 2688 1424 2752
rect 1104 1664 1424 2688
rect 1104 1600 1112 1664
rect 1176 1600 1192 1664
rect 1256 1600 1272 1664
rect 1336 1600 1352 1664
rect 1416 1600 1424 1664
rect 1104 1040 1424 1600
rect 2000 3296 2320 3856
rect 2000 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2168 3296
rect 2232 3232 2248 3296
rect 2312 3232 2320 3296
rect 2000 2208 2320 3232
rect 2000 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2168 2208
rect 2232 2144 2248 2208
rect 2312 2144 2320 2208
rect 2000 1120 2320 2144
rect 2000 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2168 1120
rect 2232 1056 2248 1120
rect 2312 1056 2320 1120
rect 2000 1040 2320 1056
rect 2897 3840 3217 3856
rect 2897 3776 2905 3840
rect 2969 3776 2985 3840
rect 3049 3776 3065 3840
rect 3129 3776 3145 3840
rect 3209 3776 3217 3840
rect 2897 2752 3217 3776
rect 2897 2688 2905 2752
rect 2969 2688 2985 2752
rect 3049 2688 3065 2752
rect 3129 2688 3145 2752
rect 3209 2688 3217 2752
rect 2897 1664 3217 2688
rect 2897 1600 2905 1664
rect 2969 1600 2985 1664
rect 3049 1600 3065 1664
rect 3129 1600 3145 1664
rect 3209 1600 3217 1664
rect 2897 1040 3217 1600
rect 3793 3296 4113 3856
rect 3793 3232 3801 3296
rect 3865 3232 3881 3296
rect 3945 3232 3961 3296
rect 4025 3232 4041 3296
rect 4105 3232 4113 3296
rect 3793 2208 4113 3232
rect 3793 2144 3801 2208
rect 3865 2144 3881 2208
rect 3945 2144 3961 2208
rect 4025 2144 4041 2208
rect 4105 2144 4113 2208
rect 3793 1120 4113 2144
rect 3793 1056 3801 1120
rect 3865 1056 3881 1120
rect 3945 1056 3961 1120
rect 4025 1056 4041 1120
rect 4105 1056 4113 1120
rect 3793 1040 4113 1056
rect 4690 3840 5010 3856
rect 4690 3776 4698 3840
rect 4762 3776 4778 3840
rect 4842 3776 4858 3840
rect 4922 3776 4938 3840
rect 5002 3776 5010 3840
rect 4690 2752 5010 3776
rect 4690 2688 4698 2752
rect 4762 2688 4778 2752
rect 4842 2688 4858 2752
rect 4922 2688 4938 2752
rect 5002 2688 5010 2752
rect 4690 1664 5010 2688
rect 4690 1600 4698 1664
rect 4762 1600 4778 1664
rect 4842 1600 4858 1664
rect 4922 1600 4938 1664
rect 5002 1600 5010 1664
rect 4690 1040 5010 1600
rect 5586 3296 5906 3856
rect 5586 3232 5594 3296
rect 5658 3232 5674 3296
rect 5738 3232 5754 3296
rect 5818 3232 5834 3296
rect 5898 3232 5906 3296
rect 5586 2208 5906 3232
rect 5586 2144 5594 2208
rect 5658 2144 5674 2208
rect 5738 2144 5754 2208
rect 5818 2144 5834 2208
rect 5898 2144 5906 2208
rect 5586 1120 5906 2144
rect 5586 1056 5594 1120
rect 5658 1056 5674 1120
rect 5738 1056 5754 1120
rect 5818 1056 5834 1120
rect 5898 1056 5906 1120
rect 5586 1040 5906 1056
rect 6483 3840 6803 3856
rect 6483 3776 6491 3840
rect 6555 3776 6571 3840
rect 6635 3776 6651 3840
rect 6715 3776 6731 3840
rect 6795 3776 6803 3840
rect 6483 2752 6803 3776
rect 6483 2688 6491 2752
rect 6555 2688 6571 2752
rect 6635 2688 6651 2752
rect 6715 2688 6731 2752
rect 6795 2688 6803 2752
rect 6483 1664 6803 2688
rect 6483 1600 6491 1664
rect 6555 1600 6571 1664
rect 6635 1600 6651 1664
rect 6715 1600 6731 1664
rect 6795 1600 6803 1664
rect 6483 1040 6803 1600
rect 7379 3296 7699 3856
rect 7379 3232 7387 3296
rect 7451 3232 7467 3296
rect 7531 3232 7547 3296
rect 7611 3232 7627 3296
rect 7691 3232 7699 3296
rect 7379 2208 7699 3232
rect 7379 2144 7387 2208
rect 7451 2144 7467 2208
rect 7531 2144 7547 2208
rect 7611 2144 7627 2208
rect 7691 2144 7699 2208
rect 7379 1120 7699 2144
rect 7379 1056 7387 1120
rect 7451 1056 7467 1120
rect 7531 1056 7547 1120
rect 7611 1056 7627 1120
rect 7691 1056 7699 1120
rect 7379 1040 7699 1056
use sky130_fd_sc_hd__clkbuf_8  BUF\[0\] OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1104 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[1\]
timestamp 1665323087
transform 1 0 1104 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[2\]
timestamp 1665323087
transform -1 0 1932 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[3\]
timestamp 1665323087
transform 1 0 1840 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[4\]
timestamp 1665323087
transform -1 0 2760 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[5\]
timestamp 1665323087
transform -1 0 3312 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[6\]
timestamp 1665323087
transform 1 0 3220 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[7\]
timestamp 1665323087
transform 1 0 3680 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[8\]
timestamp 1665323087
transform 1 0 4140 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[9\]
timestamp 1665323087
transform 1 0 5520 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[10\]
timestamp 1665323087
transform 1 0 5796 0 -1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[11\]
timestamp 1665323087
transform 1 0 5796 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[12\]
timestamp 1665323087
transform -1 0 6808 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[13\]
timestamp 1665323087
transform -1 0 6808 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[14\]
timestamp 1665323087
transform -1 0 5336 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 1012 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2116 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1665323087
transform 1 0 2852 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 3036 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 4140 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1665323087
transform 1 0 5336 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1665323087
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1665323087
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1665323087
transform 1 0 7176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1665323087
transform 1 0 1932 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1665323087
transform 1 0 3312 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1665323087
transform 1 0 4692 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1665323087
transform 1 0 5428 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1665323087
transform 1 0 5612 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_70
timestamp 1665323087
transform 1 0 6808 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_74
timestamp 1665323087
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1665323087
transform 1 0 644 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1665323087
transform 1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1665323087
transform 1 0 3036 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1665323087
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_67
timestamp 1665323087
transform 1 0 6532 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1665323087
transform 1 0 644 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1665323087
transform 1 0 1748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1665323087
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_42
timestamp 1665323087
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1665323087
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1665323087
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1665323087
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_74
timestamp 1665323087
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1665323087
transform 1 0 644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1665323087
transform 1 0 1012 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1665323087
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1665323087
transform 1 0 2852 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1665323087
transform 1 0 3036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1665323087
transform 1 0 4140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 1665323087
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1665323087
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1665323087
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_74
timestamp 1665323087
transform 1 0 7176 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1665323087
transform 1 0 368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1665323087
transform -1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1665323087
transform 1 0 368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1665323087
transform -1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1665323087
transform 1 0 368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1665323087
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1665323087
transform 1 0 368 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1665323087
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1665323087
transform 1 0 368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1665323087
transform -1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_10 OL_LATEST/OpenLane/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1665323087
transform 1 0 2944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_11
timestamp 1665323087
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12
timestamp 1665323087
transform 1 0 5520 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1665323087
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1665323087
transform 1 0 5520 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1665323087
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1665323087
transform 1 0 5520 0 1 3264
box -38 -48 130 592
<< labels >>
flabel metal4 s 2000 1040 2320 3856 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3793 1040 4113 3856 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 5586 1040 5906 3856 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7379 1040 7699 3856 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1104 1040 1424 3856 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 2897 1040 3217 3856 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4690 1040 5010 3856 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6483 1040 6803 3856 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2134 4200 2190 5000 0 FreeSans 224 90 0 0 in_n[0]
port 2 nsew signal input
flabel metal2 s 6734 4200 6790 5000 0 FreeSans 224 90 0 0 in_n[10]
port 3 nsew signal input
flabel metal2 s 7194 4200 7250 5000 0 FreeSans 224 90 0 0 in_n[11]
port 4 nsew signal input
flabel metal2 s 2594 4200 2650 5000 0 FreeSans 224 90 0 0 in_n[1]
port 5 nsew signal input
flabel metal2 s 3054 4200 3110 5000 0 FreeSans 224 90 0 0 in_n[2]
port 6 nsew signal input
flabel metal2 s 3514 4200 3570 5000 0 FreeSans 224 90 0 0 in_n[3]
port 7 nsew signal input
flabel metal2 s 3974 4200 4030 5000 0 FreeSans 224 90 0 0 in_n[4]
port 8 nsew signal input
flabel metal2 s 4434 4200 4490 5000 0 FreeSans 224 90 0 0 in_n[5]
port 9 nsew signal input
flabel metal2 s 4894 4200 4950 5000 0 FreeSans 224 90 0 0 in_n[6]
port 10 nsew signal input
flabel metal2 s 5354 4200 5410 5000 0 FreeSans 224 90 0 0 in_n[7]
port 11 nsew signal input
flabel metal2 s 5814 4200 5870 5000 0 FreeSans 224 90 0 0 in_n[8]
port 12 nsew signal input
flabel metal2 s 6274 4200 6330 5000 0 FreeSans 224 90 0 0 in_n[9]
port 13 nsew signal input
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 in_s[0]
port 14 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 in_s[1]
port 15 nsew signal input
flabel metal2 s 1674 0 1730 800 0 FreeSans 224 90 0 0 in_s[2]
port 16 nsew signal input
flabel metal2 s 754 4200 810 5000 0 FreeSans 224 90 0 0 out_n[0]
port 17 nsew signal tristate
flabel metal2 s 1214 4200 1270 5000 0 FreeSans 224 90 0 0 out_n[1]
port 18 nsew signal tristate
flabel metal2 s 1674 4200 1730 5000 0 FreeSans 224 90 0 0 out_n[2]
port 19 nsew signal tristate
flabel metal2 s 2134 0 2190 800 0 FreeSans 224 90 0 0 out_s[0]
port 20 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 out_s[10]
port 21 nsew signal tristate
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 out_s[11]
port 22 nsew signal tristate
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 out_s[1]
port 23 nsew signal tristate
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 out_s[2]
port 24 nsew signal tristate
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 out_s[3]
port 25 nsew signal tristate
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 out_s[4]
port 26 nsew signal tristate
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 out_s[5]
port 27 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 out_s[6]
port 28 nsew signal tristate
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 out_s[7]
port 29 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 out_s[8]
port 30 nsew signal tristate
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 out_s[9]
port 31 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 8000 5000
<< end >>
