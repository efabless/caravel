* NGSPICE file created from gpio_kogic_high.ext - technology: sky130A


* Top level circuit gpio_kogic_high

.end

