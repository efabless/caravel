magic
tech sky130A
magscale 1 2
timestamp 1606502073
<< metal4 >>
rect -3179 3059 3179 3100
rect -3179 -3059 2923 3059
rect 3159 -3059 3179 3059
rect -3179 -3100 3179 -3059
<< via4 >>
rect 2923 -3059 3159 3059
<< mimcap2 >>
rect -3079 2960 2921 3000
rect -3079 -2960 -3039 2960
rect 2289 -2960 2921 2960
rect -3079 -3000 2921 -2960
<< mimcap2contact >>
rect -3039 -2960 2289 2960
<< metal5 >>
rect 2881 3059 3201 3101
rect -3063 2960 2313 2984
rect -3063 -2960 -3039 2960
rect 2289 -2960 2313 2960
rect -3063 -2984 2313 -2960
rect 2881 -3059 2923 3059
rect 3159 -3059 3201 3059
rect 2881 -3101 3201 -3059
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_2
string FIXED_BBOX -3179 -3100 3021 3100
string parameters w 30.00 l 30.00 val 920.4 carea 1.00 cperi 0.17 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov +90
string library sky130
<< end >>
