* NGSPICE file created from spare_logic_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbp_1 abstract view
.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

.subckt spare_logic_block spare_xfq[0] spare_xfq[1] spare_xfqn[0] spare_xfqn[1] spare_xi[0]
+ spare_xi[1] spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0]
+ spare_xna[1] spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12]
+ spare_xz[13] spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19]
+ spare_xz[1] spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25]
+ spare_xz[26] spare_xz[2] spare_xz[3] spare_xz[4] spare_xz[5] spare_xz[6] spare_xz[7]
+ spare_xz[8] spare_xz[9] vccd vssd
XFILLER_0_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_const\[8\] vssd vssd vccd vccd spare_logic_const\[8\]/HI spare_xz[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_nor\[0\] spare_xz[9] spare_xz[11] vssd vssd vccd vccd spare_xno[0] sky130_fd_sc_hd__nor2_2
Xspare_logic_const\[22\] vssd vssd vccd vccd spare_logic_const\[22\]/HI spare_xz[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[15\] vssd vssd vccd vccd spare_logic_const\[15\]/HI spare_xz[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[6\] vssd vssd vccd vccd spare_logic_const\[6\]/HI spare_xz[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[20\] vssd vssd vccd vccd spare_logic_const\[20\]/HI spare_xz[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[13\] vssd vssd vccd vccd spare_logic_const\[13\]/HI spare_xz[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[4\] vssd vssd vccd vccd spare_logic_const\[4\]/HI spare_xz[4]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_flop\[0\] spare_xz[21] spare_xz[19] spare_xz[25] spare_xz[23] vssd vssd
+ vccd vccd spare_xfq[0] spare_xfqn[0] sky130_fd_sc_hd__dfbbp_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_mux\[1\] spare_xz[14] spare_xz[16] spare_xz[18] vssd vssd vccd vccd spare_xmx[1]
+ sky130_fd_sc_hd__mux2_2
Xspare_logic_const\[11\] vssd vssd vccd vccd spare_logic_const\[11\]/HI spare_xz[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[2\] vssd vssd vccd vccd spare_logic_const\[2\]/HI spare_xz[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_44 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[3\] spare_xz[3] vssd vssd vccd vccd spare_xi[3] sky130_fd_sc_hd__inv_2
XFILLER_10_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[0\] vssd vssd vccd vccd spare_logic_const\[0\]/HI spare_xz[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_7_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[1\] spare_xz[1] vssd vssd vccd vccd spare_xi[1] sky130_fd_sc_hd__inv_2
XFILLER_4_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_69 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[25\] vssd vssd vccd vccd spare_logic_const\[25\]/HI spare_xz[25]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_nand\[1\] spare_xz[6] spare_xz[8] vssd vssd vccd vccd spare_xna[1] sky130_fd_sc_hd__nand2_2
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[18\] vssd vssd vccd vccd spare_logic_const\[18\]/HI spare_xz[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[9\] vssd vssd vccd vccd spare_logic_const\[9\]/HI spare_xz[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_8_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xspare_logic_nor\[1\] spare_xz[10] spare_xz[12] vssd vssd vccd vccd spare_xno[1] sky130_fd_sc_hd__nor2_2
XFILLER_7_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[23\] vssd vssd vccd vccd spare_logic_const\[23\]/HI spare_xz[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_30 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xspare_logic_const\[16\] vssd vssd vccd vccd spare_logic_const\[16\]/HI spare_xz[16]
+ sky130_fd_sc_hd__conb_1
XTAP_31 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_32 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xspare_logic_const\[7\] vssd vssd vccd vccd spare_logic_const\[7\]/HI spare_xz[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_biginv spare_xz[4] vssd vssd vccd vccd spare_xib sky130_fd_sc_hd__inv_8
XFILLER_8_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[21\] vssd vssd vccd vccd spare_logic_const\[21\]/HI spare_xz[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XTAP_33 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XTAP_34 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xspare_logic_const\[14\] vssd vssd vccd vccd spare_logic_const\[14\]/HI spare_xz[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_35 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xspare_logic_const\[5\] vssd vssd vccd vccd spare_logic_const\[5\]/HI spare_xz[5]
+ sky130_fd_sc_hd__conb_1
XTAP_24 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_36 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_25 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_flop\[1\] spare_xz[22] spare_xz[20] spare_xz[26] spare_xz[24] vssd vssd
+ vccd vccd spare_xfq[1] spare_xfqn[1] sky130_fd_sc_hd__dfbbp_1
XFILLER_5_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_37 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[12\] vssd vssd vccd vccd spare_logic_const\[12\]/HI spare_xz[12]
+ sky130_fd_sc_hd__conb_1
XTAP_26 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_27 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[3\] vssd vssd vccd vccd spare_logic_const\[3\]/HI spare_xz[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XTAP_28 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xspare_logic_mux\[0\] spare_xz[13] spare_xz[15] spare_xz[17] vssd vssd vccd vccd spare_xmx[0]
+ sky130_fd_sc_hd__mux2_2
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_29 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[10\] vssd vssd vccd vccd spare_logic_const\[10\]/HI spare_xz[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[1\] vssd vssd vccd vccd spare_logic_const\[1\]/HI spare_xz[1]
+ sky130_fd_sc_hd__conb_1
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[2\] spare_xz[2] vssd vssd vccd vccd spare_xi[2] sky130_fd_sc_hd__inv_2
XFILLER_8_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[26\] vssd vssd vccd vccd spare_logic_const\[26\]/HI spare_xz[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[19\] vssd vssd vccd vccd spare_logic_const\[19\]/HI spare_xz[19]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[0\] spare_xz[0] vssd vssd vccd vccd spare_xi[0] sky130_fd_sc_hd__inv_2
XFILLER_9_20 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[24\] vssd vssd vccd vccd spare_logic_const\[24\]/HI spare_xz[24]
+ sky130_fd_sc_hd__conb_1
XFILLER_6_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_nand\[0\] spare_xz[5] spare_xz[7] vssd vssd vccd vccd spare_xna[0] sky130_fd_sc_hd__nand2_2
XFILLER_3_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[17\] vssd vssd vccd vccd spare_logic_const\[17\]/HI spare_xz[17]
+ sky130_fd_sc_hd__conb_1
.ends

