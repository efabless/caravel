VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_signal_buffering
  CLASS BLOCK ;
  FOREIGN gpio_signal_buffering ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN mgmt_io_in_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2082.940 4983.335 2084.530 4983.535 ;
      LAYER mcon ;
        RECT 2082.940 4983.365 2084.030 4983.535 ;
      LAYER met1 ;
        RECT 2082.880 4983.315 2084.090 4983.575 ;
        RECT 2083.245 4976.935 2083.565 4977.055 ;
        RECT 2079.535 4976.795 2083.565 4976.935 ;
      LAYER via ;
        RECT 2082.940 4983.315 2084.030 4983.575 ;
        RECT 2083.275 4976.795 2083.535 4977.055 ;
      LAYER met2 ;
        RECT 2082.940 4983.285 2084.030 4983.605 ;
        RECT 2083.395 4977.085 2083.535 4983.285 ;
        RECT 2083.275 4976.765 2083.535 4977.085 ;
        RECT 2083.395 4976.065 2083.535 4976.765 ;
    END
  END mgmt_io_in_unbuf[11]
  PIN mgmt_io_out_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2084.265 4986.965 2084.435 4987.445 ;
        RECT 2085.105 4986.965 2085.275 4987.445 ;
        RECT 2085.945 4986.965 2086.115 4987.445 ;
        RECT 2086.785 4986.965 2086.955 4987.445 ;
        RECT 2084.265 4986.795 2086.955 4986.965 ;
        RECT 2084.265 4986.255 2084.520 4986.795 ;
        RECT 2084.265 4986.085 2086.955 4986.255 ;
        RECT 2084.265 4985.235 2084.435 4986.085 ;
        RECT 2085.105 4985.235 2085.275 4986.085 ;
        RECT 2085.945 4985.235 2086.115 4986.085 ;
        RECT 2086.785 4985.235 2086.955 4986.085 ;
      LAYER mcon ;
        RECT 2084.350 4986.085 2084.520 4986.935 ;
      LAYER met1 ;
        RECT 2084.310 4986.025 2084.570 4986.995 ;
        RECT 2084.215 4976.375 2084.535 4976.495 ;
        RECT 2080.535 4976.235 2084.535 4976.375 ;
      LAYER via ;
        RECT 2084.310 4986.085 2084.570 4986.935 ;
        RECT 2084.245 4976.235 2084.505 4976.495 ;
      LAYER met2 ;
        RECT 2084.280 4986.085 2084.600 4986.935 ;
        RECT 2084.365 4976.525 2084.505 4986.085 ;
        RECT 2084.245 4976.205 2084.505 4976.525 ;
        RECT 2084.365 4976.065 2084.505 4976.205 ;
    END
  END mgmt_io_out_buf[11]
  PIN mgmt_io_out_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3317.250 4986.555 3317.420 4987.035 ;
        RECT 3318.090 4986.555 3318.260 4987.035 ;
        RECT 3318.930 4986.555 3319.100 4987.035 ;
        RECT 3319.770 4986.555 3319.940 4987.035 ;
        RECT 3317.250 4986.385 3319.940 4986.555 ;
        RECT 3317.250 4985.845 3317.505 4986.385 ;
        RECT 3317.250 4985.675 3319.940 4985.845 ;
        RECT 3317.250 4984.825 3317.420 4985.675 ;
        RECT 3318.090 4984.825 3318.260 4985.675 ;
        RECT 3318.930 4984.825 3319.100 4985.675 ;
        RECT 3319.770 4984.825 3319.940 4985.675 ;
      LAYER mcon ;
        RECT 3317.335 4985.675 3317.505 4986.525 ;
      LAYER met1 ;
        RECT 3317.295 4985.615 3317.555 4986.585 ;
        RECT 3317.200 4975.395 3317.520 4975.515 ;
        RECT 3306.120 4975.255 3317.520 4975.395 ;
        RECT 3306.120 4975.115 3306.260 4975.255 ;
        RECT 3302.615 4974.975 3306.260 4975.115 ;
      LAYER via ;
        RECT 3317.295 4985.675 3317.555 4986.525 ;
        RECT 3317.230 4975.255 3317.490 4975.515 ;
      LAYER met2 ;
        RECT 3317.265 4985.675 3317.585 4986.525 ;
        RECT 3317.350 4975.545 3317.490 4985.675 ;
        RECT 3317.230 4975.225 3317.490 4975.545 ;
        RECT 3317.350 4972.845 3317.490 4975.225 ;
    END
  END mgmt_io_out_buf[10]
  PIN mgmt_io_out_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3323.230 4986.555 3323.400 4987.035 ;
        RECT 3324.070 4986.555 3324.240 4987.035 ;
        RECT 3324.910 4986.555 3325.080 4987.035 ;
        RECT 3325.750 4986.555 3325.920 4987.035 ;
        RECT 3323.230 4986.385 3325.920 4986.555 ;
        RECT 3323.230 4985.845 3323.485 4986.385 ;
        RECT 3323.230 4985.675 3325.920 4985.845 ;
        RECT 3323.230 4984.825 3323.400 4985.675 ;
        RECT 3324.070 4984.825 3324.240 4985.675 ;
        RECT 3324.910 4984.825 3325.080 4985.675 ;
        RECT 3325.750 4984.825 3325.920 4985.675 ;
      LAYER mcon ;
        RECT 3323.315 4985.675 3323.485 4986.525 ;
      LAYER met1 ;
        RECT 3323.275 4985.615 3323.535 4986.585 ;
        RECT 3323.180 4974.275 3323.500 4974.395 ;
        RECT 3308.350 4974.135 3323.500 4974.275 ;
        RECT 3308.350 4973.995 3308.490 4974.135 ;
        RECT 3304.615 4973.855 3308.490 4973.995 ;
      LAYER via ;
        RECT 3323.275 4985.675 3323.535 4986.525 ;
        RECT 3323.210 4974.135 3323.470 4974.395 ;
      LAYER met2 ;
        RECT 3323.245 4985.675 3323.565 4986.525 ;
        RECT 3323.330 4974.425 3323.470 4985.675 ;
        RECT 3323.210 4974.105 3323.470 4974.425 ;
        RECT 3323.330 4972.845 3323.470 4974.105 ;
    END
  END mgmt_io_out_buf[9]
  PIN mgmt_io_in_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3315.925 4982.925 3317.515 4983.125 ;
      LAYER mcon ;
        RECT 3315.925 4982.955 3317.015 4983.125 ;
      LAYER met1 ;
        RECT 3315.865 4982.905 3317.075 4983.165 ;
        RECT 3316.230 4975.675 3316.550 4975.795 ;
        RECT 3301.615 4975.535 3316.550 4975.675 ;
      LAYER via ;
        RECT 3315.925 4982.905 3317.015 4983.165 ;
        RECT 3316.260 4975.535 3316.520 4975.795 ;
      LAYER met2 ;
        RECT 3315.925 4982.875 3317.015 4983.195 ;
        RECT 3316.380 4975.825 3316.520 4982.875 ;
        RECT 3316.260 4975.505 3316.520 4975.825 ;
        RECT 3316.380 4972.845 3316.520 4975.505 ;
    END
  END mgmt_io_in_unbuf[10]
  PIN mgmt_io_in_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3321.905 4982.925 3323.495 4983.125 ;
      LAYER mcon ;
        RECT 3321.905 4982.955 3322.995 4983.125 ;
      LAYER met1 ;
        RECT 3321.845 4982.905 3323.055 4983.165 ;
        RECT 3322.210 4974.555 3322.530 4974.675 ;
        RECT 3303.615 4974.415 3322.530 4974.555 ;
      LAYER via ;
        RECT 3321.905 4982.905 3322.995 4983.165 ;
        RECT 3322.240 4974.415 3322.500 4974.675 ;
      LAYER met2 ;
        RECT 3321.905 4982.875 3322.995 4983.195 ;
        RECT 3322.360 4974.705 3322.500 4982.875 ;
        RECT 3322.240 4974.385 3322.500 4974.705 ;
        RECT 3322.360 4972.845 3322.500 4974.385 ;
    END
  END mgmt_io_in_unbuf[9]
  PIN mgmt_io_in_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3327.885 4982.925 3329.475 4983.125 ;
      LAYER mcon ;
        RECT 3327.885 4982.955 3328.975 4983.125 ;
      LAYER met1 ;
        RECT 3327.825 4982.905 3329.035 4983.165 ;
        RECT 3328.190 4973.435 3328.510 4973.555 ;
        RECT 3305.615 4973.295 3328.510 4973.435 ;
      LAYER via ;
        RECT 3327.885 4982.905 3328.975 4983.165 ;
        RECT 3328.220 4973.295 3328.480 4973.555 ;
      LAYER met2 ;
        RECT 3327.885 4982.875 3328.975 4983.195 ;
        RECT 3328.340 4973.585 3328.480 4982.875 ;
        RECT 3328.220 4973.265 3328.480 4973.585 ;
        RECT 3328.340 4972.845 3328.480 4973.265 ;
    END
  END mgmt_io_in_unbuf[8]
  PIN mgmt_io_out_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3329.210 4986.555 3329.380 4987.035 ;
        RECT 3330.050 4986.555 3330.220 4987.035 ;
        RECT 3330.890 4986.555 3331.060 4987.035 ;
        RECT 3331.730 4986.555 3331.900 4987.035 ;
        RECT 3329.210 4986.385 3331.900 4986.555 ;
        RECT 3329.210 4985.845 3329.465 4986.385 ;
        RECT 3329.210 4985.675 3331.900 4985.845 ;
        RECT 3329.210 4984.825 3329.380 4985.675 ;
        RECT 3330.050 4984.825 3330.220 4985.675 ;
        RECT 3330.890 4984.825 3331.060 4985.675 ;
        RECT 3331.730 4984.825 3331.900 4985.675 ;
      LAYER mcon ;
        RECT 3329.295 4985.675 3329.465 4986.525 ;
      LAYER met1 ;
        RECT 3329.255 4985.615 3329.515 4986.585 ;
        RECT 3329.160 4973.155 3329.480 4973.275 ;
        RECT 3310.170 4973.015 3329.480 4973.155 ;
        RECT 3310.170 4972.875 3310.310 4973.015 ;
        RECT 3306.615 4972.735 3310.310 4972.875 ;
      LAYER via ;
        RECT 3329.255 4985.675 3329.515 4986.525 ;
        RECT 3329.190 4973.015 3329.450 4973.275 ;
      LAYER met2 ;
        RECT 3329.225 4985.675 3329.545 4986.525 ;
        RECT 3329.310 4973.305 3329.450 4985.675 ;
        RECT 3329.190 4972.985 3329.450 4973.305 ;
        RECT 3329.310 4972.845 3329.450 4972.985 ;
    END
  END mgmt_io_out_buf[8]
  PIN mgmt_io_in_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 3612.780 3381.860 3614.370 ;
      LAYER mcon ;
        RECT 3381.690 3613.280 3381.860 3614.370 ;
      LAYER met1 ;
        RECT 3371.900 3614.065 3372.040 3643.605 ;
        RECT 3371.900 3613.745 3372.160 3614.065 ;
        RECT 3381.640 3613.220 3381.900 3614.430 ;
      LAYER via ;
        RECT 3371.900 3613.775 3372.160 3614.035 ;
        RECT 3381.640 3613.280 3381.900 3614.370 ;
      LAYER met2 ;
        RECT 3371.870 3613.915 3372.190 3614.035 ;
        RECT 3381.610 3613.915 3381.930 3614.370 ;
        RECT 3369.210 3613.775 3381.930 3613.915 ;
        RECT 3381.610 3613.280 3381.930 3613.775 ;
    END
  END mgmt_io_in_unbuf[7]
  PIN mgmt_io_in_unbuf[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 3606.800 3381.860 3608.390 ;
      LAYER mcon ;
        RECT 3381.690 3607.300 3381.860 3608.390 ;
      LAYER met1 ;
        RECT 3370.780 3608.085 3370.920 3641.605 ;
        RECT 3370.780 3607.765 3371.040 3608.085 ;
        RECT 3381.640 3607.240 3381.900 3608.450 ;
      LAYER via ;
        RECT 3370.780 3607.795 3371.040 3608.055 ;
        RECT 3381.640 3607.300 3381.900 3608.390 ;
      LAYER met2 ;
        RECT 3370.750 3607.935 3371.070 3608.055 ;
        RECT 3381.610 3607.935 3381.930 3608.390 ;
        RECT 3370.330 3607.795 3381.930 3607.935 ;
        RECT 3381.610 3607.300 3381.930 3607.795 ;
    END
  END mgmt_io_in_unbuf[6]
  PIN mgmt_io_out_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 3612.875 3385.770 3613.045 ;
        RECT 3384.410 3612.790 3385.290 3612.875 ;
        RECT 3384.410 3612.205 3384.580 3612.790 ;
        RECT 3383.560 3612.035 3384.580 3612.205 ;
        RECT 3384.410 3611.365 3384.580 3612.035 ;
        RECT 3383.560 3611.195 3384.580 3611.365 ;
        RECT 3384.410 3610.525 3384.580 3611.195 ;
        RECT 3383.560 3610.355 3384.580 3610.525 ;
        RECT 3385.120 3612.205 3385.290 3612.790 ;
        RECT 3385.120 3612.035 3385.770 3612.205 ;
        RECT 3385.120 3611.365 3385.290 3612.035 ;
        RECT 3385.120 3611.195 3385.770 3611.365 ;
        RECT 3385.120 3610.525 3385.290 3611.195 ;
        RECT 3385.120 3610.355 3385.770 3610.525 ;
      LAYER met1 ;
        RECT 3371.340 3639.950 3371.480 3642.605 ;
        RECT 3371.340 3639.810 3371.760 3639.950 ;
        RECT 3371.620 3613.095 3371.760 3639.810 ;
        RECT 3371.620 3612.775 3371.880 3613.095 ;
        RECT 3384.350 3612.740 3385.320 3613.000 ;
      LAYER via ;
        RECT 3371.620 3612.805 3371.880 3613.065 ;
        RECT 3384.410 3612.740 3385.260 3613.000 ;
      LAYER met2 ;
        RECT 3371.590 3612.945 3371.910 3613.065 ;
        RECT 3384.410 3612.945 3385.260 3613.030 ;
        RECT 3369.210 3612.805 3385.260 3612.945 ;
        RECT 3384.410 3612.710 3385.260 3612.805 ;
    END
  END mgmt_io_out_buf[7]
  PIN mgmt_io_out_buf[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 3606.895 3385.770 3607.065 ;
        RECT 3384.410 3606.810 3385.290 3606.895 ;
        RECT 3384.410 3606.225 3384.580 3606.810 ;
        RECT 3383.560 3606.055 3384.580 3606.225 ;
        RECT 3384.410 3605.385 3384.580 3606.055 ;
        RECT 3383.560 3605.215 3384.580 3605.385 ;
        RECT 3384.410 3604.545 3384.580 3605.215 ;
        RECT 3383.560 3604.375 3384.580 3604.545 ;
        RECT 3385.120 3606.225 3385.290 3606.810 ;
        RECT 3385.120 3606.055 3385.770 3606.225 ;
        RECT 3385.120 3605.385 3385.290 3606.055 ;
        RECT 3385.120 3605.215 3385.770 3605.385 ;
        RECT 3385.120 3604.545 3385.290 3605.215 ;
        RECT 3385.120 3604.375 3385.770 3604.545 ;
      LAYER met1 ;
        RECT 3370.220 3638.040 3370.360 3640.605 ;
        RECT 3370.220 3637.900 3370.640 3638.040 ;
        RECT 3370.500 3607.115 3370.640 3637.900 ;
        RECT 3370.500 3606.795 3370.760 3607.115 ;
        RECT 3384.350 3606.760 3385.320 3607.020 ;
      LAYER via ;
        RECT 3370.500 3606.825 3370.760 3607.085 ;
        RECT 3384.410 3606.760 3385.260 3607.020 ;
      LAYER met2 ;
        RECT 3370.470 3606.965 3370.790 3607.085 ;
        RECT 3384.410 3606.965 3385.260 3607.050 ;
        RECT 3370.330 3606.825 3385.260 3606.965 ;
        RECT 3384.410 3606.730 3385.260 3606.825 ;
    END
  END mgmt_io_out_buf[6]
  PIN mgmt_io_in_unbuf[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2230.700 3381.860 2232.290 ;
      LAYER mcon ;
        RECT 3381.690 2231.200 3381.860 2232.290 ;
      LAYER met1 ;
        RECT 3369.800 2231.985 3369.940 2281.275 ;
        RECT 3369.800 2231.665 3370.060 2231.985 ;
        RECT 3381.640 2231.140 3381.900 2232.350 ;
      LAYER via ;
        RECT 3369.800 2231.695 3370.060 2231.955 ;
        RECT 3381.640 2231.200 3381.900 2232.290 ;
      LAYER met2 ;
        RECT 3369.770 2231.835 3370.090 2231.955 ;
        RECT 3381.610 2231.835 3381.930 2232.290 ;
        RECT 3365.990 2231.695 3381.930 2231.835 ;
        RECT 3381.610 2231.200 3381.930 2231.695 ;
    END
  END mgmt_io_in_unbuf[5]
  PIN mgmt_io_in_unbuf[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2224.720 3381.860 2226.310 ;
      LAYER mcon ;
        RECT 3381.690 2225.220 3381.860 2226.310 ;
      LAYER met1 ;
        RECT 3368.680 2226.005 3368.820 2279.275 ;
        RECT 3368.680 2225.685 3368.940 2226.005 ;
        RECT 3381.640 2225.160 3381.900 2226.370 ;
      LAYER via ;
        RECT 3368.680 2225.715 3368.940 2225.975 ;
        RECT 3381.640 2225.220 3381.900 2226.310 ;
      LAYER met2 ;
        RECT 3368.650 2225.855 3368.970 2225.975 ;
        RECT 3381.610 2225.855 3381.930 2226.310 ;
        RECT 3365.990 2225.715 3381.930 2225.855 ;
        RECT 3381.610 2225.220 3381.930 2225.715 ;
    END
  END mgmt_io_in_unbuf[4]
  PIN mgmt_io_in_unbuf[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2218.740 3381.860 2220.330 ;
      LAYER mcon ;
        RECT 3381.690 2219.240 3381.860 2220.330 ;
      LAYER met1 ;
        RECT 3367.560 2220.025 3367.700 2277.275 ;
        RECT 3367.560 2219.705 3367.820 2220.025 ;
        RECT 3381.640 2219.180 3381.900 2220.390 ;
      LAYER via ;
        RECT 3367.560 2219.735 3367.820 2219.995 ;
        RECT 3381.640 2219.240 3381.900 2220.330 ;
      LAYER met2 ;
        RECT 3367.530 2219.875 3367.850 2219.995 ;
        RECT 3381.610 2219.875 3381.930 2220.330 ;
        RECT 3365.990 2219.735 3381.930 2219.875 ;
        RECT 3381.610 2219.240 3381.930 2219.735 ;
    END
  END mgmt_io_in_unbuf[3]
  PIN mgmt_io_in_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2212.760 3381.860 2214.350 ;
      LAYER mcon ;
        RECT 3381.690 2213.260 3381.860 2214.350 ;
      LAYER met1 ;
        RECT 3366.440 2214.045 3366.580 2275.275 ;
        RECT 3366.440 2213.725 3366.700 2214.045 ;
        RECT 3381.640 2213.200 3381.900 2214.410 ;
      LAYER via ;
        RECT 3366.440 2213.755 3366.700 2214.015 ;
        RECT 3381.640 2213.260 3381.900 2214.350 ;
      LAYER met2 ;
        RECT 3366.410 2213.895 3366.730 2214.015 ;
        RECT 3381.610 2213.895 3381.930 2214.350 ;
        RECT 3365.990 2213.755 3381.930 2213.895 ;
        RECT 3381.610 2213.260 3381.930 2213.755 ;
    END
  END mgmt_io_in_unbuf[2]
  PIN mgmt_io_in_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2206.780 3381.860 2208.370 ;
      LAYER mcon ;
        RECT 3381.690 2207.280 3381.860 2208.370 ;
      LAYER met1 ;
        RECT 3365.320 2208.065 3365.460 2273.275 ;
        RECT 3365.320 2207.745 3365.580 2208.065 ;
        RECT 3381.640 2207.220 3381.900 2208.430 ;
      LAYER via ;
        RECT 3365.320 2207.775 3365.580 2208.035 ;
        RECT 3381.640 2207.280 3381.900 2208.370 ;
      LAYER met2 ;
        RECT 3365.290 2207.915 3365.610 2208.035 ;
        RECT 3381.610 2207.915 3381.930 2208.370 ;
        RECT 3364.865 2207.775 3381.930 2207.915 ;
        RECT 3381.610 2207.280 3381.930 2207.775 ;
    END
  END mgmt_io_in_unbuf[1]
  PIN mgmt_io_in_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3381.660 2200.800 3381.860 2202.390 ;
      LAYER mcon ;
        RECT 3381.690 2201.300 3381.860 2202.390 ;
      LAYER met1 ;
        RECT 3364.200 2202.085 3364.340 2271.275 ;
        RECT 3364.200 2201.765 3364.460 2202.085 ;
        RECT 3381.640 2201.240 3381.900 2202.450 ;
      LAYER via ;
        RECT 3364.200 2201.795 3364.460 2202.055 ;
        RECT 3381.640 2201.300 3381.900 2202.390 ;
      LAYER met2 ;
        RECT 3364.170 2201.935 3364.490 2202.055 ;
        RECT 3381.610 2201.935 3381.930 2202.390 ;
        RECT 3363.750 2201.795 3381.930 2201.935 ;
        RECT 3381.610 2201.300 3381.930 2201.795 ;
    END
  END mgmt_io_in_unbuf[0]
  PIN mgmt_io_out_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2200.895 3385.770 2201.065 ;
        RECT 3384.410 2200.810 3385.290 2200.895 ;
        RECT 3384.410 2200.225 3384.580 2200.810 ;
        RECT 3383.560 2200.055 3384.580 2200.225 ;
        RECT 3384.410 2199.385 3384.580 2200.055 ;
        RECT 3383.560 2199.215 3384.580 2199.385 ;
        RECT 3384.410 2198.545 3384.580 2199.215 ;
        RECT 3383.560 2198.375 3384.580 2198.545 ;
        RECT 3385.120 2200.225 3385.290 2200.810 ;
        RECT 3385.120 2200.055 3385.770 2200.225 ;
        RECT 3385.120 2199.385 3385.290 2200.055 ;
        RECT 3385.120 2199.215 3385.770 2199.385 ;
        RECT 3385.120 2198.545 3385.290 2199.215 ;
        RECT 3385.120 2198.375 3385.770 2198.545 ;
      LAYER met1 ;
        RECT 3363.640 2266.850 3363.780 2270.275 ;
        RECT 3363.640 2266.710 3364.060 2266.850 ;
        RECT 3363.920 2201.115 3364.060 2266.710 ;
        RECT 3363.920 2200.795 3364.180 2201.115 ;
        RECT 3384.350 2200.760 3385.320 2201.020 ;
      LAYER via ;
        RECT 3363.920 2200.825 3364.180 2201.085 ;
        RECT 3384.410 2200.760 3385.260 2201.020 ;
      LAYER met2 ;
        RECT 3363.890 2200.965 3364.210 2201.085 ;
        RECT 3384.410 2200.965 3385.260 2201.050 ;
        RECT 3363.750 2200.825 3385.260 2200.965 ;
        RECT 3384.410 2200.730 3385.260 2200.825 ;
    END
  END mgmt_io_out_buf[0]
  PIN mgmt_io_out_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2206.875 3385.770 2207.045 ;
        RECT 3384.410 2206.790 3385.290 2206.875 ;
        RECT 3384.410 2206.205 3384.580 2206.790 ;
        RECT 3383.560 2206.035 3384.580 2206.205 ;
        RECT 3384.410 2205.365 3384.580 2206.035 ;
        RECT 3383.560 2205.195 3384.580 2205.365 ;
        RECT 3384.410 2204.525 3384.580 2205.195 ;
        RECT 3383.560 2204.355 3384.580 2204.525 ;
        RECT 3385.120 2206.205 3385.290 2206.790 ;
        RECT 3385.120 2206.035 3385.770 2206.205 ;
        RECT 3385.120 2205.365 3385.290 2206.035 ;
        RECT 3385.120 2205.195 3385.770 2205.365 ;
        RECT 3385.120 2204.525 3385.290 2205.195 ;
        RECT 3385.120 2204.355 3385.770 2204.525 ;
      LAYER met1 ;
        RECT 3364.760 2268.790 3364.900 2272.275 ;
        RECT 3364.760 2268.650 3365.180 2268.790 ;
        RECT 3365.040 2207.095 3365.180 2268.650 ;
        RECT 3365.040 2206.775 3365.300 2207.095 ;
        RECT 3384.350 2206.740 3385.320 2207.000 ;
      LAYER via ;
        RECT 3365.040 2206.805 3365.300 2207.065 ;
        RECT 3384.410 2206.740 3385.260 2207.000 ;
      LAYER met2 ;
        RECT 3365.010 2206.945 3365.330 2207.065 ;
        RECT 3384.410 2206.945 3385.260 2207.030 ;
        RECT 3364.865 2206.805 3385.260 2206.945 ;
        RECT 3384.410 2206.710 3385.260 2206.805 ;
    END
  END mgmt_io_out_buf[1]
  PIN mgmt_io_out_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2212.855 3385.770 2213.025 ;
        RECT 3384.410 2212.770 3385.290 2212.855 ;
        RECT 3384.410 2212.185 3384.580 2212.770 ;
        RECT 3383.560 2212.015 3384.580 2212.185 ;
        RECT 3384.410 2211.345 3384.580 2212.015 ;
        RECT 3383.560 2211.175 3384.580 2211.345 ;
        RECT 3384.410 2210.505 3384.580 2211.175 ;
        RECT 3383.560 2210.335 3384.580 2210.505 ;
        RECT 3385.120 2212.185 3385.290 2212.770 ;
        RECT 3385.120 2212.015 3385.770 2212.185 ;
        RECT 3385.120 2211.345 3385.290 2212.015 ;
        RECT 3385.120 2211.175 3385.770 2211.345 ;
        RECT 3385.120 2210.505 3385.290 2211.175 ;
        RECT 3385.120 2210.335 3385.770 2210.505 ;
      LAYER met1 ;
        RECT 3365.880 2270.900 3366.020 2274.275 ;
        RECT 3365.880 2270.760 3366.300 2270.900 ;
        RECT 3366.160 2213.075 3366.300 2270.760 ;
        RECT 3366.160 2212.755 3366.420 2213.075 ;
        RECT 3384.350 2212.720 3385.320 2212.980 ;
      LAYER via ;
        RECT 3366.160 2212.785 3366.420 2213.045 ;
        RECT 3384.410 2212.720 3385.260 2212.980 ;
      LAYER met2 ;
        RECT 3366.130 2212.925 3366.450 2213.045 ;
        RECT 3384.410 2212.925 3385.260 2213.010 ;
        RECT 3365.990 2212.785 3385.260 2212.925 ;
        RECT 3384.410 2212.690 3385.260 2212.785 ;
    END
  END mgmt_io_out_buf[2]
  PIN mgmt_io_out_buf[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2218.835 3385.770 2219.005 ;
        RECT 3384.410 2218.750 3385.290 2218.835 ;
        RECT 3384.410 2218.165 3384.580 2218.750 ;
        RECT 3383.560 2217.995 3384.580 2218.165 ;
        RECT 3384.410 2217.325 3384.580 2217.995 ;
        RECT 3383.560 2217.155 3384.580 2217.325 ;
        RECT 3384.410 2216.485 3384.580 2217.155 ;
        RECT 3383.560 2216.315 3384.580 2216.485 ;
        RECT 3385.120 2218.165 3385.290 2218.750 ;
        RECT 3385.120 2217.995 3385.770 2218.165 ;
        RECT 3385.120 2217.325 3385.290 2217.995 ;
        RECT 3385.120 2217.155 3385.770 2217.325 ;
        RECT 3385.120 2216.485 3385.290 2217.155 ;
        RECT 3385.120 2216.315 3385.770 2216.485 ;
      LAYER met1 ;
        RECT 3367.000 2273.110 3367.140 2276.275 ;
        RECT 3367.000 2272.970 3367.420 2273.110 ;
        RECT 3367.280 2219.055 3367.420 2272.970 ;
        RECT 3367.280 2218.735 3367.540 2219.055 ;
        RECT 3384.350 2218.700 3385.320 2218.960 ;
      LAYER via ;
        RECT 3367.280 2218.765 3367.540 2219.025 ;
        RECT 3384.410 2218.700 3385.260 2218.960 ;
      LAYER met2 ;
        RECT 3367.250 2218.905 3367.570 2219.025 ;
        RECT 3384.410 2218.905 3385.260 2218.990 ;
        RECT 3365.990 2218.765 3385.260 2218.905 ;
        RECT 3384.410 2218.670 3385.260 2218.765 ;
    END
  END mgmt_io_out_buf[3]
  PIN mgmt_io_out_buf[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2224.815 3385.770 2224.985 ;
        RECT 3384.410 2224.730 3385.290 2224.815 ;
        RECT 3384.410 2224.145 3384.580 2224.730 ;
        RECT 3383.560 2223.975 3384.580 2224.145 ;
        RECT 3384.410 2223.305 3384.580 2223.975 ;
        RECT 3383.560 2223.135 3384.580 2223.305 ;
        RECT 3384.410 2222.465 3384.580 2223.135 ;
        RECT 3383.560 2222.295 3384.580 2222.465 ;
        RECT 3385.120 2224.145 3385.290 2224.730 ;
        RECT 3385.120 2223.975 3385.770 2224.145 ;
        RECT 3385.120 2223.305 3385.290 2223.975 ;
        RECT 3385.120 2223.135 3385.770 2223.305 ;
        RECT 3385.120 2222.465 3385.290 2223.135 ;
        RECT 3385.120 2222.295 3385.770 2222.465 ;
      LAYER met1 ;
        RECT 3368.120 2275.010 3368.260 2278.275 ;
        RECT 3368.120 2274.870 3368.540 2275.010 ;
        RECT 3368.400 2225.035 3368.540 2274.870 ;
        RECT 3368.400 2224.715 3368.660 2225.035 ;
        RECT 3384.350 2224.680 3385.320 2224.940 ;
      LAYER via ;
        RECT 3368.400 2224.745 3368.660 2225.005 ;
        RECT 3384.410 2224.680 3385.260 2224.940 ;
      LAYER met2 ;
        RECT 3368.370 2224.885 3368.690 2225.005 ;
        RECT 3384.410 2224.885 3385.260 2224.970 ;
        RECT 3365.990 2224.745 3385.260 2224.885 ;
        RECT 3384.410 2224.650 3385.260 2224.745 ;
    END
  END mgmt_io_out_buf[4]
  PIN mgmt_io_out_buf[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.560 2230.795 3385.770 2230.965 ;
        RECT 3384.410 2230.710 3385.290 2230.795 ;
        RECT 3384.410 2230.125 3384.580 2230.710 ;
        RECT 3383.560 2229.955 3384.580 2230.125 ;
        RECT 3384.410 2229.285 3384.580 2229.955 ;
        RECT 3383.560 2229.115 3384.580 2229.285 ;
        RECT 3384.410 2228.445 3384.580 2229.115 ;
        RECT 3383.560 2228.275 3384.580 2228.445 ;
        RECT 3385.120 2230.125 3385.290 2230.710 ;
        RECT 3385.120 2229.955 3385.770 2230.125 ;
        RECT 3385.120 2229.285 3385.290 2229.955 ;
        RECT 3385.120 2229.115 3385.770 2229.285 ;
        RECT 3385.120 2228.445 3385.290 2229.115 ;
        RECT 3385.120 2228.275 3385.770 2228.445 ;
      LAYER met1 ;
        RECT 3369.240 2276.890 3369.380 2280.275 ;
        RECT 3369.240 2276.750 3369.660 2276.890 ;
        RECT 3369.520 2231.015 3369.660 2276.750 ;
        RECT 3369.520 2230.695 3369.780 2231.015 ;
        RECT 3384.350 2230.660 3385.320 2230.920 ;
      LAYER via ;
        RECT 3369.520 2230.725 3369.780 2230.985 ;
        RECT 3384.410 2230.660 3385.260 2230.920 ;
      LAYER met2 ;
        RECT 3369.490 2230.865 3369.810 2230.985 ;
        RECT 3384.410 2230.865 3385.260 2230.950 ;
        RECT 3365.990 2230.725 3385.260 2230.865 ;
        RECT 3384.410 2230.630 3385.260 2230.725 ;
    END
  END mgmt_io_out_buf[5]
  PIN mgmt_io_out_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2196.660 3384.950 2197.760 ;
      LAYER mcon ;
        RECT 3384.750 2196.670 3384.920 2197.760 ;
      LAYER met1 ;
        RECT 3363.940 2196.930 3364.200 2197.250 ;
        RECT 3364.060 1194.240 3364.200 2196.930 ;
        RECT 3384.700 2196.610 3384.960 2197.820 ;
        RECT 3363.780 1194.100 3364.200 1194.240 ;
        RECT 3363.780 1190.250 3363.920 1194.100 ;
      LAYER via ;
        RECT 3363.940 2196.960 3364.200 2197.220 ;
        RECT 3384.700 2196.670 3384.960 2197.760 ;
      LAYER met2 ;
        RECT 3363.910 2197.100 3364.230 2197.220 ;
        RECT 3384.670 2197.100 3384.990 2197.760 ;
        RECT 3363.750 2196.960 3384.990 2197.100 ;
        RECT 3384.670 2196.670 3384.990 2196.960 ;
    END
  END mgmt_io_out_unbuf[0]
  PIN mgmt_io_out_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2202.640 3384.950 2203.740 ;
      LAYER mcon ;
        RECT 3384.750 2202.650 3384.920 2203.740 ;
      LAYER met1 ;
        RECT 3365.060 2202.910 3365.320 2203.230 ;
        RECT 3365.180 1191.800 3365.320 2202.910 ;
        RECT 3384.700 2202.590 3384.960 2203.800 ;
        RECT 3364.900 1191.660 3365.320 1191.800 ;
        RECT 3364.900 1188.250 3365.040 1191.660 ;
      LAYER via ;
        RECT 3365.060 2202.940 3365.320 2203.200 ;
        RECT 3384.700 2202.650 3384.960 2203.740 ;
      LAYER met2 ;
        RECT 3365.030 2203.080 3365.350 2203.200 ;
        RECT 3384.670 2203.080 3384.990 2203.740 ;
        RECT 3364.900 2202.940 3384.990 2203.080 ;
        RECT 3384.670 2202.650 3384.990 2202.940 ;
    END
  END mgmt_io_out_unbuf[1]
  PIN mgmt_io_out_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2208.620 3384.950 2209.720 ;
      LAYER mcon ;
        RECT 3384.750 2208.630 3384.920 2209.720 ;
      LAYER met1 ;
        RECT 3366.180 2208.890 3366.440 2209.210 ;
        RECT 3366.300 1190.070 3366.440 2208.890 ;
        RECT 3384.700 2208.570 3384.960 2209.780 ;
        RECT 3366.020 1189.930 3366.440 1190.070 ;
        RECT 3366.020 1186.250 3366.160 1189.930 ;
      LAYER via ;
        RECT 3366.180 2208.920 3366.440 2209.180 ;
        RECT 3384.700 2208.630 3384.960 2209.720 ;
      LAYER met2 ;
        RECT 3366.150 2209.060 3366.470 2209.180 ;
        RECT 3384.670 2209.060 3384.990 2209.720 ;
        RECT 3365.990 2208.920 3384.990 2209.060 ;
        RECT 3384.670 2208.630 3384.990 2208.920 ;
    END
  END mgmt_io_out_unbuf[2]
  PIN mgmt_io_out_unbuf[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2214.600 3384.950 2215.700 ;
      LAYER mcon ;
        RECT 3384.750 2214.610 3384.920 2215.700 ;
      LAYER met1 ;
        RECT 3367.300 2214.870 3367.560 2215.190 ;
        RECT 3367.420 1188.240 3367.560 2214.870 ;
        RECT 3384.700 2214.550 3384.960 2215.760 ;
        RECT 3367.140 1188.100 3367.560 1188.240 ;
        RECT 3367.140 1184.250 3367.280 1188.100 ;
      LAYER via ;
        RECT 3367.300 2214.900 3367.560 2215.160 ;
        RECT 3384.700 2214.610 3384.960 2215.700 ;
      LAYER met2 ;
        RECT 3367.270 2215.040 3367.590 2215.160 ;
        RECT 3384.670 2215.040 3384.990 2215.700 ;
        RECT 3365.990 2214.900 3384.990 2215.040 ;
        RECT 3384.670 2214.610 3384.990 2214.900 ;
    END
  END mgmt_io_out_unbuf[3]
  PIN mgmt_io_out_unbuf[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2220.580 3384.950 2221.680 ;
      LAYER mcon ;
        RECT 3384.750 2220.590 3384.920 2221.680 ;
      LAYER met1 ;
        RECT 3368.420 2220.850 3368.680 2221.170 ;
        RECT 3368.540 1186.020 3368.680 2220.850 ;
        RECT 3384.700 2220.530 3384.960 2221.740 ;
        RECT 3368.260 1185.880 3368.680 1186.020 ;
        RECT 3368.260 1182.250 3368.400 1185.880 ;
      LAYER via ;
        RECT 3368.420 2220.880 3368.680 2221.140 ;
        RECT 3384.700 2220.590 3384.960 2221.680 ;
      LAYER met2 ;
        RECT 3368.390 2221.020 3368.710 2221.140 ;
        RECT 3384.670 2221.020 3384.990 2221.680 ;
        RECT 3365.990 2220.880 3384.990 2221.020 ;
        RECT 3384.670 2220.590 3384.990 2220.880 ;
    END
  END mgmt_io_out_unbuf[4]
  PIN mgmt_io_out_unbuf[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2226.560 3384.950 2227.660 ;
      LAYER mcon ;
        RECT 3384.750 2226.570 3384.920 2227.660 ;
      LAYER met1 ;
        RECT 3369.540 2226.830 3369.800 2227.150 ;
        RECT 3369.660 1183.990 3369.800 2226.830 ;
        RECT 3384.700 2226.510 3384.960 2227.720 ;
        RECT 3369.380 1183.850 3369.800 1183.990 ;
        RECT 3369.380 1180.250 3369.520 1183.850 ;
      LAYER via ;
        RECT 3369.540 2226.860 3369.800 2227.120 ;
        RECT 3384.700 2226.570 3384.960 2227.660 ;
      LAYER met2 ;
        RECT 3369.510 2227.000 3369.830 2227.120 ;
        RECT 3384.670 2227.000 3384.990 2227.660 ;
        RECT 3365.990 2226.860 3384.990 2227.000 ;
        RECT 3384.670 2226.570 3384.990 2226.860 ;
    END
  END mgmt_io_out_unbuf[5]
  PIN mgmt_io_out_unbuf[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2232.540 3384.950 2233.640 ;
      LAYER mcon ;
        RECT 3384.750 2232.550 3384.920 2233.640 ;
      LAYER met1 ;
        RECT 3370.660 2232.810 3370.920 2233.130 ;
        RECT 3370.780 1182.000 3370.920 2232.810 ;
        RECT 3384.700 2232.490 3384.960 2233.700 ;
        RECT 3370.500 1181.860 3370.920 1182.000 ;
        RECT 3370.500 1178.250 3370.640 1181.860 ;
      LAYER via ;
        RECT 3370.660 2232.840 3370.920 2233.100 ;
        RECT 3384.700 2232.550 3384.960 2233.640 ;
      LAYER met2 ;
        RECT 3370.630 2232.980 3370.950 2233.100 ;
        RECT 3384.670 2232.980 3384.990 2233.640 ;
        RECT 3365.990 2232.840 3384.990 2232.980 ;
        RECT 3384.670 2232.550 3384.990 2232.840 ;
    END
  END mgmt_io_out_unbuf[6]
  PIN mgmt_io_out_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2238.520 3384.950 2239.620 ;
      LAYER mcon ;
        RECT 3384.750 2238.530 3384.920 2239.620 ;
      LAYER met1 ;
        RECT 3371.780 2238.790 3372.040 2239.110 ;
        RECT 3371.900 1180.110 3372.040 2238.790 ;
        RECT 3384.700 2238.470 3384.960 2239.680 ;
        RECT 3371.620 1179.970 3372.040 1180.110 ;
        RECT 3371.620 1176.250 3371.760 1179.970 ;
      LAYER via ;
        RECT 3371.780 2238.820 3372.040 2239.080 ;
        RECT 3384.700 2238.530 3384.960 2239.620 ;
      LAYER met2 ;
        RECT 3371.750 2238.960 3372.070 2239.080 ;
        RECT 3384.670 2238.960 3384.990 2239.620 ;
        RECT 3365.990 2238.820 3384.990 2238.960 ;
        RECT 3384.670 2238.530 3384.990 2238.820 ;
    END
  END mgmt_io_out_unbuf[7]
  PIN mgmt_io_out_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2244.500 3384.950 2245.600 ;
      LAYER mcon ;
        RECT 3384.750 2244.510 3384.920 2245.600 ;
      LAYER met1 ;
        RECT 3372.900 2244.770 3373.160 2245.090 ;
        RECT 3373.020 1178.200 3373.160 2244.770 ;
        RECT 3384.700 2244.450 3384.960 2245.660 ;
        RECT 3372.740 1178.060 3373.160 1178.200 ;
        RECT 3372.740 1174.250 3372.880 1178.060 ;
      LAYER via ;
        RECT 3372.900 2244.800 3373.160 2245.060 ;
        RECT 3384.700 2244.510 3384.960 2245.600 ;
      LAYER met2 ;
        RECT 3372.870 2244.940 3373.190 2245.060 ;
        RECT 3384.670 2244.940 3384.990 2245.600 ;
        RECT 3365.990 2244.800 3384.990 2244.940 ;
        RECT 3384.670 2244.510 3384.990 2244.800 ;
    END
  END mgmt_io_out_unbuf[8]
  PIN mgmt_io_out_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2250.480 3384.950 2251.580 ;
      LAYER mcon ;
        RECT 3384.750 2250.490 3384.920 2251.580 ;
      LAYER met1 ;
        RECT 3374.020 2250.750 3374.280 2251.070 ;
        RECT 3374.140 1176.270 3374.280 2250.750 ;
        RECT 3384.700 2250.430 3384.960 2251.640 ;
        RECT 3373.860 1176.130 3374.280 1176.270 ;
        RECT 3373.860 1172.250 3374.000 1176.130 ;
      LAYER via ;
        RECT 3374.020 2250.780 3374.280 2251.040 ;
        RECT 3384.700 2250.490 3384.960 2251.580 ;
      LAYER met2 ;
        RECT 3373.990 2250.920 3374.310 2251.040 ;
        RECT 3384.670 2250.920 3384.990 2251.580 ;
        RECT 3365.990 2250.780 3384.990 2250.920 ;
        RECT 3384.670 2250.490 3384.990 2250.780 ;
    END
  END mgmt_io_out_unbuf[9]
  PIN mgmt_io_out_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2256.460 3384.950 2257.560 ;
      LAYER mcon ;
        RECT 3384.750 2256.470 3384.920 2257.560 ;
      LAYER met1 ;
        RECT 3375.140 2256.730 3375.400 2257.050 ;
        RECT 3375.260 1174.180 3375.400 2256.730 ;
        RECT 3384.700 2256.410 3384.960 2257.620 ;
        RECT 3374.980 1174.040 3375.400 1174.180 ;
        RECT 3374.980 1170.250 3375.120 1174.040 ;
      LAYER via ;
        RECT 3375.140 2256.760 3375.400 2257.020 ;
        RECT 3384.700 2256.470 3384.960 2257.560 ;
      LAYER met2 ;
        RECT 3375.110 2256.900 3375.430 2257.020 ;
        RECT 3384.670 2256.900 3384.990 2257.560 ;
        RECT 3365.990 2256.760 3384.990 2256.900 ;
        RECT 3384.670 2256.470 3384.990 2256.760 ;
    END
  END mgmt_io_out_unbuf[10]
  PIN mgmt_io_out_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.750 2262.440 3384.950 2263.540 ;
      LAYER mcon ;
        RECT 3384.750 2262.450 3384.920 2263.540 ;
      LAYER met1 ;
        RECT 3376.400 2262.710 3376.660 2263.030 ;
        RECT 3376.520 1172.180 3376.660 2262.710 ;
        RECT 3384.700 2262.390 3384.960 2263.600 ;
        RECT 3376.240 1172.040 3376.660 1172.180 ;
        RECT 3376.240 1168.250 3376.380 1172.040 ;
      LAYER via ;
        RECT 3376.400 2262.740 3376.660 2263.000 ;
        RECT 3384.700 2262.450 3384.960 2263.540 ;
      LAYER met2 ;
        RECT 3376.370 2262.880 3376.690 2263.000 ;
        RECT 3384.670 2262.880 3384.990 2263.540 ;
        RECT 3376.040 2262.740 3384.990 2262.880 ;
        RECT 3384.670 2262.450 3384.990 2262.740 ;
    END
  END mgmt_io_out_unbuf[11]
  PIN mgmt_io_in_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2265.795 3381.490 2265.965 ;
        RECT 3381.320 2265.125 3381.490 2265.795 ;
        RECT 3380.840 2264.955 3381.490 2265.125 ;
        RECT 3381.320 2264.285 3381.490 2264.955 ;
        RECT 3380.840 2264.115 3381.490 2264.285 ;
        RECT 3381.320 2263.530 3381.490 2264.115 ;
        RECT 3382.030 2265.795 3383.050 2265.965 ;
        RECT 3382.030 2265.125 3382.200 2265.795 ;
        RECT 3382.030 2264.955 3383.050 2265.125 ;
        RECT 3382.030 2264.285 3382.200 2264.955 ;
        RECT 3382.030 2264.115 3383.050 2264.285 ;
        RECT 3382.030 2263.530 3382.200 2264.115 ;
        RECT 3381.320 2263.445 3382.200 2263.530 ;
        RECT 3380.840 2263.275 3383.050 2263.445 ;
      LAYER mcon ;
        RECT 3381.350 2263.360 3382.200 2263.530 ;
      LAYER met1 ;
        RECT 3376.680 2263.330 3376.940 2263.650 ;
        RECT 3376.800 1167.250 3376.940 2263.330 ;
        RECT 3381.290 2263.310 3382.260 2263.570 ;
      LAYER via ;
        RECT 3376.680 2263.360 3376.940 2263.620 ;
        RECT 3381.350 2263.310 3382.200 2263.570 ;
      LAYER met2 ;
        RECT 3376.650 2263.500 3376.970 2263.620 ;
        RECT 3381.350 2263.500 3382.200 2263.600 ;
        RECT 3365.990 2263.360 3382.200 2263.500 ;
        RECT 3381.350 2263.280 3382.200 2263.360 ;
    END
  END mgmt_io_in_buf[11]
  PIN mgmt_io_in_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2259.815 3381.490 2259.985 ;
        RECT 3381.320 2259.145 3381.490 2259.815 ;
        RECT 3380.840 2258.975 3381.490 2259.145 ;
        RECT 3381.320 2258.305 3381.490 2258.975 ;
        RECT 3380.840 2258.135 3381.490 2258.305 ;
        RECT 3381.320 2257.550 3381.490 2258.135 ;
        RECT 3382.030 2259.815 3383.050 2259.985 ;
        RECT 3382.030 2259.145 3382.200 2259.815 ;
        RECT 3382.030 2258.975 3383.050 2259.145 ;
        RECT 3382.030 2258.305 3382.200 2258.975 ;
        RECT 3382.030 2258.135 3383.050 2258.305 ;
        RECT 3382.030 2257.550 3382.200 2258.135 ;
        RECT 3381.320 2257.465 3382.200 2257.550 ;
        RECT 3380.840 2257.295 3383.050 2257.465 ;
      LAYER mcon ;
        RECT 3381.350 2257.380 3382.200 2257.550 ;
      LAYER met1 ;
        RECT 3375.420 2257.350 3375.680 2257.670 ;
        RECT 3375.540 1169.250 3375.680 2257.350 ;
        RECT 3381.290 2257.330 3382.260 2257.590 ;
      LAYER via ;
        RECT 3375.420 2257.380 3375.680 2257.640 ;
        RECT 3381.350 2257.330 3382.200 2257.590 ;
      LAYER met2 ;
        RECT 3375.390 2257.520 3375.710 2257.640 ;
        RECT 3381.350 2257.520 3382.200 2257.620 ;
        RECT 3365.990 2257.380 3382.200 2257.520 ;
        RECT 3381.350 2257.300 3382.200 2257.380 ;
    END
  END mgmt_io_in_buf[10]
  PIN mgmt_io_in_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2253.835 3381.490 2254.005 ;
        RECT 3381.320 2253.165 3381.490 2253.835 ;
        RECT 3380.840 2252.995 3381.490 2253.165 ;
        RECT 3381.320 2252.325 3381.490 2252.995 ;
        RECT 3380.840 2252.155 3381.490 2252.325 ;
        RECT 3381.320 2251.570 3381.490 2252.155 ;
        RECT 3382.030 2253.835 3383.050 2254.005 ;
        RECT 3382.030 2253.165 3382.200 2253.835 ;
        RECT 3382.030 2252.995 3383.050 2253.165 ;
        RECT 3382.030 2252.325 3382.200 2252.995 ;
        RECT 3382.030 2252.155 3383.050 2252.325 ;
        RECT 3382.030 2251.570 3382.200 2252.155 ;
        RECT 3381.320 2251.485 3382.200 2251.570 ;
        RECT 3380.840 2251.315 3383.050 2251.485 ;
      LAYER mcon ;
        RECT 3381.350 2251.400 3382.200 2251.570 ;
      LAYER met1 ;
        RECT 3374.300 2251.370 3374.560 2251.690 ;
        RECT 3374.420 1171.250 3374.560 2251.370 ;
        RECT 3381.290 2251.350 3382.260 2251.610 ;
      LAYER via ;
        RECT 3374.300 2251.400 3374.560 2251.660 ;
        RECT 3381.350 2251.350 3382.200 2251.610 ;
      LAYER met2 ;
        RECT 3374.270 2251.540 3374.590 2251.660 ;
        RECT 3381.350 2251.540 3382.200 2251.640 ;
        RECT 3365.990 2251.400 3382.200 2251.540 ;
        RECT 3381.350 2251.320 3382.200 2251.400 ;
    END
  END mgmt_io_in_buf[9]
  PIN mgmt_io_in_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2247.855 3381.490 2248.025 ;
        RECT 3381.320 2247.185 3381.490 2247.855 ;
        RECT 3380.840 2247.015 3381.490 2247.185 ;
        RECT 3381.320 2246.345 3381.490 2247.015 ;
        RECT 3380.840 2246.175 3381.490 2246.345 ;
        RECT 3381.320 2245.590 3381.490 2246.175 ;
        RECT 3382.030 2247.855 3383.050 2248.025 ;
        RECT 3382.030 2247.185 3382.200 2247.855 ;
        RECT 3382.030 2247.015 3383.050 2247.185 ;
        RECT 3382.030 2246.345 3382.200 2247.015 ;
        RECT 3382.030 2246.175 3383.050 2246.345 ;
        RECT 3382.030 2245.590 3382.200 2246.175 ;
        RECT 3381.320 2245.505 3382.200 2245.590 ;
        RECT 3380.840 2245.335 3383.050 2245.505 ;
      LAYER mcon ;
        RECT 3381.350 2245.420 3382.200 2245.590 ;
      LAYER met1 ;
        RECT 3373.180 2245.390 3373.440 2245.710 ;
        RECT 3373.300 1173.250 3373.440 2245.390 ;
        RECT 3381.290 2245.370 3382.260 2245.630 ;
      LAYER via ;
        RECT 3373.180 2245.420 3373.440 2245.680 ;
        RECT 3381.350 2245.370 3382.200 2245.630 ;
      LAYER met2 ;
        RECT 3373.150 2245.560 3373.470 2245.680 ;
        RECT 3381.350 2245.560 3382.200 2245.660 ;
        RECT 3365.990 2245.420 3382.200 2245.560 ;
        RECT 3381.350 2245.340 3382.200 2245.420 ;
    END
  END mgmt_io_in_buf[8]
  PIN mgmt_io_in_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2241.875 3381.490 2242.045 ;
        RECT 3381.320 2241.205 3381.490 2241.875 ;
        RECT 3380.840 2241.035 3381.490 2241.205 ;
        RECT 3381.320 2240.365 3381.490 2241.035 ;
        RECT 3380.840 2240.195 3381.490 2240.365 ;
        RECT 3381.320 2239.610 3381.490 2240.195 ;
        RECT 3382.030 2241.875 3383.050 2242.045 ;
        RECT 3382.030 2241.205 3382.200 2241.875 ;
        RECT 3382.030 2241.035 3383.050 2241.205 ;
        RECT 3382.030 2240.365 3382.200 2241.035 ;
        RECT 3382.030 2240.195 3383.050 2240.365 ;
        RECT 3382.030 2239.610 3382.200 2240.195 ;
        RECT 3381.320 2239.525 3382.200 2239.610 ;
        RECT 3380.840 2239.355 3383.050 2239.525 ;
      LAYER mcon ;
        RECT 3381.350 2239.440 3382.200 2239.610 ;
      LAYER met1 ;
        RECT 3372.060 2239.410 3372.320 2239.730 ;
        RECT 3372.180 1175.250 3372.320 2239.410 ;
        RECT 3381.290 2239.390 3382.260 2239.650 ;
      LAYER via ;
        RECT 3372.060 2239.440 3372.320 2239.700 ;
        RECT 3381.350 2239.390 3382.200 2239.650 ;
      LAYER met2 ;
        RECT 3372.030 2239.580 3372.350 2239.700 ;
        RECT 3381.350 2239.580 3382.200 2239.680 ;
        RECT 3365.990 2239.440 3382.200 2239.580 ;
        RECT 3381.350 2239.360 3382.200 2239.440 ;
    END
  END mgmt_io_in_buf[7]
  PIN mgmt_io_in_buf[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2235.895 3381.490 2236.065 ;
        RECT 3381.320 2235.225 3381.490 2235.895 ;
        RECT 3380.840 2235.055 3381.490 2235.225 ;
        RECT 3381.320 2234.385 3381.490 2235.055 ;
        RECT 3380.840 2234.215 3381.490 2234.385 ;
        RECT 3381.320 2233.630 3381.490 2234.215 ;
        RECT 3382.030 2235.895 3383.050 2236.065 ;
        RECT 3382.030 2235.225 3382.200 2235.895 ;
        RECT 3382.030 2235.055 3383.050 2235.225 ;
        RECT 3382.030 2234.385 3382.200 2235.055 ;
        RECT 3382.030 2234.215 3383.050 2234.385 ;
        RECT 3382.030 2233.630 3382.200 2234.215 ;
        RECT 3381.320 2233.545 3382.200 2233.630 ;
        RECT 3380.840 2233.375 3383.050 2233.545 ;
      LAYER mcon ;
        RECT 3381.350 2233.460 3382.200 2233.630 ;
      LAYER met1 ;
        RECT 3370.940 2233.430 3371.200 2233.750 ;
        RECT 3371.060 1177.250 3371.200 2233.430 ;
        RECT 3381.290 2233.410 3382.260 2233.670 ;
      LAYER via ;
        RECT 3370.940 2233.460 3371.200 2233.720 ;
        RECT 3381.350 2233.410 3382.200 2233.670 ;
      LAYER met2 ;
        RECT 3370.910 2233.600 3371.230 2233.720 ;
        RECT 3381.350 2233.600 3382.200 2233.700 ;
        RECT 3365.990 2233.460 3382.200 2233.600 ;
        RECT 3381.350 2233.380 3382.200 2233.460 ;
    END
  END mgmt_io_in_buf[6]
  PIN mgmt_io_in_buf[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2229.915 3381.490 2230.085 ;
        RECT 3381.320 2229.245 3381.490 2229.915 ;
        RECT 3380.840 2229.075 3381.490 2229.245 ;
        RECT 3381.320 2228.405 3381.490 2229.075 ;
        RECT 3380.840 2228.235 3381.490 2228.405 ;
        RECT 3381.320 2227.650 3381.490 2228.235 ;
        RECT 3382.030 2229.915 3383.050 2230.085 ;
        RECT 3382.030 2229.245 3382.200 2229.915 ;
        RECT 3382.030 2229.075 3383.050 2229.245 ;
        RECT 3382.030 2228.405 3382.200 2229.075 ;
        RECT 3382.030 2228.235 3383.050 2228.405 ;
        RECT 3382.030 2227.650 3382.200 2228.235 ;
        RECT 3381.320 2227.565 3382.200 2227.650 ;
        RECT 3380.840 2227.395 3383.050 2227.565 ;
      LAYER mcon ;
        RECT 3381.350 2227.480 3382.200 2227.650 ;
      LAYER met1 ;
        RECT 3369.820 2227.450 3370.080 2227.770 ;
        RECT 3369.940 1179.250 3370.080 2227.450 ;
        RECT 3381.290 2227.430 3382.260 2227.690 ;
      LAYER via ;
        RECT 3369.820 2227.480 3370.080 2227.740 ;
        RECT 3381.350 2227.430 3382.200 2227.690 ;
      LAYER met2 ;
        RECT 3369.790 2227.620 3370.110 2227.740 ;
        RECT 3381.350 2227.620 3382.200 2227.720 ;
        RECT 3365.990 2227.480 3382.200 2227.620 ;
        RECT 3381.350 2227.400 3382.200 2227.480 ;
    END
  END mgmt_io_in_buf[5]
  PIN mgmt_io_in_buf[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2223.935 3381.490 2224.105 ;
        RECT 3381.320 2223.265 3381.490 2223.935 ;
        RECT 3380.840 2223.095 3381.490 2223.265 ;
        RECT 3381.320 2222.425 3381.490 2223.095 ;
        RECT 3380.840 2222.255 3381.490 2222.425 ;
        RECT 3381.320 2221.670 3381.490 2222.255 ;
        RECT 3382.030 2223.935 3383.050 2224.105 ;
        RECT 3382.030 2223.265 3382.200 2223.935 ;
        RECT 3382.030 2223.095 3383.050 2223.265 ;
        RECT 3382.030 2222.425 3382.200 2223.095 ;
        RECT 3382.030 2222.255 3383.050 2222.425 ;
        RECT 3382.030 2221.670 3382.200 2222.255 ;
        RECT 3381.320 2221.585 3382.200 2221.670 ;
        RECT 3380.840 2221.415 3383.050 2221.585 ;
      LAYER mcon ;
        RECT 3381.350 2221.500 3382.200 2221.670 ;
      LAYER met1 ;
        RECT 3368.700 2221.470 3368.960 2221.790 ;
        RECT 3368.820 1181.250 3368.960 2221.470 ;
        RECT 3381.290 2221.450 3382.260 2221.710 ;
      LAYER via ;
        RECT 3368.700 2221.500 3368.960 2221.760 ;
        RECT 3381.350 2221.450 3382.200 2221.710 ;
      LAYER met2 ;
        RECT 3368.670 2221.640 3368.990 2221.760 ;
        RECT 3381.350 2221.640 3382.200 2221.740 ;
        RECT 3365.990 2221.500 3382.200 2221.640 ;
        RECT 3381.350 2221.420 3382.200 2221.500 ;
    END
  END mgmt_io_in_buf[4]
  PIN mgmt_io_in_buf[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2217.955 3381.490 2218.125 ;
        RECT 3381.320 2217.285 3381.490 2217.955 ;
        RECT 3380.840 2217.115 3381.490 2217.285 ;
        RECT 3381.320 2216.445 3381.490 2217.115 ;
        RECT 3380.840 2216.275 3381.490 2216.445 ;
        RECT 3381.320 2215.690 3381.490 2216.275 ;
        RECT 3382.030 2217.955 3383.050 2218.125 ;
        RECT 3382.030 2217.285 3382.200 2217.955 ;
        RECT 3382.030 2217.115 3383.050 2217.285 ;
        RECT 3382.030 2216.445 3382.200 2217.115 ;
        RECT 3382.030 2216.275 3383.050 2216.445 ;
        RECT 3382.030 2215.690 3382.200 2216.275 ;
        RECT 3381.320 2215.605 3382.200 2215.690 ;
        RECT 3380.840 2215.435 3383.050 2215.605 ;
      LAYER mcon ;
        RECT 3381.350 2215.520 3382.200 2215.690 ;
      LAYER met1 ;
        RECT 3367.580 2215.490 3367.840 2215.810 ;
        RECT 3367.700 1183.250 3367.840 2215.490 ;
        RECT 3381.290 2215.470 3382.260 2215.730 ;
      LAYER via ;
        RECT 3367.580 2215.520 3367.840 2215.780 ;
        RECT 3381.350 2215.470 3382.200 2215.730 ;
      LAYER met2 ;
        RECT 3367.550 2215.660 3367.870 2215.780 ;
        RECT 3381.350 2215.660 3382.200 2215.760 ;
        RECT 3365.990 2215.520 3382.200 2215.660 ;
        RECT 3381.350 2215.440 3382.200 2215.520 ;
    END
  END mgmt_io_in_buf[3]
  PIN mgmt_io_in_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2211.975 3381.490 2212.145 ;
        RECT 3381.320 2211.305 3381.490 2211.975 ;
        RECT 3380.840 2211.135 3381.490 2211.305 ;
        RECT 3381.320 2210.465 3381.490 2211.135 ;
        RECT 3380.840 2210.295 3381.490 2210.465 ;
        RECT 3381.320 2209.710 3381.490 2210.295 ;
        RECT 3382.030 2211.975 3383.050 2212.145 ;
        RECT 3382.030 2211.305 3382.200 2211.975 ;
        RECT 3382.030 2211.135 3383.050 2211.305 ;
        RECT 3382.030 2210.465 3382.200 2211.135 ;
        RECT 3382.030 2210.295 3383.050 2210.465 ;
        RECT 3382.030 2209.710 3382.200 2210.295 ;
        RECT 3381.320 2209.625 3382.200 2209.710 ;
        RECT 3380.840 2209.455 3383.050 2209.625 ;
      LAYER mcon ;
        RECT 3381.350 2209.540 3382.200 2209.710 ;
      LAYER met1 ;
        RECT 3366.460 2209.510 3366.720 2209.830 ;
        RECT 3366.580 1185.250 3366.720 2209.510 ;
        RECT 3381.290 2209.490 3382.260 2209.750 ;
      LAYER via ;
        RECT 3366.460 2209.540 3366.720 2209.800 ;
        RECT 3381.350 2209.490 3382.200 2209.750 ;
      LAYER met2 ;
        RECT 3366.430 2209.680 3366.750 2209.800 ;
        RECT 3381.350 2209.680 3382.200 2209.780 ;
        RECT 3365.990 2209.540 3382.200 2209.680 ;
        RECT 3381.350 2209.460 3382.200 2209.540 ;
    END
  END mgmt_io_in_buf[2]
  PIN mgmt_io_in_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2205.995 3381.490 2206.165 ;
        RECT 3381.320 2205.325 3381.490 2205.995 ;
        RECT 3380.840 2205.155 3381.490 2205.325 ;
        RECT 3381.320 2204.485 3381.490 2205.155 ;
        RECT 3380.840 2204.315 3381.490 2204.485 ;
        RECT 3381.320 2203.730 3381.490 2204.315 ;
        RECT 3382.030 2205.995 3383.050 2206.165 ;
        RECT 3382.030 2205.325 3382.200 2205.995 ;
        RECT 3382.030 2205.155 3383.050 2205.325 ;
        RECT 3382.030 2204.485 3382.200 2205.155 ;
        RECT 3382.030 2204.315 3383.050 2204.485 ;
        RECT 3382.030 2203.730 3382.200 2204.315 ;
        RECT 3381.320 2203.645 3382.200 2203.730 ;
        RECT 3380.840 2203.475 3383.050 2203.645 ;
      LAYER mcon ;
        RECT 3381.350 2203.560 3382.200 2203.730 ;
      LAYER met1 ;
        RECT 3365.340 2203.530 3365.600 2203.850 ;
        RECT 3365.460 1187.250 3365.600 2203.530 ;
        RECT 3381.290 2203.510 3382.260 2203.770 ;
      LAYER via ;
        RECT 3365.340 2203.560 3365.600 2203.820 ;
        RECT 3381.350 2203.510 3382.200 2203.770 ;
      LAYER met2 ;
        RECT 3365.310 2203.700 3365.630 2203.820 ;
        RECT 3381.350 2203.700 3382.200 2203.800 ;
        RECT 3364.900 2203.560 3382.200 2203.700 ;
        RECT 3381.350 2203.480 3382.200 2203.560 ;
    END
  END mgmt_io_in_buf[1]
  PIN mgmt_io_in_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3380.840 2200.015 3381.490 2200.185 ;
        RECT 3381.320 2199.345 3381.490 2200.015 ;
        RECT 3380.840 2199.175 3381.490 2199.345 ;
        RECT 3381.320 2198.505 3381.490 2199.175 ;
        RECT 3380.840 2198.335 3381.490 2198.505 ;
        RECT 3381.320 2197.750 3381.490 2198.335 ;
        RECT 3382.030 2200.015 3383.050 2200.185 ;
        RECT 3382.030 2199.345 3382.200 2200.015 ;
        RECT 3382.030 2199.175 3383.050 2199.345 ;
        RECT 3382.030 2198.505 3382.200 2199.175 ;
        RECT 3382.030 2198.335 3383.050 2198.505 ;
        RECT 3382.030 2197.750 3382.200 2198.335 ;
        RECT 3381.320 2197.665 3382.200 2197.750 ;
        RECT 3380.840 2197.495 3383.050 2197.665 ;
      LAYER mcon ;
        RECT 3381.350 2197.580 3382.200 2197.750 ;
      LAYER met1 ;
        RECT 3364.220 2197.550 3364.480 2197.870 ;
        RECT 3364.340 1189.250 3364.480 2197.550 ;
        RECT 3381.290 2197.530 3382.260 2197.790 ;
      LAYER via ;
        RECT 3364.220 2197.580 3364.480 2197.840 ;
        RECT 3381.350 2197.530 3382.200 2197.790 ;
      LAYER met2 ;
        RECT 3364.190 2197.720 3364.510 2197.840 ;
        RECT 3381.350 2197.720 3382.200 2197.820 ;
        RECT 3363.750 2197.580 3382.200 2197.720 ;
        RECT 3381.350 2197.500 3382.200 2197.580 ;
    END
  END mgmt_io_in_buf[0]
  PIN mgmt_io_in_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 851.350 4981.710 852.940 4981.910 ;
      LAYER mcon ;
        RECT 851.850 4981.740 852.940 4981.910 ;
      LAYER met1 ;
        RECT 851.790 4981.690 853.000 4981.950 ;
        RECT 852.315 4977.145 852.635 4977.265 ;
        RECT 852.315 4977.005 860.545 4977.145 ;
      LAYER via ;
        RECT 851.850 4981.690 852.940 4981.950 ;
        RECT 852.345 4977.005 852.605 4977.265 ;
      LAYER met2 ;
        RECT 851.850 4981.660 852.940 4981.980 ;
        RECT 852.345 4977.295 852.485 4981.660 ;
        RECT 852.345 4976.975 852.605 4977.295 ;
        RECT 852.345 4975.490 852.485 4976.975 ;
    END
  END mgmt_io_in_unbuf[12]
  PIN mgmt_io_in_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 845.370 4981.710 846.960 4981.910 ;
      LAYER mcon ;
        RECT 845.870 4981.740 846.960 4981.910 ;
      LAYER met1 ;
        RECT 845.810 4981.690 847.020 4981.950 ;
        RECT 846.215 4976.025 846.535 4976.145 ;
        RECT 846.215 4975.885 858.555 4976.025 ;
      LAYER via ;
        RECT 845.870 4981.690 846.960 4981.950 ;
        RECT 846.245 4975.885 846.505 4976.145 ;
      LAYER met2 ;
        RECT 845.870 4981.660 846.960 4981.980 ;
        RECT 846.365 4976.175 846.505 4981.660 ;
        RECT 846.245 4975.855 846.505 4976.175 ;
        RECT 846.365 4975.275 846.505 4975.855 ;
    END
  END mgmt_io_in_unbuf[13]
  PIN mgmt_io_in_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 839.390 4981.710 840.980 4981.910 ;
      LAYER mcon ;
        RECT 839.890 4981.740 840.980 4981.910 ;
      LAYER met1 ;
        RECT 839.830 4981.690 841.040 4981.950 ;
        RECT 840.355 4974.905 840.675 4975.025 ;
        RECT 840.355 4974.765 856.550 4974.905 ;
      LAYER via ;
        RECT 839.890 4981.690 840.980 4981.950 ;
        RECT 840.385 4974.765 840.645 4975.025 ;
      LAYER met2 ;
        RECT 839.890 4981.660 840.980 4981.980 ;
        RECT 840.385 4975.055 840.525 4981.660 ;
        RECT 840.385 4974.735 840.645 4975.055 ;
        RECT 840.385 4974.400 840.525 4974.735 ;
    END
  END mgmt_io_in_unbuf[14]
  PIN mgmt_io_out_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 836.965 4985.340 837.135 4985.820 ;
        RECT 837.805 4985.340 837.975 4985.820 ;
        RECT 838.645 4985.340 838.815 4985.820 ;
        RECT 839.485 4985.340 839.655 4985.820 ;
        RECT 836.965 4985.170 839.655 4985.340 ;
        RECT 839.400 4984.630 839.655 4985.170 ;
        RECT 836.965 4984.460 839.655 4984.630 ;
        RECT 836.965 4983.610 837.135 4984.460 ;
        RECT 837.805 4983.610 837.975 4984.460 ;
        RECT 838.645 4983.610 838.815 4984.460 ;
        RECT 839.485 4983.610 839.655 4984.460 ;
      LAYER mcon ;
        RECT 839.400 4984.460 839.570 4985.310 ;
      LAYER met1 ;
        RECT 839.350 4984.400 839.610 4985.370 ;
        RECT 839.385 4974.625 839.705 4974.745 ;
        RECT 839.385 4974.485 852.205 4974.625 ;
        RECT 852.065 4974.345 852.205 4974.485 ;
        RECT 852.065 4974.205 855.550 4974.345 ;
      LAYER via ;
        RECT 839.350 4984.460 839.610 4985.310 ;
        RECT 839.415 4974.485 839.675 4974.745 ;
      LAYER met2 ;
        RECT 839.320 4984.460 839.640 4985.310 ;
        RECT 839.415 4974.775 839.555 4984.460 ;
        RECT 839.415 4974.455 839.675 4974.775 ;
        RECT 839.415 4974.400 839.555 4974.455 ;
    END
  END mgmt_io_out_buf[14]
  PIN mgmt_io_out_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 842.945 4985.340 843.115 4985.820 ;
        RECT 843.785 4985.340 843.955 4985.820 ;
        RECT 844.625 4985.340 844.795 4985.820 ;
        RECT 845.465 4985.340 845.635 4985.820 ;
        RECT 842.945 4985.170 845.635 4985.340 ;
        RECT 845.380 4984.630 845.635 4985.170 ;
        RECT 842.945 4984.460 845.635 4984.630 ;
        RECT 842.945 4983.610 843.115 4984.460 ;
        RECT 843.785 4983.610 843.955 4984.460 ;
        RECT 844.625 4983.610 844.795 4984.460 ;
        RECT 845.465 4983.610 845.635 4984.460 ;
      LAYER mcon ;
        RECT 845.380 4984.460 845.550 4985.310 ;
      LAYER met1 ;
        RECT 845.330 4984.400 845.590 4985.370 ;
        RECT 845.365 4975.745 845.685 4975.865 ;
        RECT 845.365 4975.605 854.355 4975.745 ;
        RECT 854.215 4975.465 854.355 4975.605 ;
        RECT 854.215 4975.325 857.555 4975.465 ;
      LAYER via ;
        RECT 845.330 4984.460 845.590 4985.310 ;
        RECT 845.395 4975.605 845.655 4975.865 ;
      LAYER met2 ;
        RECT 845.300 4984.460 845.620 4985.310 ;
        RECT 845.395 4975.895 845.535 4984.460 ;
        RECT 845.395 4975.575 845.655 4975.895 ;
        RECT 845.395 4975.275 845.535 4975.575 ;
    END
  END mgmt_io_out_buf[13]
  PIN mgmt_io_out_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 848.925 4985.340 849.095 4985.820 ;
        RECT 849.765 4985.340 849.935 4985.820 ;
        RECT 850.605 4985.340 850.775 4985.820 ;
        RECT 851.445 4985.340 851.615 4985.820 ;
        RECT 848.925 4985.170 851.615 4985.340 ;
        RECT 851.360 4984.630 851.615 4985.170 ;
        RECT 848.925 4984.460 851.615 4984.630 ;
        RECT 848.925 4983.610 849.095 4984.460 ;
        RECT 849.765 4983.610 849.935 4984.460 ;
        RECT 850.605 4983.610 850.775 4984.460 ;
        RECT 851.445 4983.610 851.615 4984.460 ;
      LAYER mcon ;
        RECT 851.360 4984.460 851.530 4985.310 ;
      LAYER met1 ;
        RECT 851.310 4984.400 851.570 4985.370 ;
        RECT 851.345 4976.585 851.665 4976.705 ;
        RECT 851.345 4976.445 859.545 4976.585 ;
      LAYER via ;
        RECT 851.310 4984.460 851.570 4985.310 ;
        RECT 851.375 4976.445 851.635 4976.705 ;
      LAYER met2 ;
        RECT 851.280 4984.460 851.600 4985.310 ;
        RECT 851.375 4976.735 851.515 4984.460 ;
        RECT 851.375 4976.415 851.635 4976.735 ;
        RECT 851.375 4975.490 851.515 4976.415 ;
    END
  END mgmt_io_out_buf[12]
  PIN mgmt_io_out_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.100 4437.655 204.310 4437.825 ;
        RECT 202.580 4437.570 203.460 4437.655 ;
        RECT 202.580 4436.985 202.750 4437.570 ;
        RECT 202.100 4436.815 202.750 4436.985 ;
        RECT 202.580 4436.145 202.750 4436.815 ;
        RECT 202.100 4435.975 202.750 4436.145 ;
        RECT 202.580 4435.305 202.750 4435.975 ;
        RECT 202.100 4435.135 202.750 4435.305 ;
        RECT 203.290 4436.985 203.460 4437.570 ;
        RECT 203.290 4436.815 204.310 4436.985 ;
        RECT 203.290 4436.145 203.460 4436.815 ;
        RECT 203.290 4435.975 204.310 4436.145 ;
        RECT 203.290 4435.305 203.460 4435.975 ;
        RECT 203.290 4435.135 204.310 4435.305 ;
      LAYER mcon ;
        RECT 202.610 4437.570 203.460 4437.740 ;
      LAYER met1 ;
        RECT 214.815 4437.875 214.955 4461.585 ;
        RECT 202.550 4437.520 203.520 4437.780 ;
        RECT 214.695 4437.555 214.955 4437.875 ;
      LAYER via ;
        RECT 202.610 4437.520 203.460 4437.780 ;
        RECT 214.695 4437.585 214.955 4437.845 ;
      LAYER met2 ;
        RECT 202.610 4437.725 203.460 4437.810 ;
        RECT 214.665 4437.725 214.985 4437.845 ;
        RECT 202.610 4437.585 216.135 4437.725 ;
        RECT 202.610 4437.490 203.460 4437.585 ;
    END
  END mgmt_io_out_buf[15]
  PIN mgmt_io_out_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.100 4431.675 204.310 4431.845 ;
        RECT 202.580 4431.590 203.460 4431.675 ;
        RECT 202.580 4431.005 202.750 4431.590 ;
        RECT 202.100 4430.835 202.750 4431.005 ;
        RECT 202.580 4430.165 202.750 4430.835 ;
        RECT 202.100 4429.995 202.750 4430.165 ;
        RECT 202.580 4429.325 202.750 4429.995 ;
        RECT 202.100 4429.155 202.750 4429.325 ;
        RECT 203.290 4431.005 203.460 4431.590 ;
        RECT 203.290 4430.835 204.310 4431.005 ;
        RECT 203.290 4430.165 203.460 4430.835 ;
        RECT 203.290 4429.995 204.310 4430.165 ;
        RECT 203.290 4429.325 203.460 4429.995 ;
        RECT 203.290 4429.155 204.310 4429.325 ;
      LAYER mcon ;
        RECT 202.610 4431.590 203.460 4431.760 ;
      LAYER met1 ;
        RECT 215.935 4431.895 216.075 4459.585 ;
        RECT 202.550 4431.540 203.520 4431.800 ;
        RECT 215.815 4431.575 216.075 4431.895 ;
      LAYER via ;
        RECT 202.610 4431.540 203.460 4431.800 ;
        RECT 215.815 4431.605 216.075 4431.865 ;
      LAYER met2 ;
        RECT 202.610 4431.745 203.460 4431.830 ;
        RECT 215.785 4431.745 216.105 4431.865 ;
        RECT 202.610 4431.605 216.135 4431.745 ;
        RECT 202.610 4431.510 203.460 4431.605 ;
    END
  END mgmt_io_out_buf[16]
  PIN mgmt_io_in_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.010 4431.580 206.210 4433.170 ;
      LAYER mcon ;
        RECT 206.010 4432.080 206.180 4433.170 ;
      LAYER met1 ;
        RECT 215.375 4458.380 215.515 4460.585 ;
        RECT 215.375 4458.240 215.795 4458.380 ;
        RECT 205.970 4432.020 206.230 4433.230 ;
        RECT 215.655 4432.865 215.795 4458.240 ;
        RECT 215.535 4432.545 215.795 4432.865 ;
      LAYER via ;
        RECT 205.970 4432.080 206.230 4433.170 ;
        RECT 215.535 4432.575 215.795 4432.835 ;
      LAYER met2 ;
        RECT 205.940 4432.715 206.260 4433.170 ;
        RECT 215.505 4432.715 215.825 4432.835 ;
        RECT 205.940 4432.575 216.135 4432.715 ;
        RECT 205.940 4432.080 206.260 4432.575 ;
    END
  END mgmt_io_in_unbuf[16]
  PIN mgmt_io_in_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.010 4437.560 206.210 4439.150 ;
      LAYER mcon ;
        RECT 206.010 4438.060 206.180 4439.150 ;
      LAYER met1 ;
        RECT 214.255 4460.415 214.395 4462.585 ;
        RECT 214.255 4460.275 214.675 4460.415 ;
        RECT 205.970 4438.000 206.230 4439.210 ;
        RECT 214.535 4438.725 214.675 4460.275 ;
        RECT 214.415 4438.405 214.675 4438.725 ;
      LAYER via ;
        RECT 205.970 4438.060 206.230 4439.150 ;
        RECT 214.415 4438.435 214.675 4438.695 ;
      LAYER met2 ;
        RECT 205.940 4438.695 206.260 4439.150 ;
        RECT 205.940 4438.555 216.135 4438.695 ;
        RECT 205.940 4438.060 206.260 4438.555 ;
        RECT 214.385 4438.435 214.705 4438.555 ;
    END
  END mgmt_io_in_unbuf[15]
  PIN mgmt_io_out_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3019.465 204.435 3019.635 ;
        RECT 202.705 3019.380 203.585 3019.465 ;
        RECT 202.705 3018.795 202.875 3019.380 ;
        RECT 202.225 3018.625 202.875 3018.795 ;
        RECT 202.705 3017.955 202.875 3018.625 ;
        RECT 202.225 3017.785 202.875 3017.955 ;
        RECT 202.705 3017.115 202.875 3017.785 ;
        RECT 202.225 3016.945 202.875 3017.115 ;
        RECT 203.415 3018.795 203.585 3019.380 ;
        RECT 203.415 3018.625 204.435 3018.795 ;
        RECT 203.415 3017.955 203.585 3018.625 ;
        RECT 203.415 3017.785 204.435 3017.955 ;
        RECT 203.415 3017.115 203.585 3017.785 ;
        RECT 203.415 3016.945 204.435 3017.115 ;
      LAYER mcon ;
        RECT 202.735 3019.380 203.585 3019.550 ;
      LAYER met1 ;
        RECT 216.915 3019.685 217.055 3063.780 ;
        RECT 202.675 3019.330 203.645 3019.590 ;
        RECT 216.795 3019.365 217.055 3019.685 ;
      LAYER via ;
        RECT 202.735 3019.330 203.585 3019.590 ;
        RECT 216.795 3019.395 217.055 3019.655 ;
      LAYER met2 ;
        RECT 202.735 3019.535 203.585 3019.620 ;
        RECT 216.765 3019.535 217.085 3019.655 ;
        RECT 202.735 3019.395 221.600 3019.535 ;
        RECT 202.735 3019.300 203.585 3019.395 ;
    END
  END mgmt_io_out_buf[17]
  PIN mgmt_io_out_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3013.485 204.435 3013.655 ;
        RECT 202.705 3013.400 203.585 3013.485 ;
        RECT 202.705 3012.815 202.875 3013.400 ;
        RECT 202.225 3012.645 202.875 3012.815 ;
        RECT 202.705 3011.975 202.875 3012.645 ;
        RECT 202.225 3011.805 202.875 3011.975 ;
        RECT 202.705 3011.135 202.875 3011.805 ;
        RECT 202.225 3010.965 202.875 3011.135 ;
        RECT 203.415 3012.815 203.585 3013.400 ;
        RECT 203.415 3012.645 204.435 3012.815 ;
        RECT 203.415 3011.975 203.585 3012.645 ;
        RECT 203.415 3011.805 204.435 3011.975 ;
        RECT 203.415 3011.135 203.585 3011.805 ;
        RECT 203.415 3010.965 204.435 3011.135 ;
      LAYER mcon ;
        RECT 202.735 3013.400 203.585 3013.570 ;
      LAYER met1 ;
        RECT 218.035 3013.705 218.175 3061.780 ;
        RECT 202.675 3013.350 203.645 3013.610 ;
        RECT 217.915 3013.385 218.175 3013.705 ;
      LAYER via ;
        RECT 202.735 3013.350 203.585 3013.610 ;
        RECT 217.915 3013.415 218.175 3013.675 ;
      LAYER met2 ;
        RECT 202.735 3013.555 203.585 3013.640 ;
        RECT 217.885 3013.555 218.205 3013.675 ;
        RECT 202.735 3013.415 221.600 3013.555 ;
        RECT 202.735 3013.320 203.585 3013.415 ;
    END
  END mgmt_io_out_buf[18]
  PIN mgmt_io_out_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3007.505 204.435 3007.675 ;
        RECT 202.705 3007.420 203.585 3007.505 ;
        RECT 202.705 3006.835 202.875 3007.420 ;
        RECT 202.225 3006.665 202.875 3006.835 ;
        RECT 202.705 3005.995 202.875 3006.665 ;
        RECT 202.225 3005.825 202.875 3005.995 ;
        RECT 202.705 3005.155 202.875 3005.825 ;
        RECT 202.225 3004.985 202.875 3005.155 ;
        RECT 203.415 3006.835 203.585 3007.420 ;
        RECT 203.415 3006.665 204.435 3006.835 ;
        RECT 203.415 3005.995 203.585 3006.665 ;
        RECT 203.415 3005.825 204.435 3005.995 ;
        RECT 203.415 3005.155 203.585 3005.825 ;
        RECT 203.415 3004.985 204.435 3005.155 ;
      LAYER mcon ;
        RECT 202.735 3007.420 203.585 3007.590 ;
      LAYER met1 ;
        RECT 219.155 3007.725 219.295 3059.780 ;
        RECT 202.675 3007.370 203.645 3007.630 ;
        RECT 219.035 3007.405 219.295 3007.725 ;
      LAYER via ;
        RECT 202.735 3007.370 203.585 3007.630 ;
        RECT 219.035 3007.435 219.295 3007.695 ;
      LAYER met2 ;
        RECT 202.735 3007.575 203.585 3007.660 ;
        RECT 219.005 3007.575 219.325 3007.695 ;
        RECT 202.735 3007.435 221.600 3007.575 ;
        RECT 202.735 3007.340 203.585 3007.435 ;
    END
  END mgmt_io_out_buf[19]
  PIN mgmt_io_out_buf[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 3001.525 204.435 3001.695 ;
        RECT 202.705 3001.440 203.585 3001.525 ;
        RECT 202.705 3000.855 202.875 3001.440 ;
        RECT 202.225 3000.685 202.875 3000.855 ;
        RECT 202.705 3000.015 202.875 3000.685 ;
        RECT 202.225 2999.845 202.875 3000.015 ;
        RECT 202.705 2999.175 202.875 2999.845 ;
        RECT 202.225 2999.005 202.875 2999.175 ;
        RECT 203.415 3000.855 203.585 3001.440 ;
        RECT 203.415 3000.685 204.435 3000.855 ;
        RECT 203.415 3000.015 203.585 3000.685 ;
        RECT 203.415 2999.845 204.435 3000.015 ;
        RECT 203.415 2999.175 203.585 2999.845 ;
        RECT 203.415 2999.005 204.435 2999.175 ;
      LAYER mcon ;
        RECT 202.735 3001.440 203.585 3001.610 ;
      LAYER met1 ;
        RECT 220.275 3001.745 220.415 3057.780 ;
        RECT 202.675 3001.390 203.645 3001.650 ;
        RECT 220.155 3001.425 220.415 3001.745 ;
      LAYER via ;
        RECT 202.735 3001.390 203.585 3001.650 ;
        RECT 220.155 3001.455 220.415 3001.715 ;
      LAYER met2 ;
        RECT 202.735 3001.595 203.585 3001.680 ;
        RECT 220.125 3001.595 220.445 3001.715 ;
        RECT 202.735 3001.455 221.600 3001.595 ;
        RECT 202.735 3001.360 203.585 3001.455 ;
    END
  END mgmt_io_out_buf[20]
  PIN mgmt_io_out_buf[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 2995.545 204.435 2995.715 ;
        RECT 202.705 2995.460 203.585 2995.545 ;
        RECT 202.705 2994.875 202.875 2995.460 ;
        RECT 202.225 2994.705 202.875 2994.875 ;
        RECT 202.705 2994.035 202.875 2994.705 ;
        RECT 202.225 2993.865 202.875 2994.035 ;
        RECT 202.705 2993.195 202.875 2993.865 ;
        RECT 202.225 2993.025 202.875 2993.195 ;
        RECT 203.415 2994.875 203.585 2995.460 ;
        RECT 203.415 2994.705 204.435 2994.875 ;
        RECT 203.415 2994.035 203.585 2994.705 ;
        RECT 203.415 2993.865 204.435 2994.035 ;
        RECT 203.415 2993.195 203.585 2993.865 ;
        RECT 203.415 2993.025 204.435 2993.195 ;
      LAYER mcon ;
        RECT 202.735 2995.460 203.585 2995.630 ;
      LAYER met1 ;
        RECT 221.395 2995.765 221.535 3055.780 ;
        RECT 202.675 2995.410 203.645 2995.670 ;
        RECT 221.275 2995.445 221.535 2995.765 ;
      LAYER via ;
        RECT 202.735 2995.410 203.585 2995.670 ;
        RECT 221.275 2995.475 221.535 2995.735 ;
      LAYER met2 ;
        RECT 202.735 2995.615 203.585 2995.700 ;
        RECT 221.245 2995.615 221.565 2995.735 ;
        RECT 202.735 2995.475 221.605 2995.615 ;
        RECT 202.735 2995.380 203.585 2995.475 ;
    END
  END mgmt_io_out_buf[21]
  PIN mgmt_io_out_buf[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.225 2989.565 204.435 2989.735 ;
        RECT 202.705 2989.480 203.585 2989.565 ;
        RECT 202.705 2988.895 202.875 2989.480 ;
        RECT 202.225 2988.725 202.875 2988.895 ;
        RECT 202.705 2988.055 202.875 2988.725 ;
        RECT 202.225 2987.885 202.875 2988.055 ;
        RECT 202.705 2987.215 202.875 2987.885 ;
        RECT 202.225 2987.045 202.875 2987.215 ;
        RECT 203.415 2988.895 203.585 2989.480 ;
        RECT 203.415 2988.725 204.435 2988.895 ;
        RECT 203.415 2988.055 203.585 2988.725 ;
        RECT 203.415 2987.885 204.435 2988.055 ;
        RECT 203.415 2987.215 203.585 2987.885 ;
        RECT 203.415 2987.045 204.435 2987.215 ;
      LAYER mcon ;
        RECT 202.735 2989.480 203.585 2989.650 ;
      LAYER met1 ;
        RECT 222.515 2989.785 222.655 3053.780 ;
        RECT 202.675 2989.430 203.645 2989.690 ;
        RECT 222.395 2989.465 222.655 2989.785 ;
      LAYER via ;
        RECT 202.735 2989.430 203.585 2989.690 ;
        RECT 222.395 2989.495 222.655 2989.755 ;
      LAYER met2 ;
        RECT 202.735 2989.635 203.585 2989.720 ;
        RECT 222.365 2989.635 222.685 2989.755 ;
        RECT 202.735 2989.495 222.720 2989.635 ;
        RECT 202.735 2989.400 203.585 2989.495 ;
    END
  END mgmt_io_out_buf[22]
  PIN mgmt_io_in_unbuf[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 2989.470 206.335 2991.060 ;
      LAYER mcon ;
        RECT 206.135 2989.970 206.305 2991.060 ;
      LAYER met1 ;
        RECT 221.955 3051.605 222.095 3054.780 ;
        RECT 221.955 3051.465 222.375 3051.605 ;
        RECT 206.095 2989.910 206.355 2991.120 ;
        RECT 222.235 2990.755 222.375 3051.465 ;
        RECT 222.115 2990.435 222.375 2990.755 ;
      LAYER via ;
        RECT 206.095 2989.970 206.355 2991.060 ;
        RECT 222.115 2990.465 222.375 2990.725 ;
      LAYER met2 ;
        RECT 206.065 2990.605 206.385 2991.060 ;
        RECT 222.085 2990.605 222.405 2990.725 ;
        RECT 206.065 2990.465 222.720 2990.605 ;
        RECT 206.065 2989.970 206.385 2990.465 ;
    END
  END mgmt_io_in_unbuf[22]
  PIN mgmt_io_in_unbuf[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 2995.450 206.335 2997.040 ;
      LAYER mcon ;
        RECT 206.135 2995.950 206.305 2997.040 ;
      LAYER met1 ;
        RECT 220.835 3053.795 220.975 3056.780 ;
        RECT 220.835 3053.655 221.255 3053.795 ;
        RECT 206.095 2995.890 206.355 2997.100 ;
        RECT 221.115 2996.735 221.255 3053.655 ;
        RECT 220.995 2996.415 221.255 2996.735 ;
      LAYER via ;
        RECT 206.095 2995.950 206.355 2997.040 ;
        RECT 220.995 2996.445 221.255 2996.705 ;
      LAYER met2 ;
        RECT 206.065 2996.585 206.385 2997.040 ;
        RECT 220.965 2996.585 221.285 2996.705 ;
        RECT 206.065 2996.445 221.605 2996.585 ;
        RECT 206.065 2995.950 206.385 2996.445 ;
    END
  END mgmt_io_in_unbuf[21]
  PIN mgmt_io_in_unbuf[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3001.430 206.335 3003.020 ;
      LAYER mcon ;
        RECT 206.135 3001.930 206.305 3003.020 ;
      LAYER met1 ;
        RECT 219.715 3055.785 219.855 3058.780 ;
        RECT 219.715 3055.645 220.135 3055.785 ;
        RECT 206.095 3001.870 206.355 3003.080 ;
        RECT 219.995 3002.715 220.135 3055.645 ;
        RECT 219.875 3002.395 220.135 3002.715 ;
      LAYER via ;
        RECT 206.095 3001.930 206.355 3003.020 ;
        RECT 219.875 3002.425 220.135 3002.685 ;
      LAYER met2 ;
        RECT 206.065 3002.565 206.385 3003.020 ;
        RECT 219.845 3002.565 220.165 3002.685 ;
        RECT 206.065 3002.425 221.600 3002.565 ;
        RECT 206.065 3001.930 206.385 3002.425 ;
    END
  END mgmt_io_in_unbuf[20]
  PIN mgmt_io_in_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3007.410 206.335 3009.000 ;
      LAYER mcon ;
        RECT 206.135 3007.910 206.305 3009.000 ;
      LAYER met1 ;
        RECT 218.595 3057.670 218.735 3060.780 ;
        RECT 218.595 3057.530 219.015 3057.670 ;
        RECT 206.095 3007.850 206.355 3009.060 ;
        RECT 218.875 3008.695 219.015 3057.530 ;
        RECT 218.755 3008.375 219.015 3008.695 ;
      LAYER via ;
        RECT 206.095 3007.910 206.355 3009.000 ;
        RECT 218.755 3008.405 219.015 3008.665 ;
      LAYER met2 ;
        RECT 206.065 3008.545 206.385 3009.000 ;
        RECT 218.725 3008.545 219.045 3008.665 ;
        RECT 206.065 3008.405 221.600 3008.545 ;
        RECT 206.065 3007.910 206.385 3008.405 ;
    END
  END mgmt_io_in_unbuf[19]
  PIN mgmt_io_in_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3013.390 206.335 3014.980 ;
      LAYER mcon ;
        RECT 206.135 3013.890 206.305 3014.980 ;
      LAYER met1 ;
        RECT 217.475 3059.685 217.615 3062.780 ;
        RECT 217.475 3059.545 217.895 3059.685 ;
        RECT 206.095 3013.830 206.355 3015.040 ;
        RECT 217.755 3014.675 217.895 3059.545 ;
        RECT 217.635 3014.355 217.895 3014.675 ;
      LAYER via ;
        RECT 206.095 3013.890 206.355 3014.980 ;
        RECT 217.635 3014.385 217.895 3014.645 ;
      LAYER met2 ;
        RECT 206.065 3014.525 206.385 3014.980 ;
        RECT 217.605 3014.525 217.925 3014.645 ;
        RECT 206.065 3014.385 221.600 3014.525 ;
        RECT 206.065 3013.890 206.385 3014.385 ;
    END
  END mgmt_io_in_unbuf[18]
  PIN mgmt_io_in_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.135 3019.370 206.335 3020.960 ;
      LAYER mcon ;
        RECT 206.135 3019.870 206.305 3020.960 ;
      LAYER met1 ;
        RECT 216.355 3061.745 216.495 3064.780 ;
        RECT 216.355 3061.605 216.775 3061.745 ;
        RECT 206.095 3019.810 206.355 3021.020 ;
        RECT 216.635 3020.655 216.775 3061.605 ;
        RECT 216.515 3020.335 216.775 3020.655 ;
      LAYER via ;
        RECT 206.095 3019.870 206.355 3020.960 ;
        RECT 216.515 3020.365 216.775 3020.625 ;
      LAYER met2 ;
        RECT 206.065 3020.505 206.385 3020.960 ;
        RECT 216.485 3020.505 216.805 3020.625 ;
        RECT 206.065 3020.365 221.600 3020.505 ;
        RECT 206.065 3019.870 206.385 3020.365 ;
    END
  END mgmt_io_in_unbuf[17]
  PIN mgmt_io_out_buf[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1695.680 204.545 1695.850 ;
        RECT 202.815 1695.595 203.695 1695.680 ;
        RECT 202.815 1695.010 202.985 1695.595 ;
        RECT 202.335 1694.840 202.985 1695.010 ;
        RECT 202.815 1694.170 202.985 1694.840 ;
        RECT 202.335 1694.000 202.985 1694.170 ;
        RECT 202.815 1693.330 202.985 1694.000 ;
        RECT 202.335 1693.160 202.985 1693.330 ;
        RECT 203.525 1695.010 203.695 1695.595 ;
        RECT 203.525 1694.840 204.545 1695.010 ;
        RECT 203.525 1694.170 203.695 1694.840 ;
        RECT 203.525 1694.000 204.545 1694.170 ;
        RECT 203.525 1693.330 203.695 1694.000 ;
        RECT 203.525 1693.160 204.545 1693.330 ;
      LAYER mcon ;
        RECT 202.845 1695.595 203.695 1695.765 ;
      LAYER met1 ;
        RECT 223.495 1695.900 223.635 1772.650 ;
        RECT 202.785 1695.545 203.755 1695.805 ;
        RECT 223.375 1695.580 223.635 1695.900 ;
      LAYER via ;
        RECT 202.845 1695.545 203.695 1695.805 ;
        RECT 223.375 1695.610 223.635 1695.870 ;
      LAYER met2 ;
        RECT 202.845 1695.750 203.695 1695.835 ;
        RECT 223.345 1695.750 223.665 1695.870 ;
        RECT 202.845 1695.610 223.840 1695.750 ;
        RECT 202.845 1695.515 203.695 1695.610 ;
    END
  END mgmt_io_out_buf[23]
  PIN mgmt_io_out_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1689.700 204.545 1689.870 ;
        RECT 202.815 1689.615 203.695 1689.700 ;
        RECT 202.815 1689.030 202.985 1689.615 ;
        RECT 202.335 1688.860 202.985 1689.030 ;
        RECT 202.815 1688.190 202.985 1688.860 ;
        RECT 202.335 1688.020 202.985 1688.190 ;
        RECT 202.815 1687.350 202.985 1688.020 ;
        RECT 202.335 1687.180 202.985 1687.350 ;
        RECT 203.525 1689.030 203.695 1689.615 ;
        RECT 203.525 1688.860 204.545 1689.030 ;
        RECT 203.525 1688.190 203.695 1688.860 ;
        RECT 203.525 1688.020 204.545 1688.190 ;
        RECT 203.525 1687.350 203.695 1688.020 ;
        RECT 203.525 1687.180 204.545 1687.350 ;
      LAYER mcon ;
        RECT 202.845 1689.615 203.695 1689.785 ;
      LAYER met1 ;
        RECT 224.615 1689.920 224.755 1770.650 ;
        RECT 202.785 1689.565 203.755 1689.825 ;
        RECT 224.495 1689.600 224.755 1689.920 ;
      LAYER via ;
        RECT 202.845 1689.565 203.695 1689.825 ;
        RECT 224.495 1689.630 224.755 1689.890 ;
      LAYER met2 ;
        RECT 202.845 1689.770 203.695 1689.855 ;
        RECT 224.465 1689.770 224.785 1689.890 ;
        RECT 202.845 1689.630 224.910 1689.770 ;
        RECT 202.845 1689.535 203.695 1689.630 ;
    END
  END mgmt_io_out_buf[24]
  PIN mgmt_io_out_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1683.720 204.545 1683.890 ;
        RECT 202.815 1683.635 203.695 1683.720 ;
        RECT 202.815 1683.050 202.985 1683.635 ;
        RECT 202.335 1682.880 202.985 1683.050 ;
        RECT 202.815 1682.210 202.985 1682.880 ;
        RECT 202.335 1682.040 202.985 1682.210 ;
        RECT 202.815 1681.370 202.985 1682.040 ;
        RECT 202.335 1681.200 202.985 1681.370 ;
        RECT 203.525 1683.050 203.695 1683.635 ;
        RECT 203.525 1682.880 204.545 1683.050 ;
        RECT 203.525 1682.210 203.695 1682.880 ;
        RECT 203.525 1682.040 204.545 1682.210 ;
        RECT 203.525 1681.370 203.695 1682.040 ;
        RECT 203.525 1681.200 204.545 1681.370 ;
      LAYER mcon ;
        RECT 202.845 1683.635 203.695 1683.805 ;
      LAYER met1 ;
        RECT 225.735 1683.940 225.875 1768.650 ;
        RECT 202.785 1683.585 203.755 1683.845 ;
        RECT 225.615 1683.620 225.875 1683.940 ;
      LAYER via ;
        RECT 202.845 1683.585 203.695 1683.845 ;
        RECT 225.615 1683.650 225.875 1683.910 ;
      LAYER met2 ;
        RECT 202.845 1683.790 203.695 1683.875 ;
        RECT 225.585 1683.790 225.905 1683.910 ;
        RECT 202.845 1683.650 225.975 1683.790 ;
        RECT 202.845 1683.555 203.695 1683.650 ;
    END
  END mgmt_io_out_buf[25]
  PIN mgmt_io_out_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.335 1677.740 204.545 1677.910 ;
        RECT 202.815 1677.655 203.695 1677.740 ;
        RECT 202.815 1677.070 202.985 1677.655 ;
        RECT 202.335 1676.900 202.985 1677.070 ;
        RECT 202.815 1676.230 202.985 1676.900 ;
        RECT 202.335 1676.060 202.985 1676.230 ;
        RECT 202.815 1675.390 202.985 1676.060 ;
        RECT 202.335 1675.220 202.985 1675.390 ;
        RECT 203.525 1677.070 203.695 1677.655 ;
        RECT 203.525 1676.900 204.545 1677.070 ;
        RECT 203.525 1676.230 203.695 1676.900 ;
        RECT 203.525 1676.060 204.545 1676.230 ;
        RECT 203.525 1675.390 203.695 1676.060 ;
        RECT 203.525 1675.220 204.545 1675.390 ;
      LAYER mcon ;
        RECT 202.845 1677.655 203.695 1677.825 ;
      LAYER met1 ;
        RECT 226.855 1677.960 226.995 1766.650 ;
        RECT 202.785 1677.605 203.755 1677.865 ;
        RECT 226.735 1677.640 226.995 1677.960 ;
      LAYER via ;
        RECT 202.845 1677.605 203.695 1677.865 ;
        RECT 226.735 1677.670 226.995 1677.930 ;
      LAYER met2 ;
        RECT 202.845 1677.810 203.695 1677.895 ;
        RECT 226.705 1677.810 227.025 1677.930 ;
        RECT 202.845 1677.670 227.100 1677.810 ;
        RECT 202.845 1677.575 203.695 1677.670 ;
    END
  END mgmt_io_out_buf[26]
  PIN mgmt_io_in_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1677.645 206.445 1679.235 ;
      LAYER mcon ;
        RECT 206.245 1678.145 206.415 1679.235 ;
      LAYER met1 ;
        RECT 226.295 1764.910 226.435 1767.650 ;
        RECT 226.295 1764.770 226.715 1764.910 ;
        RECT 206.205 1678.085 206.465 1679.295 ;
        RECT 226.575 1678.930 226.715 1764.770 ;
        RECT 226.455 1678.610 226.715 1678.930 ;
      LAYER via ;
        RECT 206.205 1678.145 206.465 1679.235 ;
        RECT 226.455 1678.640 226.715 1678.900 ;
      LAYER met2 ;
        RECT 206.175 1678.780 206.495 1679.235 ;
        RECT 226.425 1678.780 226.745 1678.900 ;
        RECT 206.175 1678.640 227.100 1678.780 ;
        RECT 206.175 1678.145 206.495 1678.640 ;
    END
  END mgmt_io_in_unbuf[26]
  PIN mgmt_io_in_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1683.625 206.445 1685.215 ;
      LAYER mcon ;
        RECT 206.245 1684.125 206.415 1685.215 ;
      LAYER met1 ;
        RECT 225.175 1766.915 225.315 1769.650 ;
        RECT 225.175 1766.775 225.595 1766.915 ;
        RECT 206.205 1684.065 206.465 1685.275 ;
        RECT 225.455 1684.790 225.595 1766.775 ;
        RECT 225.335 1684.470 225.595 1684.790 ;
      LAYER via ;
        RECT 206.205 1684.125 206.465 1685.215 ;
        RECT 225.335 1684.500 225.595 1684.760 ;
      LAYER met2 ;
        RECT 206.175 1684.760 206.495 1685.215 ;
        RECT 206.175 1684.620 225.975 1684.760 ;
        RECT 206.175 1684.125 206.495 1684.620 ;
        RECT 225.305 1684.500 225.625 1684.620 ;
    END
  END mgmt_io_in_unbuf[25]
  PIN mgmt_io_in_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1689.605 206.445 1691.195 ;
      LAYER mcon ;
        RECT 206.245 1690.105 206.415 1691.195 ;
      LAYER met1 ;
        RECT 224.055 1768.975 224.195 1771.650 ;
        RECT 224.055 1768.835 224.475 1768.975 ;
        RECT 206.205 1690.045 206.465 1691.255 ;
        RECT 224.335 1690.890 224.475 1768.835 ;
        RECT 224.215 1690.570 224.475 1690.890 ;
      LAYER via ;
        RECT 206.205 1690.105 206.465 1691.195 ;
        RECT 224.215 1690.600 224.475 1690.860 ;
      LAYER met2 ;
        RECT 206.175 1690.740 206.495 1691.195 ;
        RECT 224.185 1690.740 224.505 1690.860 ;
        RECT 206.175 1690.600 224.910 1690.740 ;
        RECT 206.175 1690.105 206.495 1690.600 ;
    END
  END mgmt_io_in_unbuf[24]
  PIN mgmt_io_in_unbuf[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 206.245 1695.585 206.445 1697.175 ;
      LAYER mcon ;
        RECT 206.245 1696.085 206.415 1697.175 ;
      LAYER met1 ;
        RECT 222.935 1770.850 223.075 1773.650 ;
        RECT 222.935 1770.710 223.355 1770.850 ;
        RECT 206.205 1696.025 206.465 1697.235 ;
        RECT 223.215 1696.870 223.355 1770.710 ;
        RECT 223.095 1696.550 223.355 1696.870 ;
      LAYER via ;
        RECT 206.205 1696.085 206.465 1697.175 ;
        RECT 223.095 1696.580 223.355 1696.840 ;
      LAYER met2 ;
        RECT 206.175 1696.720 206.495 1697.175 ;
        RECT 223.065 1696.720 223.385 1696.840 ;
        RECT 206.175 1696.580 223.840 1696.720 ;
        RECT 206.175 1696.085 206.495 1696.580 ;
    END
  END mgmt_io_in_unbuf[23]
  PIN mgmt_io_out_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 760.135 216.390 760.305 216.870 ;
        RECT 760.975 216.390 761.145 216.870 ;
        RECT 761.815 216.390 761.985 216.870 ;
        RECT 762.655 216.390 762.825 216.870 ;
        RECT 760.135 216.220 762.825 216.390 ;
        RECT 760.135 215.680 760.390 216.220 ;
        RECT 760.135 215.510 762.825 215.680 ;
        RECT 760.135 214.660 760.305 215.510 ;
        RECT 760.975 214.660 761.145 215.510 ;
        RECT 761.815 214.660 761.985 215.510 ;
        RECT 762.655 214.660 762.825 215.510 ;
      LAYER mcon ;
        RECT 760.220 215.510 760.390 216.360 ;
      LAYER met1 ;
        RECT 760.190 225.380 760.510 225.500 ;
        RECT 655.615 225.240 760.510 225.380 ;
        RECT 760.170 215.450 760.430 216.420 ;
      LAYER via ;
        RECT 760.220 225.240 760.480 225.500 ;
        RECT 760.170 215.510 760.430 216.360 ;
      LAYER met2 ;
        RECT 760.220 225.530 760.360 232.345 ;
        RECT 760.220 225.210 760.480 225.530 ;
        RECT 760.220 216.360 760.360 225.210 ;
        RECT 760.140 215.510 760.460 216.360 ;
    END
  END mgmt_io_out_buf[27]
  PIN mgmt_io_out_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 766.115 216.390 766.285 216.870 ;
        RECT 766.955 216.390 767.125 216.870 ;
        RECT 767.795 216.390 767.965 216.870 ;
        RECT 768.635 216.390 768.805 216.870 ;
        RECT 766.115 216.220 768.805 216.390 ;
        RECT 766.115 215.680 766.370 216.220 ;
        RECT 766.115 215.510 768.805 215.680 ;
        RECT 766.115 214.660 766.285 215.510 ;
        RECT 766.955 214.660 767.125 215.510 ;
        RECT 767.795 214.660 767.965 215.510 ;
        RECT 768.635 214.660 768.805 215.510 ;
      LAYER mcon ;
        RECT 766.200 215.510 766.370 216.360 ;
      LAYER met1 ;
        RECT 766.170 224.540 766.490 224.660 ;
        RECT 657.615 224.400 766.490 224.540 ;
        RECT 766.150 215.450 766.410 216.420 ;
      LAYER via ;
        RECT 766.200 224.400 766.460 224.660 ;
        RECT 766.150 215.510 766.410 216.360 ;
      LAYER met2 ;
        RECT 766.200 224.690 766.340 232.345 ;
        RECT 766.200 224.370 766.460 224.690 ;
        RECT 766.200 216.360 766.340 224.370 ;
        RECT 766.120 215.510 766.440 216.360 ;
    END
  END mgmt_io_out_buf[28]
  PIN mgmt_io_out_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 772.095 216.390 772.265 216.870 ;
        RECT 772.935 216.390 773.105 216.870 ;
        RECT 773.775 216.390 773.945 216.870 ;
        RECT 774.615 216.390 774.785 216.870 ;
        RECT 772.095 216.220 774.785 216.390 ;
        RECT 772.095 215.680 772.350 216.220 ;
        RECT 772.095 215.510 774.785 215.680 ;
        RECT 772.095 214.660 772.265 215.510 ;
        RECT 772.935 214.660 773.105 215.510 ;
        RECT 773.775 214.660 773.945 215.510 ;
        RECT 774.615 214.660 774.785 215.510 ;
      LAYER mcon ;
        RECT 772.180 215.510 772.350 216.360 ;
      LAYER met1 ;
        RECT 772.150 223.700 772.470 223.820 ;
        RECT 659.615 223.560 772.470 223.700 ;
        RECT 772.130 215.450 772.390 216.420 ;
      LAYER via ;
        RECT 772.180 223.560 772.440 223.820 ;
        RECT 772.130 215.510 772.390 216.360 ;
      LAYER met2 ;
        RECT 772.180 223.850 772.320 232.345 ;
        RECT 772.180 223.530 772.440 223.850 ;
        RECT 772.180 216.360 772.320 223.530 ;
        RECT 772.100 215.510 772.420 216.360 ;
    END
  END mgmt_io_out_buf[29]
  PIN mgmt_io_out_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 778.075 216.390 778.245 216.870 ;
        RECT 778.915 216.390 779.085 216.870 ;
        RECT 779.755 216.390 779.925 216.870 ;
        RECT 780.595 216.390 780.765 216.870 ;
        RECT 778.075 216.220 780.765 216.390 ;
        RECT 778.075 215.680 778.330 216.220 ;
        RECT 778.075 215.510 780.765 215.680 ;
        RECT 778.075 214.660 778.245 215.510 ;
        RECT 778.915 214.660 779.085 215.510 ;
        RECT 779.755 214.660 779.925 215.510 ;
        RECT 780.595 214.660 780.765 215.510 ;
      LAYER mcon ;
        RECT 778.160 215.510 778.330 216.360 ;
      LAYER met1 ;
        RECT 778.130 222.860 778.450 222.980 ;
        RECT 661.615 222.720 778.450 222.860 ;
        RECT 778.110 215.450 778.370 216.420 ;
      LAYER via ;
        RECT 778.160 222.720 778.420 222.980 ;
        RECT 778.110 215.510 778.370 216.360 ;
      LAYER met2 ;
        RECT 778.160 223.010 778.300 232.345 ;
        RECT 778.160 222.690 778.420 223.010 ;
        RECT 778.160 216.360 778.300 222.690 ;
        RECT 778.080 215.510 778.400 216.360 ;
    END
  END mgmt_io_out_buf[30]
  PIN mgmt_io_in_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 783.220 212.760 784.320 212.960 ;
      LAYER mcon ;
        RECT 783.230 212.790 784.320 212.960 ;
      LAYER met1 ;
        RECT 783.490 222.580 783.810 222.700 ;
        RECT 666.300 222.440 783.810 222.580 ;
        RECT 662.755 222.300 666.440 222.440 ;
        RECT 783.170 212.750 784.380 213.010 ;
      LAYER via ;
        RECT 783.520 222.440 783.780 222.700 ;
        RECT 783.230 212.750 784.320 213.010 ;
      LAYER met2 ;
        RECT 783.520 222.730 783.660 232.345 ;
        RECT 783.520 222.410 783.780 222.730 ;
        RECT 783.520 213.040 783.660 222.410 ;
        RECT 783.230 212.720 784.320 213.040 ;
    END
  END mgmt_io_in_unbuf[30]
  PIN mgmt_io_in_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 777.240 212.760 778.340 212.960 ;
      LAYER mcon ;
        RECT 777.250 212.790 778.340 212.960 ;
      LAYER met1 ;
        RECT 777.510 223.420 777.830 223.540 ;
        RECT 664.260 223.280 777.830 223.420 ;
        RECT 660.755 223.140 664.400 223.280 ;
        RECT 777.190 212.750 778.400 213.010 ;
      LAYER via ;
        RECT 777.540 223.280 777.800 223.540 ;
        RECT 777.250 212.750 778.340 213.010 ;
      LAYER met2 ;
        RECT 777.540 223.570 777.680 232.345 ;
        RECT 777.540 223.250 777.800 223.570 ;
        RECT 777.540 213.040 777.680 223.250 ;
        RECT 777.250 212.720 778.340 213.040 ;
    END
  END mgmt_io_in_unbuf[29]
  PIN mgmt_io_in_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 771.260 212.760 772.360 212.960 ;
      LAYER mcon ;
        RECT 771.270 212.790 772.360 212.960 ;
      LAYER met1 ;
        RECT 771.530 224.260 771.850 224.380 ;
        RECT 662.235 224.120 771.850 224.260 ;
        RECT 658.755 223.980 662.375 224.120 ;
        RECT 771.210 212.750 772.420 213.010 ;
      LAYER via ;
        RECT 771.560 224.120 771.820 224.380 ;
        RECT 771.270 212.750 772.360 213.010 ;
      LAYER met2 ;
        RECT 771.560 224.410 771.700 232.345 ;
        RECT 771.560 224.090 771.820 224.410 ;
        RECT 771.560 213.040 771.700 224.090 ;
        RECT 771.270 212.720 772.360 213.040 ;
    END
  END mgmt_io_in_unbuf[28]
  PIN mgmt_io_in_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 765.280 212.760 766.380 212.960 ;
      LAYER mcon ;
        RECT 765.290 212.790 766.380 212.960 ;
      LAYER met1 ;
        RECT 765.550 225.100 765.870 225.220 ;
        RECT 660.230 224.960 765.870 225.100 ;
        RECT 656.755 224.820 660.370 224.960 ;
        RECT 765.230 212.750 766.440 213.010 ;
      LAYER via ;
        RECT 765.580 224.960 765.840 225.220 ;
        RECT 765.290 212.750 766.380 213.010 ;
      LAYER met2 ;
        RECT 765.580 225.250 765.720 232.345 ;
        RECT 765.580 224.930 765.840 225.250 ;
        RECT 765.580 213.040 765.720 224.930 ;
        RECT 765.290 212.720 766.380 213.040 ;
    END
  END mgmt_io_in_unbuf[27]
  PIN mgmt_io_oeb_buf[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 784.055 216.390 784.225 216.870 ;
        RECT 784.895 216.390 785.065 216.870 ;
        RECT 785.735 216.390 785.905 216.870 ;
        RECT 786.575 216.390 786.745 216.870 ;
        RECT 784.055 216.220 786.745 216.390 ;
        RECT 784.055 215.680 784.310 216.220 ;
        RECT 784.055 215.510 786.745 215.680 ;
        RECT 784.055 214.660 784.225 215.510 ;
        RECT 784.895 214.660 785.065 215.510 ;
        RECT 785.735 214.660 785.905 215.510 ;
        RECT 786.575 214.660 786.745 215.510 ;
      LAYER mcon ;
        RECT 784.140 215.510 784.310 216.360 ;
      LAYER met1 ;
        RECT 784.110 222.020 784.430 222.140 ;
        RECT 667.215 221.880 784.430 222.020 ;
        RECT 663.755 221.740 667.355 221.880 ;
        RECT 784.090 215.450 784.350 216.420 ;
      LAYER via ;
        RECT 784.140 221.880 784.400 222.140 ;
        RECT 784.090 215.510 784.350 216.360 ;
      LAYER met2 ;
        RECT 784.140 222.170 784.280 232.345 ;
        RECT 784.140 221.850 784.400 222.170 ;
        RECT 784.140 216.360 784.280 221.850 ;
        RECT 784.060 215.510 784.380 216.360 ;
    END
  END mgmt_io_oeb_buf[0]
  PIN mgmt_io_oeb_buf[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 213.300 790.205 214.150 ;
        RECT 790.875 213.300 791.045 214.150 ;
        RECT 791.715 213.300 791.885 214.150 ;
        RECT 792.555 213.300 792.725 214.150 ;
        RECT 790.035 213.130 792.725 213.300 ;
        RECT 790.035 212.590 790.290 213.130 ;
        RECT 790.035 212.420 792.725 212.590 ;
        RECT 790.035 211.940 790.205 212.420 ;
        RECT 790.875 211.940 791.045 212.420 ;
        RECT 791.715 211.940 791.885 212.420 ;
        RECT 792.555 211.940 792.725 212.420 ;
      LAYER mcon ;
        RECT 790.120 212.450 790.290 213.300 ;
      LAYER met1 ;
        RECT 789.470 221.460 789.790 221.580 ;
        RECT 668.245 221.320 789.790 221.460 ;
        RECT 664.755 221.180 668.385 221.320 ;
        RECT 790.080 212.390 790.340 213.360 ;
      LAYER via ;
        RECT 789.500 221.320 789.760 221.580 ;
        RECT 790.080 212.450 790.340 213.300 ;
      LAYER met2 ;
        RECT 789.500 221.610 789.640 232.345 ;
        RECT 789.500 221.290 789.760 221.610 ;
        RECT 789.500 214.240 789.640 221.290 ;
        RECT 789.500 214.100 790.275 214.240 ;
        RECT 790.135 213.300 790.275 214.100 ;
        RECT 790.050 212.450 790.370 213.300 ;
    END
  END mgmt_io_oeb_buf[1]
  PIN mgmt_io_oeb_buf[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 216.390 790.205 216.870 ;
        RECT 790.875 216.390 791.045 216.870 ;
        RECT 791.715 216.390 791.885 216.870 ;
        RECT 792.555 216.390 792.725 216.870 ;
        RECT 790.035 216.220 792.725 216.390 ;
        RECT 790.035 215.680 790.290 216.220 ;
        RECT 790.035 215.510 792.725 215.680 ;
        RECT 790.035 214.660 790.205 215.510 ;
        RECT 790.875 214.660 791.045 215.510 ;
        RECT 791.715 214.660 791.885 215.510 ;
        RECT 792.555 214.660 792.725 215.510 ;
      LAYER mcon ;
        RECT 790.120 215.510 790.290 216.360 ;
      LAYER met1 ;
        RECT 790.090 220.900 790.410 221.020 ;
        RECT 669.190 220.760 790.410 220.900 ;
        RECT 665.755 220.620 669.330 220.760 ;
        RECT 790.070 215.450 790.330 216.420 ;
      LAYER via ;
        RECT 790.120 220.760 790.380 221.020 ;
        RECT 790.070 215.510 790.330 216.360 ;
      LAYER met2 ;
        RECT 790.120 221.050 790.260 232.345 ;
        RECT 790.120 220.730 790.380 221.050 ;
        RECT 790.120 216.360 790.260 220.730 ;
        RECT 790.040 215.510 790.360 216.360 ;
    END
  END mgmt_io_oeb_buf[2]
  PIN mgmt_io_oeb_unbuf[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2270.340 215.850 2271.930 216.050 ;
      LAYER mcon ;
        RECT 2270.840 215.850 2271.930 216.020 ;
      LAYER met1 ;
        RECT 2271.305 221.040 2416.200 221.180 ;
        RECT 2271.305 220.920 2271.625 221.040 ;
        RECT 2270.780 215.810 2271.990 216.070 ;
        RECT 2416.060 211.780 2416.200 221.040 ;
        RECT 3377.640 212.245 3377.780 1161.450 ;
        RECT 2537.220 212.105 3377.780 212.245 ;
        RECT 2537.220 211.780 2537.360 212.105 ;
        RECT 2416.060 211.640 2537.360 211.780 ;
      LAYER via ;
        RECT 2271.335 220.920 2271.595 221.180 ;
        RECT 2270.840 215.810 2271.930 216.070 ;
      LAYER met2 ;
        RECT 2271.335 221.210 2271.475 232.485 ;
        RECT 2271.335 220.890 2271.595 221.210 ;
        RECT 2271.335 216.100 2271.475 220.890 ;
        RECT 2270.840 215.780 2271.930 216.100 ;
    END
  END mgmt_io_oeb_unbuf[2]
  PIN mgmt_io_oeb_unbuf[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2270.340 212.760 2271.440 212.960 ;
      LAYER mcon ;
        RECT 2270.340 212.790 2271.430 212.960 ;
      LAYER met1 ;
        RECT 2270.335 221.600 2417.040 221.740 ;
        RECT 2270.335 221.480 2270.655 221.600 ;
        RECT 2270.280 212.750 2271.490 213.010 ;
        RECT 2416.900 212.060 2417.040 221.600 ;
        RECT 3376.800 212.740 3376.940 1160.450 ;
        RECT 2536.380 212.600 3376.940 212.740 ;
        RECT 2536.380 212.060 2536.520 212.600 ;
        RECT 2416.900 211.920 2536.520 212.060 ;
      LAYER via ;
        RECT 2270.365 221.480 2270.625 221.740 ;
        RECT 2270.340 212.750 2271.430 213.010 ;
      LAYER met2 ;
        RECT 2270.365 221.770 2270.505 232.485 ;
        RECT 2270.365 221.450 2270.625 221.770 ;
        RECT 2270.365 214.170 2270.505 221.450 ;
        RECT 2270.365 214.030 2271.140 214.170 ;
        RECT 2271.000 213.040 2271.140 214.030 ;
        RECT 2270.340 212.720 2271.430 213.040 ;
    END
  END mgmt_io_oeb_unbuf[1]
  PIN mgmt_io_oeb_unbuf[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2264.360 215.850 2265.950 216.050 ;
      LAYER mcon ;
        RECT 2264.860 215.850 2265.950 216.020 ;
      LAYER met1 ;
        RECT 2265.205 222.160 2417.880 222.300 ;
        RECT 2265.205 222.040 2265.525 222.160 ;
        RECT 2264.800 215.810 2266.010 216.070 ;
        RECT 2417.740 212.340 2417.880 222.160 ;
        RECT 3375.960 213.300 3376.100 1159.440 ;
        RECT 2535.540 213.160 3376.100 213.300 ;
        RECT 2535.540 212.340 2535.680 213.160 ;
        RECT 2417.740 212.200 2535.680 212.340 ;
      LAYER via ;
        RECT 2265.235 222.040 2265.495 222.300 ;
        RECT 2264.860 215.810 2265.950 216.070 ;
      LAYER met2 ;
        RECT 2265.355 222.330 2265.495 232.485 ;
        RECT 2265.235 222.010 2265.495 222.330 ;
        RECT 2265.355 216.100 2265.495 222.010 ;
        RECT 2264.860 215.780 2265.950 216.100 ;
    END
  END mgmt_io_oeb_unbuf[0]
  PIN mgmt_io_in_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2261.935 213.300 2262.105 214.150 ;
        RECT 2262.775 213.300 2262.945 214.150 ;
        RECT 2263.615 213.300 2263.785 214.150 ;
        RECT 2264.455 213.300 2264.625 214.150 ;
        RECT 2261.935 213.130 2264.625 213.300 ;
        RECT 2264.370 212.590 2264.625 213.130 ;
        RECT 2261.935 212.420 2264.625 212.590 ;
        RECT 2261.935 211.940 2262.105 212.420 ;
        RECT 2262.775 211.940 2262.945 212.420 ;
        RECT 2263.615 211.940 2263.785 212.420 ;
        RECT 2264.455 211.940 2264.625 212.420 ;
      LAYER mcon ;
        RECT 2264.370 212.450 2264.540 213.300 ;
      LAYER met1 ;
        RECT 3375.400 1154.570 3375.540 1158.450 ;
        RECT 3375.120 1154.430 3375.540 1154.570 ;
        RECT 2264.355 222.720 2418.720 222.860 ;
        RECT 2264.355 222.600 2264.675 222.720 ;
        RECT 2264.320 212.390 2264.580 213.360 ;
        RECT 2418.580 212.620 2418.720 222.720 ;
        RECT 3375.120 213.860 3375.260 1154.430 ;
        RECT 2534.700 213.720 3375.260 213.860 ;
        RECT 2534.700 212.620 2534.840 213.720 ;
        RECT 2418.580 212.480 2534.840 212.620 ;
      LAYER via ;
        RECT 2264.385 222.600 2264.645 222.860 ;
        RECT 2264.320 212.450 2264.580 213.300 ;
      LAYER met2 ;
        RECT 2264.385 222.890 2264.525 232.485 ;
        RECT 2264.385 222.570 2264.645 222.890 ;
        RECT 2264.385 213.300 2264.525 222.570 ;
        RECT 2264.290 212.450 2264.610 213.300 ;
    END
  END mgmt_io_in_buf[30]
  PIN mgmt_io_in_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2255.955 213.300 2256.125 214.150 ;
        RECT 2256.795 213.300 2256.965 214.150 ;
        RECT 2257.635 213.300 2257.805 214.150 ;
        RECT 2258.475 213.300 2258.645 214.150 ;
        RECT 2255.955 213.130 2258.645 213.300 ;
        RECT 2258.390 212.590 2258.645 213.130 ;
        RECT 2255.955 212.420 2258.645 212.590 ;
        RECT 2255.955 211.940 2256.125 212.420 ;
        RECT 2256.795 211.940 2256.965 212.420 ;
        RECT 2257.635 211.940 2257.805 212.420 ;
        RECT 2258.475 211.940 2258.645 212.420 ;
      LAYER mcon ;
        RECT 2258.390 212.450 2258.560 213.300 ;
      LAYER met1 ;
        RECT 3374.280 1152.510 3374.420 1156.450 ;
        RECT 3374.000 1152.370 3374.420 1152.510 ;
        RECT 2258.375 223.560 2419.840 223.700 ;
        RECT 2258.375 223.440 2258.695 223.560 ;
        RECT 2258.340 212.390 2258.600 213.360 ;
        RECT 2419.695 213.180 2419.835 223.560 ;
        RECT 3374.000 214.700 3374.140 1152.370 ;
        RECT 2533.580 214.560 3374.140 214.700 ;
        RECT 2533.580 213.180 2533.720 214.560 ;
        RECT 2419.695 213.040 2533.720 213.180 ;
      LAYER via ;
        RECT 2258.405 223.440 2258.665 223.700 ;
        RECT 2258.340 212.450 2258.600 213.300 ;
      LAYER met2 ;
        RECT 2258.405 223.730 2258.545 232.485 ;
        RECT 2258.405 223.410 2258.665 223.730 ;
        RECT 2258.405 213.300 2258.545 223.410 ;
        RECT 2258.310 212.450 2258.630 213.300 ;
    END
  END mgmt_io_in_buf[29]
  PIN mgmt_io_in_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2249.975 213.300 2250.145 214.150 ;
        RECT 2250.815 213.300 2250.985 214.150 ;
        RECT 2251.655 213.300 2251.825 214.150 ;
        RECT 2252.495 213.300 2252.665 214.150 ;
        RECT 2249.975 213.130 2252.665 213.300 ;
        RECT 2252.410 212.590 2252.665 213.130 ;
        RECT 2249.975 212.420 2252.665 212.590 ;
        RECT 2249.975 211.940 2250.145 212.420 ;
        RECT 2250.815 211.940 2250.985 212.420 ;
        RECT 2251.655 211.940 2251.825 212.420 ;
        RECT 2252.495 211.940 2252.665 212.420 ;
      LAYER mcon ;
        RECT 2252.410 212.450 2252.580 213.300 ;
      LAYER met1 ;
        RECT 3373.160 1150.590 3373.300 1154.440 ;
        RECT 3372.880 1150.450 3373.300 1150.590 ;
        RECT 2252.395 224.400 2420.960 224.540 ;
        RECT 2252.395 224.280 2252.715 224.400 ;
        RECT 2420.820 213.740 2420.960 224.400 ;
        RECT 3372.880 215.540 3373.020 1150.450 ;
        RECT 2532.460 215.400 3373.020 215.540 ;
        RECT 2532.460 213.740 2532.600 215.400 ;
        RECT 2420.820 213.600 2532.600 213.740 ;
        RECT 2252.360 212.390 2252.620 213.360 ;
      LAYER via ;
        RECT 2252.425 224.280 2252.685 224.540 ;
        RECT 2252.360 212.450 2252.620 213.300 ;
      LAYER met2 ;
        RECT 2252.425 224.570 2252.565 232.485 ;
        RECT 2252.425 224.250 2252.685 224.570 ;
        RECT 2252.425 213.300 2252.565 224.250 ;
        RECT 2252.330 212.450 2252.650 213.300 ;
    END
  END mgmt_io_in_buf[28]
  PIN mgmt_io_in_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2243.995 213.300 2244.165 214.150 ;
        RECT 2244.835 213.300 2245.005 214.150 ;
        RECT 2245.675 213.300 2245.845 214.150 ;
        RECT 2246.515 213.300 2246.685 214.150 ;
        RECT 2243.995 213.130 2246.685 213.300 ;
        RECT 2246.430 212.590 2246.685 213.130 ;
        RECT 2243.995 212.420 2246.685 212.590 ;
        RECT 2243.995 211.940 2244.165 212.420 ;
        RECT 2244.835 211.940 2245.005 212.420 ;
        RECT 2245.675 211.940 2245.845 212.420 ;
        RECT 2246.515 211.940 2246.685 212.420 ;
      LAYER mcon ;
        RECT 2246.430 212.450 2246.600 213.300 ;
      LAYER met1 ;
        RECT 3372.040 1148.550 3372.180 1152.440 ;
        RECT 3371.760 1148.410 3372.180 1148.550 ;
        RECT 2246.415 225.240 2422.080 225.380 ;
        RECT 2246.415 225.120 2246.735 225.240 ;
        RECT 2421.940 214.300 2422.080 225.240 ;
        RECT 3371.760 216.380 3371.900 1148.410 ;
        RECT 2531.340 216.240 3371.900 216.380 ;
        RECT 2531.340 214.300 2531.480 216.240 ;
        RECT 2421.940 214.160 2531.480 214.300 ;
        RECT 2246.380 212.390 2246.640 213.360 ;
      LAYER via ;
        RECT 2246.445 225.120 2246.705 225.380 ;
        RECT 2246.380 212.450 2246.640 213.300 ;
      LAYER met2 ;
        RECT 2246.445 225.410 2246.585 232.485 ;
        RECT 2246.445 225.090 2246.705 225.410 ;
        RECT 2246.445 213.300 2246.585 225.090 ;
        RECT 2246.350 212.450 2246.670 213.300 ;
    END
  END mgmt_io_in_buf[27]
  PIN mgmt_io_out_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2240.440 215.850 2242.030 216.050 ;
      LAYER mcon ;
        RECT 2240.940 215.850 2242.030 216.020 ;
      LAYER met1 ;
        RECT 2241.405 225.520 2422.360 225.660 ;
        RECT 2241.405 225.400 2241.725 225.520 ;
        RECT 2240.880 215.810 2242.090 216.070 ;
        RECT 2422.220 214.580 2422.360 225.520 ;
        RECT 3371.480 216.660 3371.620 1151.440 ;
        RECT 2531.060 216.520 3371.620 216.660 ;
        RECT 2531.060 214.580 2531.200 216.520 ;
        RECT 2422.220 214.440 2531.200 214.580 ;
      LAYER via ;
        RECT 2241.435 225.400 2241.695 225.660 ;
        RECT 2240.940 215.810 2242.030 216.070 ;
      LAYER met2 ;
        RECT 2241.435 225.690 2241.575 232.485 ;
        RECT 2241.435 225.370 2241.695 225.690 ;
        RECT 2241.435 216.100 2241.575 225.370 ;
        RECT 2240.940 215.780 2242.030 216.100 ;
    END
  END mgmt_io_out_unbuf[27]
  PIN mgmt_io_out_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2246.420 215.850 2248.010 216.050 ;
      LAYER mcon ;
        RECT 2246.920 215.850 2248.010 216.020 ;
      LAYER met1 ;
        RECT 2247.385 224.680 2421.240 224.820 ;
        RECT 2247.385 224.560 2247.705 224.680 ;
        RECT 2246.860 215.810 2248.070 216.070 ;
        RECT 2421.100 214.020 2421.240 224.680 ;
        RECT 3372.600 215.820 3372.740 1153.450 ;
        RECT 2532.180 215.680 3372.740 215.820 ;
        RECT 2532.180 214.020 2532.320 215.680 ;
        RECT 2421.100 213.880 2532.320 214.020 ;
      LAYER via ;
        RECT 2247.415 224.560 2247.675 224.820 ;
        RECT 2246.920 215.810 2248.010 216.070 ;
      LAYER met2 ;
        RECT 2247.415 224.850 2247.555 232.485 ;
        RECT 2247.415 224.530 2247.675 224.850 ;
        RECT 2247.415 216.100 2247.555 224.530 ;
        RECT 2246.920 215.780 2248.010 216.100 ;
    END
  END mgmt_io_out_unbuf[28]
  PIN mgmt_io_out_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2252.400 215.850 2253.990 216.050 ;
      LAYER mcon ;
        RECT 2252.900 215.850 2253.990 216.020 ;
      LAYER met1 ;
        RECT 2253.245 223.840 2420.120 223.980 ;
        RECT 2253.245 223.720 2253.565 223.840 ;
        RECT 2252.840 215.810 2254.050 216.070 ;
        RECT 2419.980 213.460 2420.120 223.840 ;
        RECT 3373.720 214.980 3373.860 1155.440 ;
        RECT 2533.300 214.840 3373.860 214.980 ;
        RECT 2533.300 213.460 2533.440 214.840 ;
        RECT 2419.980 213.320 2533.440 213.460 ;
      LAYER via ;
        RECT 2253.275 223.720 2253.535 223.980 ;
        RECT 2252.900 215.810 2253.990 216.070 ;
      LAYER met2 ;
        RECT 2253.395 224.010 2253.535 232.485 ;
        RECT 2253.275 223.690 2253.535 224.010 ;
        RECT 2253.395 216.100 2253.535 223.690 ;
        RECT 2252.900 215.780 2253.990 216.100 ;
    END
  END mgmt_io_out_unbuf[29]
  PIN mgmt_io_out_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2258.380 215.850 2259.970 216.050 ;
      LAYER mcon ;
        RECT 2258.880 215.850 2259.970 216.020 ;
      LAYER met1 ;
        RECT 2259.345 223.000 2419.000 223.140 ;
        RECT 2259.345 222.880 2259.665 223.000 ;
        RECT 2258.820 215.810 2260.030 216.070 ;
        RECT 2418.860 212.900 2419.000 223.000 ;
        RECT 3374.840 214.140 3374.980 1157.450 ;
        RECT 2534.420 214.000 3374.980 214.140 ;
        RECT 2534.420 212.900 2534.560 214.000 ;
        RECT 2418.860 212.760 2534.560 212.900 ;
      LAYER via ;
        RECT 2259.375 222.880 2259.635 223.140 ;
        RECT 2258.880 215.810 2259.970 216.070 ;
      LAYER met2 ;
        RECT 2259.375 223.170 2259.515 232.485 ;
        RECT 2259.375 222.850 2259.635 223.170 ;
        RECT 2259.375 216.100 2259.515 222.850 ;
        RECT 2258.880 215.780 2259.970 216.100 ;
    END
  END mgmt_io_out_unbuf[30]
  PIN mgmt_io_out_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2150.740 215.850 2152.330 216.050 ;
      LAYER mcon ;
        RECT 2151.240 215.850 2152.330 216.020 ;
      LAYER met1 ;
        RECT 2151.705 238.120 2439.160 238.260 ;
        RECT 2151.705 238.000 2152.025 238.120 ;
        RECT 2439.020 222.980 2439.160 238.120 ;
        RECT 3354.680 229.260 3354.820 1121.750 ;
        RECT 2514.260 229.120 3354.820 229.260 ;
        RECT 2514.260 222.980 2514.400 229.120 ;
        RECT 2439.020 222.840 2514.400 222.980 ;
        RECT 2151.180 215.810 2152.390 216.070 ;
      LAYER via ;
        RECT 2151.735 238.000 2151.995 238.260 ;
        RECT 2151.240 215.810 2152.330 216.070 ;
      LAYER met2 ;
        RECT 2151.735 238.290 2151.875 238.365 ;
        RECT 2151.735 237.970 2151.995 238.290 ;
        RECT 2151.735 216.100 2151.875 237.970 ;
        RECT 2151.240 215.780 2152.330 216.100 ;
    END
  END mgmt_io_out_unbuf[26]
  PIN mgmt_io_out_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2156.720 215.850 2158.310 216.050 ;
      LAYER mcon ;
        RECT 2157.220 215.850 2158.310 216.020 ;
      LAYER met1 ;
        RECT 2157.685 237.280 2438.040 237.420 ;
        RECT 2157.685 237.160 2158.005 237.280 ;
        RECT 2437.900 222.420 2438.040 237.280 ;
        RECT 3355.800 228.420 3355.940 1123.700 ;
        RECT 2515.380 228.280 3355.940 228.420 ;
        RECT 2515.380 222.420 2515.520 228.280 ;
        RECT 2437.900 222.280 2515.520 222.420 ;
        RECT 2157.160 215.810 2158.370 216.070 ;
      LAYER via ;
        RECT 2157.715 237.160 2157.975 237.420 ;
        RECT 2157.220 215.810 2158.310 216.070 ;
      LAYER met2 ;
        RECT 2157.715 237.450 2157.855 237.575 ;
        RECT 2157.715 237.130 2157.975 237.450 ;
        RECT 2157.715 216.100 2157.855 237.130 ;
        RECT 2157.220 215.780 2158.310 216.100 ;
    END
  END mgmt_io_out_unbuf[25]
  PIN mgmt_io_out_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2162.700 215.850 2164.290 216.050 ;
      LAYER mcon ;
        RECT 2163.200 215.850 2164.290 216.020 ;
      LAYER met1 ;
        RECT 2163.665 236.440 2436.920 236.580 ;
        RECT 2163.665 236.320 2163.985 236.440 ;
        RECT 2436.780 221.860 2436.920 236.440 ;
        RECT 3356.920 227.580 3357.060 1125.690 ;
        RECT 2516.500 227.440 3357.060 227.580 ;
        RECT 2516.500 221.860 2516.640 227.440 ;
        RECT 2436.780 221.720 2516.640 221.860 ;
        RECT 2163.140 215.810 2164.350 216.070 ;
      LAYER via ;
        RECT 2163.695 236.320 2163.955 236.580 ;
        RECT 2163.200 215.810 2164.290 216.070 ;
      LAYER met2 ;
        RECT 2163.695 236.610 2163.835 236.720 ;
        RECT 2163.695 236.290 2163.955 236.610 ;
        RECT 2163.695 216.100 2163.835 236.290 ;
        RECT 2163.200 215.780 2164.290 216.100 ;
    END
  END mgmt_io_out_unbuf[24]
  PIN mgmt_io_out_unbuf[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2168.680 215.850 2170.270 216.050 ;
      LAYER mcon ;
        RECT 2169.180 215.850 2170.270 216.020 ;
      LAYER met1 ;
        RECT 2169.645 235.600 2435.800 235.740 ;
        RECT 2169.645 235.480 2169.965 235.600 ;
        RECT 2435.660 221.300 2435.800 235.600 ;
        RECT 3358.040 226.740 3358.180 1127.710 ;
        RECT 2517.620 226.600 3358.180 226.740 ;
        RECT 2517.620 221.300 2517.760 226.600 ;
        RECT 2435.660 221.160 2517.760 221.300 ;
        RECT 2169.120 215.810 2170.330 216.070 ;
      LAYER via ;
        RECT 2169.675 235.480 2169.935 235.740 ;
        RECT 2169.180 215.810 2170.270 216.070 ;
      LAYER met2 ;
        RECT 2169.675 235.770 2169.815 235.930 ;
        RECT 2169.675 235.450 2169.935 235.770 ;
        RECT 2169.675 216.100 2169.815 235.450 ;
        RECT 2169.180 215.780 2170.270 216.100 ;
    END
  END mgmt_io_out_unbuf[23]
  PIN mgmt_io_out_unbuf[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2174.660 215.850 2176.250 216.050 ;
      LAYER mcon ;
        RECT 2175.160 215.850 2176.250 216.020 ;
      LAYER met1 ;
        RECT 2175.625 234.760 2434.680 234.900 ;
        RECT 2175.625 234.640 2175.945 234.760 ;
        RECT 2434.540 220.740 2434.680 234.760 ;
        RECT 3359.160 225.900 3359.300 1129.680 ;
        RECT 2518.740 225.760 3359.300 225.900 ;
        RECT 2518.740 220.740 2518.880 225.760 ;
        RECT 2434.540 220.600 2518.880 220.740 ;
        RECT 2175.100 215.810 2176.310 216.070 ;
      LAYER via ;
        RECT 2175.655 234.640 2175.915 234.900 ;
        RECT 2175.160 215.810 2176.250 216.070 ;
      LAYER met2 ;
        RECT 2175.655 234.930 2175.795 235.010 ;
        RECT 2175.655 234.610 2175.915 234.930 ;
        RECT 2175.655 216.100 2175.795 234.610 ;
        RECT 2175.160 215.780 2176.250 216.100 ;
    END
  END mgmt_io_out_unbuf[22]
  PIN mgmt_io_out_unbuf[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2180.640 215.850 2182.230 216.050 ;
      LAYER mcon ;
        RECT 2181.140 215.850 2182.230 216.020 ;
      LAYER met1 ;
        RECT 2181.485 233.920 2433.560 234.060 ;
        RECT 2181.485 233.800 2181.805 233.920 ;
        RECT 2433.420 220.180 2433.560 233.920 ;
        RECT 3360.280 225.060 3360.420 1131.700 ;
        RECT 2519.860 224.920 3360.420 225.060 ;
        RECT 2519.860 220.180 2520.000 224.920 ;
        RECT 2433.420 220.040 2520.000 220.180 ;
        RECT 2181.080 215.810 2182.290 216.070 ;
      LAYER via ;
        RECT 2181.515 233.800 2181.775 234.060 ;
        RECT 2181.140 215.810 2182.230 216.070 ;
      LAYER met2 ;
        RECT 2181.635 234.090 2181.775 234.200 ;
        RECT 2181.515 233.770 2181.775 234.090 ;
        RECT 2181.635 216.100 2181.775 233.770 ;
        RECT 2181.140 215.780 2182.230 216.100 ;
    END
  END mgmt_io_out_unbuf[21]
  PIN mgmt_io_out_unbuf[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2186.620 215.850 2188.210 216.050 ;
      LAYER mcon ;
        RECT 2187.120 215.850 2188.210 216.020 ;
      LAYER met1 ;
        RECT 2187.585 233.080 2432.440 233.220 ;
        RECT 2187.585 232.960 2187.905 233.080 ;
        RECT 2432.300 219.620 2432.440 233.080 ;
        RECT 3361.400 224.220 3361.540 1133.690 ;
        RECT 2520.980 224.080 3361.540 224.220 ;
        RECT 2520.980 219.620 2521.120 224.080 ;
        RECT 2432.300 219.480 2521.120 219.620 ;
        RECT 2187.060 215.810 2188.270 216.070 ;
      LAYER via ;
        RECT 2187.615 232.960 2187.875 233.220 ;
        RECT 2187.120 215.810 2188.210 216.070 ;
      LAYER met2 ;
        RECT 2187.615 233.250 2187.755 233.365 ;
        RECT 2187.615 232.930 2187.875 233.250 ;
        RECT 2187.615 216.100 2187.755 232.930 ;
        RECT 2187.120 215.780 2188.210 216.100 ;
    END
  END mgmt_io_out_unbuf[20]
  PIN mgmt_io_out_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2192.600 215.850 2194.190 216.050 ;
      LAYER mcon ;
        RECT 2193.100 215.850 2194.190 216.020 ;
      LAYER met1 ;
        RECT 2193.445 232.240 2431.320 232.380 ;
        RECT 2193.445 232.120 2193.765 232.240 ;
        RECT 2431.180 219.060 2431.320 232.240 ;
        RECT 3362.520 223.380 3362.660 1135.690 ;
        RECT 2522.100 223.240 3362.660 223.380 ;
        RECT 2522.100 219.060 2522.240 223.240 ;
        RECT 2431.180 218.920 2522.240 219.060 ;
        RECT 2193.040 215.810 2194.250 216.070 ;
      LAYER via ;
        RECT 2193.475 232.120 2193.735 232.380 ;
        RECT 2193.100 215.810 2194.190 216.070 ;
      LAYER met2 ;
        RECT 2193.595 232.410 2193.735 232.485 ;
        RECT 2193.475 232.090 2193.735 232.410 ;
        RECT 2193.595 216.100 2193.735 232.090 ;
        RECT 2193.100 215.780 2194.190 216.100 ;
    END
  END mgmt_io_out_unbuf[19]
  PIN mgmt_io_out_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2198.580 215.850 2200.170 216.050 ;
      LAYER mcon ;
        RECT 2199.080 215.850 2200.170 216.020 ;
      LAYER met1 ;
        RECT 2199.545 231.400 2430.200 231.540 ;
        RECT 2199.545 231.280 2199.865 231.400 ;
        RECT 2430.060 218.500 2430.200 231.400 ;
        RECT 3363.640 222.540 3363.780 1137.690 ;
        RECT 2523.220 222.400 3363.780 222.540 ;
        RECT 2523.220 218.500 2523.360 222.400 ;
        RECT 2430.060 218.360 2523.360 218.500 ;
        RECT 2199.020 215.810 2200.230 216.070 ;
      LAYER via ;
        RECT 2199.575 231.280 2199.835 231.540 ;
        RECT 2199.080 215.810 2200.170 216.070 ;
      LAYER met2 ;
        RECT 2199.575 231.570 2199.715 232.485 ;
        RECT 2199.575 231.250 2199.835 231.570 ;
        RECT 2199.575 216.100 2199.715 231.250 ;
        RECT 2199.080 215.780 2200.170 216.100 ;
    END
  END mgmt_io_out_unbuf[18]
  PIN mgmt_io_out_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2204.560 215.850 2206.150 216.050 ;
      LAYER mcon ;
        RECT 2205.060 215.850 2206.150 216.020 ;
      LAYER met1 ;
        RECT 2205.525 230.560 2429.080 230.700 ;
        RECT 2205.525 230.440 2205.845 230.560 ;
        RECT 2428.940 217.940 2429.080 230.560 ;
        RECT 3364.760 221.700 3364.900 1139.690 ;
        RECT 2524.340 221.560 3364.900 221.700 ;
        RECT 2524.340 217.940 2524.480 221.560 ;
        RECT 2428.940 217.800 2524.480 217.940 ;
        RECT 2205.000 215.810 2206.210 216.070 ;
      LAYER via ;
        RECT 2205.555 230.440 2205.815 230.700 ;
        RECT 2205.060 215.810 2206.150 216.070 ;
      LAYER met2 ;
        RECT 2205.555 230.730 2205.695 232.485 ;
        RECT 2205.555 230.410 2205.815 230.730 ;
        RECT 2205.555 216.100 2205.695 230.410 ;
        RECT 2205.060 215.780 2206.150 216.100 ;
    END
  END mgmt_io_out_unbuf[17]
  PIN mgmt_io_out_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2210.540 215.850 2212.130 216.050 ;
      LAYER mcon ;
        RECT 2211.040 215.850 2212.130 216.020 ;
      LAYER met1 ;
        RECT 2211.505 229.720 2427.960 229.860 ;
        RECT 2211.505 229.600 2211.825 229.720 ;
        RECT 2427.820 217.380 2427.960 229.720 ;
        RECT 3365.880 220.860 3366.020 1141.690 ;
        RECT 2525.460 220.720 3366.020 220.860 ;
        RECT 2525.460 217.380 2525.600 220.720 ;
        RECT 2427.820 217.240 2525.600 217.380 ;
        RECT 2210.980 215.810 2212.190 216.070 ;
      LAYER via ;
        RECT 2211.535 229.600 2211.795 229.860 ;
        RECT 2211.040 215.810 2212.130 216.070 ;
      LAYER met2 ;
        RECT 2211.535 229.890 2211.675 232.485 ;
        RECT 2211.535 229.570 2211.795 229.890 ;
        RECT 2211.535 216.100 2211.675 229.570 ;
        RECT 2211.040 215.780 2212.130 216.100 ;
    END
  END mgmt_io_out_unbuf[16]
  PIN mgmt_io_out_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2216.520 215.850 2218.110 216.050 ;
      LAYER mcon ;
        RECT 2217.020 215.850 2218.110 216.020 ;
      LAYER met1 ;
        RECT 2217.485 228.880 2426.840 229.020 ;
        RECT 2217.485 228.760 2217.805 228.880 ;
        RECT 2426.700 216.820 2426.840 228.880 ;
        RECT 3367.000 220.020 3367.140 1143.680 ;
        RECT 2526.580 219.880 3367.140 220.020 ;
        RECT 2526.580 216.820 2526.720 219.880 ;
        RECT 2426.700 216.680 2526.720 216.820 ;
        RECT 2216.960 215.810 2218.170 216.070 ;
      LAYER via ;
        RECT 2217.515 228.760 2217.775 229.020 ;
        RECT 2217.020 215.810 2218.110 216.070 ;
      LAYER met2 ;
        RECT 2217.515 229.050 2217.655 232.485 ;
        RECT 2217.515 228.730 2217.775 229.050 ;
        RECT 2217.515 216.100 2217.655 228.730 ;
        RECT 2217.020 215.780 2218.110 216.100 ;
    END
  END mgmt_io_out_unbuf[15]
  PIN mgmt_io_out_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2222.500 215.850 2224.090 216.050 ;
      LAYER mcon ;
        RECT 2223.000 215.850 2224.090 216.020 ;
      LAYER met1 ;
        RECT 2223.465 228.040 2425.720 228.180 ;
        RECT 2223.465 227.920 2223.785 228.040 ;
        RECT 2425.580 216.260 2425.720 228.040 ;
        RECT 3368.120 219.180 3368.260 1145.690 ;
        RECT 2527.700 219.040 3368.260 219.180 ;
        RECT 2527.700 216.260 2527.840 219.040 ;
        RECT 2425.580 216.120 2527.840 216.260 ;
        RECT 2222.940 215.810 2224.150 216.070 ;
      LAYER via ;
        RECT 2223.495 227.920 2223.755 228.180 ;
        RECT 2223.000 215.810 2224.090 216.070 ;
      LAYER met2 ;
        RECT 2223.495 228.210 2223.635 232.485 ;
        RECT 2223.495 227.890 2223.755 228.210 ;
        RECT 2223.495 216.100 2223.635 227.890 ;
        RECT 2223.000 215.780 2224.090 216.100 ;
    END
  END mgmt_io_out_unbuf[14]
  PIN mgmt_io_out_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2228.480 215.850 2230.070 216.050 ;
      LAYER mcon ;
        RECT 2228.980 215.850 2230.070 216.020 ;
      LAYER met1 ;
        RECT 2229.445 227.200 2424.600 227.340 ;
        RECT 2229.445 227.080 2229.765 227.200 ;
        RECT 2228.920 215.810 2230.130 216.070 ;
        RECT 2424.460 215.700 2424.600 227.200 ;
        RECT 3369.240 218.340 3369.380 1147.670 ;
        RECT 2528.820 218.200 3369.380 218.340 ;
        RECT 2528.820 215.700 2528.960 218.200 ;
        RECT 2424.460 215.560 2528.960 215.700 ;
      LAYER via ;
        RECT 2229.475 227.080 2229.735 227.340 ;
        RECT 2228.980 215.810 2230.070 216.070 ;
      LAYER met2 ;
        RECT 2229.475 227.370 2229.615 232.485 ;
        RECT 2229.475 227.050 2229.735 227.370 ;
        RECT 2229.475 216.100 2229.615 227.050 ;
        RECT 2228.980 215.780 2230.070 216.100 ;
    END
  END mgmt_io_out_unbuf[13]
  PIN mgmt_io_out_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2234.460 215.850 2236.050 216.050 ;
      LAYER mcon ;
        RECT 2234.960 215.850 2236.050 216.020 ;
      LAYER met1 ;
        RECT 2235.425 226.360 2423.480 226.500 ;
        RECT 2235.425 226.240 2235.745 226.360 ;
        RECT 2234.900 215.810 2236.110 216.070 ;
        RECT 2423.340 215.140 2423.480 226.360 ;
        RECT 3370.360 217.500 3370.500 1149.680 ;
        RECT 2529.940 217.360 3370.500 217.500 ;
        RECT 2529.940 215.140 2530.080 217.360 ;
        RECT 2423.340 215.000 2530.080 215.140 ;
      LAYER via ;
        RECT 2235.455 226.240 2235.715 226.500 ;
        RECT 2234.960 215.810 2236.050 216.070 ;
      LAYER met2 ;
        RECT 2235.455 226.530 2235.595 232.485 ;
        RECT 2235.455 226.210 2235.715 226.530 ;
        RECT 2235.455 216.100 2235.595 226.210 ;
        RECT 2234.960 215.780 2236.050 216.100 ;
    END
  END mgmt_io_out_unbuf[12]
  PIN mgmt_io_in_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2238.015 213.300 2238.185 214.150 ;
        RECT 2238.855 213.300 2239.025 214.150 ;
        RECT 2239.695 213.300 2239.865 214.150 ;
        RECT 2240.535 213.300 2240.705 214.150 ;
        RECT 2238.015 213.130 2240.705 213.300 ;
        RECT 2240.450 212.590 2240.705 213.130 ;
        RECT 2238.015 212.420 2240.705 212.590 ;
        RECT 2238.015 211.940 2238.185 212.420 ;
        RECT 2238.855 211.940 2239.025 212.420 ;
        RECT 2239.695 211.940 2239.865 212.420 ;
        RECT 2240.535 211.940 2240.705 212.420 ;
      LAYER mcon ;
        RECT 2240.450 212.450 2240.620 213.300 ;
      LAYER met1 ;
        RECT 3370.920 1146.470 3371.060 1150.680 ;
        RECT 3370.640 1146.330 3371.060 1146.470 ;
        RECT 2240.435 226.080 2423.200 226.220 ;
        RECT 2240.435 225.960 2240.755 226.080 ;
        RECT 2423.060 214.860 2423.200 226.080 ;
        RECT 3370.640 217.220 3370.780 1146.330 ;
        RECT 2530.220 217.080 3370.780 217.220 ;
        RECT 2530.220 214.860 2530.360 217.080 ;
        RECT 2423.060 214.720 2530.360 214.860 ;
        RECT 2240.400 212.390 2240.660 213.360 ;
      LAYER via ;
        RECT 2240.465 225.960 2240.725 226.220 ;
        RECT 2240.400 212.450 2240.660 213.300 ;
      LAYER met2 ;
        RECT 2240.465 226.250 2240.605 232.485 ;
        RECT 2240.465 225.930 2240.725 226.250 ;
        RECT 2240.465 213.300 2240.605 225.930 ;
        RECT 2240.370 212.450 2240.690 213.300 ;
    END
  END mgmt_io_in_buf[12]
  PIN mgmt_io_in_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2232.035 213.300 2232.205 214.150 ;
        RECT 2232.875 213.300 2233.045 214.150 ;
        RECT 2233.715 213.300 2233.885 214.150 ;
        RECT 2234.555 213.300 2234.725 214.150 ;
        RECT 2232.035 213.130 2234.725 213.300 ;
        RECT 2234.470 212.590 2234.725 213.130 ;
        RECT 2232.035 212.420 2234.725 212.590 ;
        RECT 2232.035 211.940 2232.205 212.420 ;
        RECT 2232.875 211.940 2233.045 212.420 ;
        RECT 2233.715 211.940 2233.885 212.420 ;
        RECT 2234.555 211.940 2234.725 212.420 ;
      LAYER mcon ;
        RECT 2234.470 212.450 2234.640 213.300 ;
      LAYER met1 ;
        RECT 3369.800 1144.700 3369.940 1148.680 ;
        RECT 3369.520 1144.560 3369.940 1144.700 ;
        RECT 2234.455 226.920 2424.320 227.060 ;
        RECT 2234.455 226.800 2234.775 226.920 ;
        RECT 2424.180 215.420 2424.320 226.920 ;
        RECT 3369.520 218.060 3369.660 1144.560 ;
        RECT 2529.100 217.920 3369.660 218.060 ;
        RECT 2529.100 215.420 2529.240 217.920 ;
        RECT 2424.180 215.280 2529.240 215.420 ;
        RECT 2234.420 212.390 2234.680 213.360 ;
      LAYER via ;
        RECT 2234.485 226.800 2234.745 227.060 ;
        RECT 2234.420 212.450 2234.680 213.300 ;
      LAYER met2 ;
        RECT 2234.485 227.090 2234.625 232.485 ;
        RECT 2234.485 226.770 2234.745 227.090 ;
        RECT 2234.485 213.300 2234.625 226.770 ;
        RECT 2234.390 212.450 2234.710 213.300 ;
    END
  END mgmt_io_in_buf[13]
  PIN mgmt_io_in_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2226.055 213.300 2226.225 214.150 ;
        RECT 2226.895 213.300 2227.065 214.150 ;
        RECT 2227.735 213.300 2227.905 214.150 ;
        RECT 2228.575 213.300 2228.745 214.150 ;
        RECT 2226.055 213.130 2228.745 213.300 ;
        RECT 2228.490 212.590 2228.745 213.130 ;
        RECT 2226.055 212.420 2228.745 212.590 ;
        RECT 2226.055 211.940 2226.225 212.420 ;
        RECT 2226.895 211.940 2227.065 212.420 ;
        RECT 2227.735 211.940 2227.905 212.420 ;
        RECT 2228.575 211.940 2228.745 212.420 ;
      LAYER mcon ;
        RECT 2228.490 212.450 2228.660 213.300 ;
      LAYER met1 ;
        RECT 3368.680 1142.570 3368.820 1146.670 ;
        RECT 3368.400 1142.430 3368.820 1142.570 ;
        RECT 2228.475 227.760 2425.440 227.900 ;
        RECT 2228.475 227.640 2228.795 227.760 ;
        RECT 2425.300 215.980 2425.440 227.760 ;
        RECT 3368.400 218.900 3368.540 1142.430 ;
        RECT 2527.980 218.760 3368.540 218.900 ;
        RECT 2527.980 215.980 2528.120 218.760 ;
        RECT 2425.300 215.840 2528.120 215.980 ;
        RECT 2228.440 212.390 2228.700 213.360 ;
      LAYER via ;
        RECT 2228.505 227.640 2228.765 227.900 ;
        RECT 2228.440 212.450 2228.700 213.300 ;
      LAYER met2 ;
        RECT 2228.505 227.930 2228.645 232.485 ;
        RECT 2228.505 227.610 2228.765 227.930 ;
        RECT 2228.505 213.300 2228.645 227.610 ;
        RECT 2228.410 212.450 2228.730 213.300 ;
    END
  END mgmt_io_in_buf[14]
  PIN mgmt_io_in_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2220.075 213.300 2220.245 214.150 ;
        RECT 2220.915 213.300 2221.085 214.150 ;
        RECT 2221.755 213.300 2221.925 214.150 ;
        RECT 2222.595 213.300 2222.765 214.150 ;
        RECT 2220.075 213.130 2222.765 213.300 ;
        RECT 2222.510 212.590 2222.765 213.130 ;
        RECT 2220.075 212.420 2222.765 212.590 ;
        RECT 2220.075 211.940 2220.245 212.420 ;
        RECT 2220.915 211.940 2221.085 212.420 ;
        RECT 2221.755 211.940 2221.925 212.420 ;
        RECT 2222.595 211.940 2222.765 212.420 ;
      LAYER mcon ;
        RECT 2222.510 212.450 2222.680 213.300 ;
      LAYER met1 ;
        RECT 3367.560 1140.840 3367.700 1144.690 ;
        RECT 3367.280 1140.700 3367.700 1140.840 ;
        RECT 2222.495 228.600 2426.560 228.740 ;
        RECT 2222.495 228.480 2222.815 228.600 ;
        RECT 2426.420 216.540 2426.560 228.600 ;
        RECT 3367.280 219.740 3367.420 1140.700 ;
        RECT 2526.860 219.600 3367.420 219.740 ;
        RECT 2526.860 216.540 2527.000 219.600 ;
        RECT 2426.420 216.400 2527.000 216.540 ;
        RECT 2222.460 212.390 2222.720 213.360 ;
      LAYER via ;
        RECT 2222.525 228.480 2222.785 228.740 ;
        RECT 2222.460 212.450 2222.720 213.300 ;
      LAYER met2 ;
        RECT 2222.525 228.770 2222.665 232.485 ;
        RECT 2222.525 228.450 2222.785 228.770 ;
        RECT 2222.525 213.300 2222.665 228.450 ;
        RECT 2222.430 212.450 2222.750 213.300 ;
    END
  END mgmt_io_in_buf[15]
  PIN mgmt_io_in_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2214.095 213.300 2214.265 214.150 ;
        RECT 2214.935 213.300 2215.105 214.150 ;
        RECT 2215.775 213.300 2215.945 214.150 ;
        RECT 2216.615 213.300 2216.785 214.150 ;
        RECT 2214.095 213.130 2216.785 213.300 ;
        RECT 2216.530 212.590 2216.785 213.130 ;
        RECT 2214.095 212.420 2216.785 212.590 ;
        RECT 2214.095 211.940 2214.265 212.420 ;
        RECT 2214.935 211.940 2215.105 212.420 ;
        RECT 2215.775 211.940 2215.945 212.420 ;
        RECT 2216.615 211.940 2216.785 212.420 ;
      LAYER mcon ;
        RECT 2216.530 212.450 2216.700 213.300 ;
      LAYER met1 ;
        RECT 3366.440 1138.790 3366.580 1142.700 ;
        RECT 3366.160 1138.650 3366.580 1138.790 ;
        RECT 2216.515 229.440 2427.680 229.580 ;
        RECT 2216.515 229.320 2216.835 229.440 ;
        RECT 2427.540 217.100 2427.680 229.440 ;
        RECT 3366.160 220.580 3366.300 1138.650 ;
        RECT 2525.740 220.440 3366.300 220.580 ;
        RECT 2525.740 217.100 2525.880 220.440 ;
        RECT 2427.540 216.960 2525.880 217.100 ;
        RECT 2216.480 212.390 2216.740 213.360 ;
      LAYER via ;
        RECT 2216.545 229.320 2216.805 229.580 ;
        RECT 2216.480 212.450 2216.740 213.300 ;
      LAYER met2 ;
        RECT 2216.545 229.610 2216.685 232.485 ;
        RECT 2216.545 229.290 2216.805 229.610 ;
        RECT 2216.545 213.300 2216.685 229.290 ;
        RECT 2216.450 212.450 2216.770 213.300 ;
    END
  END mgmt_io_in_buf[16]
  PIN mgmt_io_in_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2208.115 213.300 2208.285 214.150 ;
        RECT 2208.955 213.300 2209.125 214.150 ;
        RECT 2209.795 213.300 2209.965 214.150 ;
        RECT 2210.635 213.300 2210.805 214.150 ;
        RECT 2208.115 213.130 2210.805 213.300 ;
        RECT 2210.550 212.590 2210.805 213.130 ;
        RECT 2208.115 212.420 2210.805 212.590 ;
        RECT 2208.115 211.940 2208.285 212.420 ;
        RECT 2208.955 211.940 2209.125 212.420 ;
        RECT 2209.795 211.940 2209.965 212.420 ;
        RECT 2210.635 211.940 2210.805 212.420 ;
      LAYER mcon ;
        RECT 2210.550 212.450 2210.720 213.300 ;
      LAYER met1 ;
        RECT 3365.320 1137.340 3365.460 1140.690 ;
        RECT 3365.040 1137.200 3365.460 1137.340 ;
        RECT 2210.535 230.280 2428.800 230.420 ;
        RECT 2210.535 230.160 2210.855 230.280 ;
        RECT 2428.660 217.660 2428.800 230.280 ;
        RECT 3365.040 221.420 3365.180 1137.200 ;
        RECT 2524.620 221.280 3365.180 221.420 ;
        RECT 2524.620 217.660 2524.760 221.280 ;
        RECT 2428.660 217.520 2524.760 217.660 ;
        RECT 2210.500 212.390 2210.760 213.360 ;
      LAYER via ;
        RECT 2210.565 230.160 2210.825 230.420 ;
        RECT 2210.500 212.450 2210.760 213.300 ;
      LAYER met2 ;
        RECT 2210.565 230.450 2210.705 232.485 ;
        RECT 2210.565 230.130 2210.825 230.450 ;
        RECT 2210.565 213.300 2210.705 230.130 ;
        RECT 2210.470 212.450 2210.790 213.300 ;
    END
  END mgmt_io_in_buf[17]
  PIN mgmt_io_in_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2202.135 213.300 2202.305 214.150 ;
        RECT 2202.975 213.300 2203.145 214.150 ;
        RECT 2203.815 213.300 2203.985 214.150 ;
        RECT 2204.655 213.300 2204.825 214.150 ;
        RECT 2202.135 213.130 2204.825 213.300 ;
        RECT 2204.570 212.590 2204.825 213.130 ;
        RECT 2202.135 212.420 2204.825 212.590 ;
        RECT 2202.135 211.940 2202.305 212.420 ;
        RECT 2202.975 211.940 2203.145 212.420 ;
        RECT 2203.815 211.940 2203.985 212.420 ;
        RECT 2204.655 211.940 2204.825 212.420 ;
      LAYER mcon ;
        RECT 2204.570 212.450 2204.740 213.300 ;
      LAYER met1 ;
        RECT 3364.200 1135.060 3364.340 1138.680 ;
        RECT 3363.920 1134.920 3364.340 1135.060 ;
        RECT 2204.555 231.120 2429.920 231.260 ;
        RECT 2204.555 231.000 2204.875 231.120 ;
        RECT 2429.780 218.220 2429.920 231.120 ;
        RECT 3363.920 222.260 3364.060 1134.920 ;
        RECT 2523.500 222.120 3364.060 222.260 ;
        RECT 2523.500 218.220 2523.640 222.120 ;
        RECT 2429.780 218.080 2523.640 218.220 ;
        RECT 2204.520 212.390 2204.780 213.360 ;
      LAYER via ;
        RECT 2204.585 231.000 2204.845 231.260 ;
        RECT 2204.520 212.450 2204.780 213.300 ;
      LAYER met2 ;
        RECT 2204.585 231.290 2204.725 232.485 ;
        RECT 2204.585 230.970 2204.845 231.290 ;
        RECT 2204.585 213.300 2204.725 230.970 ;
        RECT 2204.490 212.450 2204.810 213.300 ;
    END
  END mgmt_io_in_buf[18]
  PIN mgmt_io_in_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2196.155 213.300 2196.325 214.150 ;
        RECT 2196.995 213.300 2197.165 214.150 ;
        RECT 2197.835 213.300 2198.005 214.150 ;
        RECT 2198.675 213.300 2198.845 214.150 ;
        RECT 2196.155 213.130 2198.845 213.300 ;
        RECT 2198.590 212.590 2198.845 213.130 ;
        RECT 2196.155 212.420 2198.845 212.590 ;
        RECT 2196.155 211.940 2196.325 212.420 ;
        RECT 2196.995 211.940 2197.165 212.420 ;
        RECT 2197.835 211.940 2198.005 212.420 ;
        RECT 2198.675 211.940 2198.845 212.420 ;
      LAYER mcon ;
        RECT 2198.590 212.450 2198.760 213.300 ;
      LAYER met1 ;
        RECT 3363.080 1133.110 3363.220 1136.680 ;
        RECT 3362.800 1132.970 3363.220 1133.110 ;
        RECT 2198.575 231.960 2431.040 232.100 ;
        RECT 2198.575 231.840 2198.895 231.960 ;
        RECT 2430.900 218.780 2431.040 231.960 ;
        RECT 3362.800 223.100 3362.940 1132.970 ;
        RECT 2522.380 222.960 3362.940 223.100 ;
        RECT 2522.380 218.780 2522.520 222.960 ;
        RECT 2430.900 218.640 2522.520 218.780 ;
        RECT 2198.540 212.390 2198.800 213.360 ;
      LAYER via ;
        RECT 2198.605 231.840 2198.865 232.100 ;
        RECT 2198.540 212.450 2198.800 213.300 ;
      LAYER met2 ;
        RECT 2198.605 232.130 2198.745 232.485 ;
        RECT 2198.605 231.810 2198.865 232.130 ;
        RECT 2198.605 213.300 2198.745 231.810 ;
        RECT 2198.510 212.450 2198.830 213.300 ;
    END
  END mgmt_io_in_buf[19]
  PIN mgmt_io_in_buf[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2190.175 213.300 2190.345 214.150 ;
        RECT 2191.015 213.300 2191.185 214.150 ;
        RECT 2191.855 213.300 2192.025 214.150 ;
        RECT 2192.695 213.300 2192.865 214.150 ;
        RECT 2190.175 213.130 2192.865 213.300 ;
        RECT 2192.610 212.590 2192.865 213.130 ;
        RECT 2190.175 212.420 2192.865 212.590 ;
        RECT 2190.175 211.940 2190.345 212.420 ;
        RECT 2191.015 211.940 2191.185 212.420 ;
        RECT 2191.855 211.940 2192.025 212.420 ;
        RECT 2192.695 211.940 2192.865 212.420 ;
      LAYER mcon ;
        RECT 2192.610 212.450 2192.780 213.300 ;
      LAYER met1 ;
        RECT 3361.960 1130.930 3362.100 1134.710 ;
        RECT 3361.680 1130.790 3362.100 1130.930 ;
        RECT 2192.595 232.800 2432.160 232.940 ;
        RECT 2192.595 232.680 2192.915 232.800 ;
        RECT 2432.020 219.340 2432.160 232.800 ;
        RECT 3361.680 223.940 3361.820 1130.790 ;
        RECT 2521.260 223.800 3361.820 223.940 ;
        RECT 2521.260 219.340 2521.400 223.800 ;
        RECT 2432.020 219.200 2521.400 219.340 ;
        RECT 2192.560 212.390 2192.820 213.360 ;
      LAYER via ;
        RECT 2192.625 232.680 2192.885 232.940 ;
        RECT 2192.560 212.450 2192.820 213.300 ;
      LAYER met2 ;
        RECT 2192.625 232.970 2192.765 233.010 ;
        RECT 2192.625 232.650 2192.885 232.970 ;
        RECT 2192.625 213.300 2192.765 232.650 ;
        RECT 2192.530 212.450 2192.850 213.300 ;
    END
  END mgmt_io_in_buf[20]
  PIN mgmt_io_in_buf[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2184.195 213.300 2184.365 214.150 ;
        RECT 2185.035 213.300 2185.205 214.150 ;
        RECT 2185.875 213.300 2186.045 214.150 ;
        RECT 2186.715 213.300 2186.885 214.150 ;
        RECT 2184.195 213.130 2186.885 213.300 ;
        RECT 2186.630 212.590 2186.885 213.130 ;
        RECT 2184.195 212.420 2186.885 212.590 ;
        RECT 2184.195 211.940 2184.365 212.420 ;
        RECT 2185.035 211.940 2185.205 212.420 ;
        RECT 2185.875 211.940 2186.045 212.420 ;
        RECT 2186.715 211.940 2186.885 212.420 ;
      LAYER mcon ;
        RECT 2186.630 212.450 2186.800 213.300 ;
      LAYER met1 ;
        RECT 3360.840 1128.910 3360.980 1132.680 ;
        RECT 3360.560 1128.770 3360.980 1128.910 ;
        RECT 2186.615 233.640 2433.280 233.780 ;
        RECT 2186.615 233.520 2186.935 233.640 ;
        RECT 2433.140 219.900 2433.280 233.640 ;
        RECT 3360.560 224.780 3360.700 1128.770 ;
        RECT 2520.140 224.640 3360.700 224.780 ;
        RECT 2520.140 219.900 2520.280 224.640 ;
        RECT 2433.140 219.760 2520.280 219.900 ;
        RECT 2186.580 212.390 2186.840 213.360 ;
      LAYER via ;
        RECT 2186.645 233.520 2186.905 233.780 ;
        RECT 2186.580 212.450 2186.840 213.300 ;
      LAYER met2 ;
        RECT 2186.645 233.810 2186.785 233.870 ;
        RECT 2186.645 233.490 2186.905 233.810 ;
        RECT 2186.645 213.300 2186.785 233.490 ;
        RECT 2186.550 212.450 2186.870 213.300 ;
    END
  END mgmt_io_in_buf[21]
  PIN mgmt_io_in_buf[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2178.215 213.300 2178.385 214.150 ;
        RECT 2179.055 213.300 2179.225 214.150 ;
        RECT 2179.895 213.300 2180.065 214.150 ;
        RECT 2180.735 213.300 2180.905 214.150 ;
        RECT 2178.215 213.130 2180.905 213.300 ;
        RECT 2180.650 212.590 2180.905 213.130 ;
        RECT 2178.215 212.420 2180.905 212.590 ;
        RECT 2178.215 211.940 2178.385 212.420 ;
        RECT 2179.055 211.940 2179.225 212.420 ;
        RECT 2179.895 211.940 2180.065 212.420 ;
        RECT 2180.735 211.940 2180.905 212.420 ;
      LAYER mcon ;
        RECT 2180.650 212.450 2180.820 213.300 ;
      LAYER met1 ;
        RECT 3359.720 1127.010 3359.860 1130.700 ;
        RECT 3359.440 1126.870 3359.860 1127.010 ;
        RECT 2180.635 234.480 2434.400 234.620 ;
        RECT 2180.635 234.360 2180.955 234.480 ;
        RECT 2434.260 220.460 2434.400 234.480 ;
        RECT 3359.440 225.620 3359.580 1126.870 ;
        RECT 2519.020 225.480 3359.580 225.620 ;
        RECT 2519.020 220.460 2519.160 225.480 ;
        RECT 2434.260 220.320 2519.160 220.460 ;
        RECT 2180.600 212.390 2180.860 213.360 ;
      LAYER via ;
        RECT 2180.665 234.360 2180.925 234.620 ;
        RECT 2180.600 212.450 2180.860 213.300 ;
      LAYER met2 ;
        RECT 2180.665 234.650 2180.805 234.705 ;
        RECT 2180.665 234.330 2180.925 234.650 ;
        RECT 2180.665 213.300 2180.805 234.330 ;
        RECT 2180.570 212.450 2180.890 213.300 ;
    END
  END mgmt_io_in_buf[22]
  PIN mgmt_io_in_buf[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2172.235 213.300 2172.405 214.150 ;
        RECT 2173.075 213.300 2173.245 214.150 ;
        RECT 2173.915 213.300 2174.085 214.150 ;
        RECT 2174.755 213.300 2174.925 214.150 ;
        RECT 2172.235 213.130 2174.925 213.300 ;
        RECT 2174.670 212.590 2174.925 213.130 ;
        RECT 2172.235 212.420 2174.925 212.590 ;
        RECT 2172.235 211.940 2172.405 212.420 ;
        RECT 2173.075 211.940 2173.245 212.420 ;
        RECT 2173.915 211.940 2174.085 212.420 ;
        RECT 2174.755 211.940 2174.925 212.420 ;
      LAYER mcon ;
        RECT 2174.670 212.450 2174.840 213.300 ;
      LAYER met1 ;
        RECT 3358.600 1125.030 3358.740 1128.720 ;
        RECT 3358.320 1124.890 3358.740 1125.030 ;
        RECT 2174.655 235.320 2435.520 235.460 ;
        RECT 2174.655 235.200 2174.975 235.320 ;
        RECT 2435.380 221.020 2435.520 235.320 ;
        RECT 3358.320 226.460 3358.460 1124.890 ;
        RECT 2517.900 226.320 3358.460 226.460 ;
        RECT 2517.900 221.020 2518.040 226.320 ;
        RECT 2435.380 220.880 2518.040 221.020 ;
        RECT 2174.620 212.390 2174.880 213.360 ;
      LAYER via ;
        RECT 2174.685 235.200 2174.945 235.460 ;
        RECT 2174.620 212.450 2174.880 213.300 ;
      LAYER met2 ;
        RECT 2174.685 235.490 2174.825 235.530 ;
        RECT 2174.685 235.170 2174.945 235.490 ;
        RECT 2174.685 213.300 2174.825 235.170 ;
        RECT 2174.590 212.450 2174.910 213.300 ;
    END
  END mgmt_io_in_buf[23]
  PIN mgmt_io_in_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2166.255 213.300 2166.425 214.150 ;
        RECT 2167.095 213.300 2167.265 214.150 ;
        RECT 2167.935 213.300 2168.105 214.150 ;
        RECT 2168.775 213.300 2168.945 214.150 ;
        RECT 2166.255 213.130 2168.945 213.300 ;
        RECT 2168.690 212.590 2168.945 213.130 ;
        RECT 2166.255 212.420 2168.945 212.590 ;
        RECT 2166.255 211.940 2166.425 212.420 ;
        RECT 2167.095 211.940 2167.265 212.420 ;
        RECT 2167.935 211.940 2168.105 212.420 ;
        RECT 2168.775 211.940 2168.945 212.420 ;
      LAYER mcon ;
        RECT 2168.690 212.450 2168.860 213.300 ;
      LAYER met1 ;
        RECT 3357.480 1123.150 3357.620 1126.740 ;
        RECT 3357.200 1123.010 3357.620 1123.150 ;
        RECT 2168.675 236.160 2436.640 236.300 ;
        RECT 2168.675 236.040 2168.995 236.160 ;
        RECT 2436.500 221.580 2436.640 236.160 ;
        RECT 3357.200 227.300 3357.340 1123.010 ;
        RECT 2516.780 227.160 3357.340 227.300 ;
        RECT 2516.780 221.580 2516.920 227.160 ;
        RECT 2436.500 221.440 2516.920 221.580 ;
        RECT 2168.640 212.390 2168.900 213.360 ;
      LAYER via ;
        RECT 2168.705 236.040 2168.965 236.300 ;
        RECT 2168.640 212.450 2168.900 213.300 ;
      LAYER met2 ;
        RECT 2168.705 236.330 2168.845 236.400 ;
        RECT 2168.705 236.010 2168.965 236.330 ;
        RECT 2168.705 213.300 2168.845 236.010 ;
        RECT 2168.610 212.450 2168.930 213.300 ;
    END
  END mgmt_io_in_buf[24]
  PIN mgmt_io_in_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2160.275 213.300 2160.445 214.150 ;
        RECT 2161.115 213.300 2161.285 214.150 ;
        RECT 2161.955 213.300 2162.125 214.150 ;
        RECT 2162.795 213.300 2162.965 214.150 ;
        RECT 2160.275 213.130 2162.965 213.300 ;
        RECT 2162.710 212.590 2162.965 213.130 ;
        RECT 2160.275 212.420 2162.965 212.590 ;
        RECT 2160.275 211.940 2160.445 212.420 ;
        RECT 2161.115 211.940 2161.285 212.420 ;
        RECT 2161.955 211.940 2162.125 212.420 ;
        RECT 2162.795 211.940 2162.965 212.420 ;
      LAYER mcon ;
        RECT 2162.710 212.450 2162.880 213.300 ;
      LAYER met1 ;
        RECT 3356.360 1121.090 3356.500 1124.690 ;
        RECT 3356.080 1120.950 3356.500 1121.090 ;
        RECT 2162.695 237.000 2437.760 237.140 ;
        RECT 2162.695 236.880 2163.015 237.000 ;
        RECT 2437.620 222.140 2437.760 237.000 ;
        RECT 3356.080 228.140 3356.220 1120.950 ;
        RECT 2515.660 228.000 3356.220 228.140 ;
        RECT 2515.660 222.140 2515.800 228.000 ;
        RECT 2437.620 222.000 2515.800 222.140 ;
        RECT 2162.660 212.390 2162.920 213.360 ;
      LAYER via ;
        RECT 2162.725 236.880 2162.985 237.140 ;
        RECT 2162.660 212.450 2162.920 213.300 ;
      LAYER met2 ;
        RECT 2162.725 237.170 2162.865 237.225 ;
        RECT 2162.725 236.850 2162.985 237.170 ;
        RECT 2162.725 213.300 2162.865 236.850 ;
        RECT 2162.630 212.450 2162.950 213.300 ;
    END
  END mgmt_io_in_buf[25]
  PIN mgmt_io_in_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2154.295 213.300 2154.465 214.150 ;
        RECT 2155.135 213.300 2155.305 214.150 ;
        RECT 2155.975 213.300 2156.145 214.150 ;
        RECT 2156.815 213.300 2156.985 214.150 ;
        RECT 2154.295 213.130 2156.985 213.300 ;
        RECT 2156.730 212.590 2156.985 213.130 ;
        RECT 2154.295 212.420 2156.985 212.590 ;
        RECT 2154.295 211.940 2154.465 212.420 ;
        RECT 2155.135 211.940 2155.305 212.420 ;
        RECT 2155.975 211.940 2156.145 212.420 ;
        RECT 2156.815 211.940 2156.985 212.420 ;
      LAYER mcon ;
        RECT 2156.730 212.450 2156.900 213.300 ;
      LAYER met1 ;
        RECT 3355.240 1118.490 3355.380 1122.730 ;
        RECT 3354.960 1118.350 3355.380 1118.490 ;
        RECT 2156.715 237.840 2438.880 237.980 ;
        RECT 2156.715 237.720 2157.035 237.840 ;
        RECT 2438.740 222.700 2438.880 237.840 ;
        RECT 3354.960 228.980 3355.100 1118.350 ;
        RECT 2514.540 228.840 3355.100 228.980 ;
        RECT 2514.540 222.700 2514.680 228.840 ;
        RECT 2438.740 222.560 2514.680 222.700 ;
        RECT 2156.680 212.390 2156.940 213.360 ;
      LAYER via ;
        RECT 2156.745 237.720 2157.005 237.980 ;
        RECT 2156.680 212.450 2156.940 213.300 ;
      LAYER met2 ;
        RECT 2156.745 238.010 2156.885 238.085 ;
        RECT 2156.745 237.690 2157.005 238.010 ;
        RECT 2156.745 213.300 2156.885 237.690 ;
        RECT 2156.650 212.450 2156.970 213.300 ;
    END
  END mgmt_io_in_buf[26]
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 2082.975 4987.615 2083.145 4987.785 ;
        RECT 2083.435 4987.615 2083.605 4987.785 ;
        RECT 2083.895 4987.615 2084.065 4987.785 ;
        RECT 2084.355 4987.615 2084.525 4987.785 ;
        RECT 2084.815 4987.615 2084.985 4987.785 ;
        RECT 2085.275 4987.615 2085.445 4987.785 ;
        RECT 2085.735 4987.615 2085.905 4987.785 ;
        RECT 2086.195 4987.615 2086.365 4987.785 ;
        RECT 2086.655 4987.615 2086.825 4987.785 ;
        RECT 2087.115 4987.615 2087.285 4987.785 ;
        RECT 2087.575 4987.615 2087.745 4987.785 ;
        RECT 2088.035 4987.615 2088.205 4987.785 ;
        RECT 2088.495 4987.615 2088.665 4987.785 ;
        RECT 2088.955 4987.615 2089.125 4987.785 ;
        RECT 2082.975 4982.175 2083.145 4982.345 ;
        RECT 2083.435 4982.175 2083.605 4982.345 ;
        RECT 2083.895 4982.175 2084.065 4982.345 ;
        RECT 2084.355 4982.175 2084.525 4982.345 ;
        RECT 2084.815 4982.175 2084.985 4982.345 ;
        RECT 2085.275 4982.175 2085.445 4982.345 ;
        RECT 2085.735 4982.175 2085.905 4982.345 ;
        RECT 2086.195 4982.175 2086.365 4982.345 ;
        RECT 2086.655 4982.175 2086.825 4982.345 ;
        RECT 2087.115 4982.175 2087.285 4982.345 ;
        RECT 2087.575 4982.175 2087.745 4982.345 ;
        RECT 2088.035 4982.175 2088.205 4982.345 ;
        RECT 2088.495 4982.175 2088.665 4982.345 ;
        RECT 2088.955 4982.175 2089.125 4982.345 ;
      LAYER met1 ;
        RECT 2082.830 4987.460 2089.270 4987.940 ;
        RECT 2082.830 4982.020 2089.270 4982.500 ;
      LAYER via ;
        RECT 2085.135 4987.535 2086.920 4987.835 ;
        RECT 2085.135 4982.125 2086.920 4982.425 ;
      LAYER met2 ;
        RECT 2085.095 4987.490 2086.960 4987.920 ;
        RECT 2085.095 4982.065 2086.960 4982.495 ;
      LAYER via2 ;
        RECT 2085.135 4987.535 2086.920 4987.835 ;
        RECT 2085.135 4982.125 2086.920 4982.425 ;
      LAYER met3 ;
        RECT 2085.090 4982.050 2086.955 4989.575 ;
    END
    PORT
      LAYER li1 ;
        RECT 834.795 4985.990 834.965 4986.160 ;
        RECT 835.255 4985.990 835.425 4986.160 ;
        RECT 835.715 4985.990 835.885 4986.160 ;
        RECT 836.175 4985.990 836.345 4986.160 ;
        RECT 836.635 4985.990 836.805 4986.160 ;
        RECT 837.095 4985.990 837.265 4986.160 ;
        RECT 837.555 4985.990 837.725 4986.160 ;
        RECT 838.015 4985.990 838.185 4986.160 ;
        RECT 838.475 4985.990 838.645 4986.160 ;
        RECT 838.935 4985.990 839.105 4986.160 ;
        RECT 839.395 4985.990 839.565 4986.160 ;
        RECT 839.855 4985.990 840.025 4986.160 ;
        RECT 840.315 4985.990 840.485 4986.160 ;
        RECT 840.775 4985.990 840.945 4986.160 ;
        RECT 841.235 4985.990 841.405 4986.160 ;
        RECT 841.695 4985.990 841.865 4986.160 ;
        RECT 842.155 4985.990 842.325 4986.160 ;
        RECT 842.615 4985.990 842.785 4986.160 ;
        RECT 843.075 4985.990 843.245 4986.160 ;
        RECT 843.535 4985.990 843.705 4986.160 ;
        RECT 843.995 4985.990 844.165 4986.160 ;
        RECT 844.455 4985.990 844.625 4986.160 ;
        RECT 844.915 4985.990 845.085 4986.160 ;
        RECT 845.375 4985.990 845.545 4986.160 ;
        RECT 845.835 4985.990 846.005 4986.160 ;
        RECT 846.295 4985.990 846.465 4986.160 ;
        RECT 846.755 4985.990 846.925 4986.160 ;
        RECT 847.215 4985.990 847.385 4986.160 ;
        RECT 847.675 4985.990 847.845 4986.160 ;
        RECT 848.135 4985.990 848.305 4986.160 ;
        RECT 848.595 4985.990 848.765 4986.160 ;
        RECT 849.055 4985.990 849.225 4986.160 ;
        RECT 849.515 4985.990 849.685 4986.160 ;
        RECT 849.975 4985.990 850.145 4986.160 ;
        RECT 850.435 4985.990 850.605 4986.160 ;
        RECT 850.895 4985.990 851.065 4986.160 ;
        RECT 851.355 4985.990 851.525 4986.160 ;
        RECT 851.815 4985.990 851.985 4986.160 ;
        RECT 852.275 4985.990 852.445 4986.160 ;
        RECT 852.735 4985.990 852.905 4986.160 ;
        RECT 834.795 4980.550 834.965 4980.720 ;
        RECT 835.255 4980.550 835.425 4980.720 ;
        RECT 835.715 4980.550 835.885 4980.720 ;
        RECT 836.175 4980.550 836.345 4980.720 ;
        RECT 836.635 4980.550 836.805 4980.720 ;
        RECT 837.095 4980.550 837.265 4980.720 ;
        RECT 837.555 4980.550 837.725 4980.720 ;
        RECT 838.015 4980.550 838.185 4980.720 ;
        RECT 838.475 4980.550 838.645 4980.720 ;
        RECT 838.935 4980.550 839.105 4980.720 ;
        RECT 839.395 4980.550 839.565 4980.720 ;
        RECT 839.855 4980.550 840.025 4980.720 ;
        RECT 840.315 4980.550 840.485 4980.720 ;
        RECT 840.775 4980.550 840.945 4980.720 ;
        RECT 841.235 4980.550 841.405 4980.720 ;
        RECT 841.695 4980.550 841.865 4980.720 ;
        RECT 842.155 4980.550 842.325 4980.720 ;
        RECT 842.615 4980.550 842.785 4980.720 ;
        RECT 843.075 4980.550 843.245 4980.720 ;
        RECT 843.535 4980.550 843.705 4980.720 ;
        RECT 843.995 4980.550 844.165 4980.720 ;
        RECT 844.455 4980.550 844.625 4980.720 ;
        RECT 844.915 4980.550 845.085 4980.720 ;
        RECT 845.375 4980.550 845.545 4980.720 ;
        RECT 845.835 4980.550 846.005 4980.720 ;
        RECT 846.295 4980.550 846.465 4980.720 ;
        RECT 846.755 4980.550 846.925 4980.720 ;
        RECT 847.215 4980.550 847.385 4980.720 ;
        RECT 847.675 4980.550 847.845 4980.720 ;
        RECT 848.135 4980.550 848.305 4980.720 ;
        RECT 848.595 4980.550 848.765 4980.720 ;
        RECT 849.055 4980.550 849.225 4980.720 ;
        RECT 849.515 4980.550 849.685 4980.720 ;
        RECT 849.975 4980.550 850.145 4980.720 ;
        RECT 850.435 4980.550 850.605 4980.720 ;
        RECT 850.895 4980.550 851.065 4980.720 ;
        RECT 851.355 4980.550 851.525 4980.720 ;
        RECT 851.815 4980.550 851.985 4980.720 ;
        RECT 852.275 4980.550 852.445 4980.720 ;
        RECT 852.735 4980.550 852.905 4980.720 ;
      LAYER met1 ;
        RECT 834.650 4985.835 853.050 4986.315 ;
        RECT 834.650 4980.395 853.050 4980.875 ;
      LAYER via ;
        RECT 842.950 4985.890 844.735 4986.190 ;
        RECT 842.950 4980.480 844.735 4980.780 ;
      LAYER met2 ;
        RECT 842.910 4985.845 844.775 4986.275 ;
        RECT 842.910 4980.420 844.775 4980.850 ;
      LAYER via2 ;
        RECT 842.950 4985.890 844.735 4986.190 ;
        RECT 842.950 4980.480 844.735 4980.780 ;
      LAYER met3 ;
        RECT 842.905 4980.405 844.770 4987.930 ;
    END
    PORT
      LAYER li1 ;
        RECT 3309.980 4987.205 3310.150 4987.375 ;
        RECT 3310.440 4987.205 3310.610 4987.375 ;
        RECT 3310.900 4987.205 3311.070 4987.375 ;
        RECT 3311.360 4987.205 3311.530 4987.375 ;
        RECT 3311.820 4987.205 3311.990 4987.375 ;
        RECT 3312.280 4987.205 3312.450 4987.375 ;
        RECT 3312.740 4987.205 3312.910 4987.375 ;
        RECT 3313.200 4987.205 3313.370 4987.375 ;
        RECT 3313.660 4987.205 3313.830 4987.375 ;
        RECT 3314.120 4987.205 3314.290 4987.375 ;
        RECT 3314.580 4987.205 3314.750 4987.375 ;
        RECT 3315.040 4987.205 3315.210 4987.375 ;
        RECT 3315.500 4987.205 3315.670 4987.375 ;
        RECT 3315.960 4987.205 3316.130 4987.375 ;
        RECT 3316.420 4987.205 3316.590 4987.375 ;
        RECT 3316.880 4987.205 3317.050 4987.375 ;
        RECT 3317.340 4987.205 3317.510 4987.375 ;
        RECT 3317.800 4987.205 3317.970 4987.375 ;
        RECT 3318.260 4987.205 3318.430 4987.375 ;
        RECT 3318.720 4987.205 3318.890 4987.375 ;
        RECT 3319.180 4987.205 3319.350 4987.375 ;
        RECT 3319.640 4987.205 3319.810 4987.375 ;
        RECT 3320.100 4987.205 3320.270 4987.375 ;
        RECT 3320.560 4987.205 3320.730 4987.375 ;
        RECT 3321.020 4987.205 3321.190 4987.375 ;
        RECT 3321.480 4987.205 3321.650 4987.375 ;
        RECT 3321.940 4987.205 3322.110 4987.375 ;
        RECT 3322.400 4987.205 3322.570 4987.375 ;
        RECT 3322.860 4987.205 3323.030 4987.375 ;
        RECT 3323.320 4987.205 3323.490 4987.375 ;
        RECT 3323.780 4987.205 3323.950 4987.375 ;
        RECT 3324.240 4987.205 3324.410 4987.375 ;
        RECT 3324.700 4987.205 3324.870 4987.375 ;
        RECT 3325.160 4987.205 3325.330 4987.375 ;
        RECT 3325.620 4987.205 3325.790 4987.375 ;
        RECT 3326.080 4987.205 3326.250 4987.375 ;
        RECT 3326.540 4987.205 3326.710 4987.375 ;
        RECT 3327.000 4987.205 3327.170 4987.375 ;
        RECT 3327.460 4987.205 3327.630 4987.375 ;
        RECT 3327.920 4987.205 3328.090 4987.375 ;
        RECT 3328.380 4987.205 3328.550 4987.375 ;
        RECT 3328.840 4987.205 3329.010 4987.375 ;
        RECT 3329.300 4987.205 3329.470 4987.375 ;
        RECT 3329.760 4987.205 3329.930 4987.375 ;
        RECT 3330.220 4987.205 3330.390 4987.375 ;
        RECT 3330.680 4987.205 3330.850 4987.375 ;
        RECT 3331.140 4987.205 3331.310 4987.375 ;
        RECT 3331.600 4987.205 3331.770 4987.375 ;
        RECT 3332.060 4987.205 3332.230 4987.375 ;
        RECT 3332.520 4987.205 3332.690 4987.375 ;
        RECT 3332.980 4987.205 3333.150 4987.375 ;
        RECT 3333.440 4987.205 3333.610 4987.375 ;
        RECT 3333.900 4987.205 3334.070 4987.375 ;
        RECT 3309.980 4981.765 3310.150 4981.935 ;
      LAYER li1 ;
        RECT 3310.295 4981.765 3315.500 4981.935 ;
        RECT 3315.670 4981.765 3315.815 4981.935 ;
      LAYER li1 ;
        RECT 3315.960 4981.765 3316.130 4981.935 ;
        RECT 3316.420 4981.765 3316.590 4981.935 ;
        RECT 3316.880 4981.765 3317.050 4981.935 ;
        RECT 3317.340 4981.765 3317.510 4981.935 ;
        RECT 3317.800 4981.765 3317.970 4981.935 ;
        RECT 3318.260 4981.765 3318.430 4981.935 ;
        RECT 3318.720 4981.765 3318.890 4981.935 ;
        RECT 3319.180 4981.765 3319.350 4981.935 ;
        RECT 3319.640 4981.765 3319.810 4981.935 ;
        RECT 3320.100 4981.765 3320.270 4981.935 ;
        RECT 3320.560 4981.765 3320.730 4981.935 ;
        RECT 3321.020 4981.765 3321.190 4981.935 ;
        RECT 3321.480 4981.765 3321.650 4981.935 ;
        RECT 3321.940 4981.765 3322.110 4981.935 ;
        RECT 3322.400 4981.765 3322.570 4981.935 ;
        RECT 3322.860 4981.765 3323.030 4981.935 ;
        RECT 3323.320 4981.765 3323.490 4981.935 ;
        RECT 3323.780 4981.765 3323.950 4981.935 ;
        RECT 3324.240 4981.765 3324.410 4981.935 ;
        RECT 3324.700 4981.765 3324.870 4981.935 ;
        RECT 3325.160 4981.765 3325.330 4981.935 ;
        RECT 3325.620 4981.765 3325.790 4981.935 ;
        RECT 3326.080 4981.765 3326.250 4981.935 ;
        RECT 3326.540 4981.765 3326.710 4981.935 ;
        RECT 3327.000 4981.765 3327.170 4981.935 ;
        RECT 3327.460 4981.765 3327.630 4981.935 ;
        RECT 3327.920 4981.765 3328.090 4981.935 ;
        RECT 3328.380 4981.765 3328.550 4981.935 ;
        RECT 3328.840 4981.765 3329.010 4981.935 ;
        RECT 3329.300 4981.765 3329.470 4981.935 ;
        RECT 3329.760 4981.765 3329.930 4981.935 ;
        RECT 3330.220 4981.765 3330.390 4981.935 ;
        RECT 3330.680 4981.765 3330.850 4981.935 ;
        RECT 3331.140 4981.765 3331.310 4981.935 ;
        RECT 3331.600 4981.765 3331.770 4981.935 ;
        RECT 3332.060 4981.765 3332.230 4981.935 ;
        RECT 3332.520 4981.765 3332.690 4981.935 ;
        RECT 3332.980 4981.765 3333.150 4981.935 ;
        RECT 3333.440 4981.765 3333.610 4981.935 ;
        RECT 3333.900 4981.765 3334.070 4981.935 ;
      LAYER li1 ;
        RECT 3310.385 4981.220 3315.730 4981.765 ;
        RECT 3313.805 4980.390 3314.145 4981.220 ;
      LAYER mcon ;
        RECT 3310.440 4981.765 3310.610 4981.935 ;
        RECT 3310.900 4981.765 3311.070 4981.935 ;
        RECT 3311.360 4981.765 3311.530 4981.935 ;
        RECT 3311.820 4981.765 3311.990 4981.935 ;
        RECT 3312.280 4981.765 3312.450 4981.935 ;
        RECT 3312.740 4981.765 3312.910 4981.935 ;
        RECT 3313.200 4981.765 3313.370 4981.935 ;
        RECT 3313.660 4981.765 3313.830 4981.935 ;
        RECT 3314.120 4981.765 3314.290 4981.935 ;
        RECT 3314.580 4981.765 3314.750 4981.935 ;
        RECT 3315.040 4981.765 3315.210 4981.935 ;
      LAYER met1 ;
        RECT 3309.835 4987.050 3334.215 4987.530 ;
        RECT 3309.835 4981.610 3334.215 4982.090 ;
      LAYER via ;
        RECT 3318.185 4987.125 3319.970 4987.425 ;
        RECT 3318.185 4981.715 3319.970 4982.015 ;
      LAYER met2 ;
        RECT 3318.145 4987.080 3320.010 4987.510 ;
        RECT 3318.145 4981.655 3320.010 4982.085 ;
      LAYER via2 ;
        RECT 3318.185 4987.125 3319.970 4987.425 ;
        RECT 3318.185 4981.715 3319.970 4982.015 ;
      LAYER met3 ;
        RECT 3318.140 4981.640 3320.005 4989.165 ;
    END
    PORT
      LAYER li1 ;
        RECT 3380.500 2267.965 3380.670 2268.135 ;
        RECT 3385.940 2267.965 3386.110 2268.135 ;
        RECT 3380.500 2267.505 3380.670 2267.675 ;
        RECT 3385.940 2267.505 3386.110 2267.675 ;
        RECT 3380.500 2267.045 3380.670 2267.215 ;
        RECT 3385.940 2267.045 3386.110 2267.215 ;
        RECT 3380.500 2266.585 3380.670 2266.755 ;
        RECT 3385.940 2266.585 3386.110 2266.755 ;
        RECT 3380.500 2266.125 3380.670 2266.295 ;
        RECT 3385.940 2266.125 3386.110 2266.295 ;
        RECT 3380.500 2265.665 3380.670 2265.835 ;
        RECT 3385.940 2265.665 3386.110 2265.835 ;
        RECT 3380.500 2265.205 3380.670 2265.375 ;
        RECT 3385.940 2265.205 3386.110 2265.375 ;
        RECT 3380.500 2264.745 3380.670 2264.915 ;
        RECT 3385.940 2264.745 3386.110 2264.915 ;
        RECT 3380.500 2264.285 3380.670 2264.455 ;
        RECT 3385.940 2264.285 3386.110 2264.455 ;
        RECT 3380.500 2263.825 3380.670 2263.995 ;
        RECT 3385.940 2263.825 3386.110 2263.995 ;
        RECT 3380.500 2263.365 3380.670 2263.535 ;
        RECT 3385.940 2263.365 3386.110 2263.535 ;
        RECT 3380.500 2262.905 3380.670 2263.075 ;
        RECT 3385.940 2262.905 3386.110 2263.075 ;
        RECT 3380.500 2262.445 3380.670 2262.615 ;
        RECT 3385.940 2262.445 3386.110 2262.615 ;
        RECT 3380.500 2261.985 3380.670 2262.155 ;
        RECT 3385.940 2261.985 3386.110 2262.155 ;
        RECT 3380.500 2261.525 3380.670 2261.695 ;
        RECT 3385.940 2261.525 3386.110 2261.695 ;
        RECT 3380.500 2261.065 3380.670 2261.235 ;
        RECT 3385.940 2261.065 3386.110 2261.235 ;
        RECT 3380.500 2260.605 3380.670 2260.775 ;
        RECT 3385.940 2260.605 3386.110 2260.775 ;
        RECT 3380.500 2260.145 3380.670 2260.315 ;
        RECT 3385.940 2260.145 3386.110 2260.315 ;
        RECT 3380.500 2259.685 3380.670 2259.855 ;
        RECT 3385.940 2259.685 3386.110 2259.855 ;
        RECT 3380.500 2259.225 3380.670 2259.395 ;
        RECT 3385.940 2259.225 3386.110 2259.395 ;
        RECT 3380.500 2258.765 3380.670 2258.935 ;
        RECT 3385.940 2258.765 3386.110 2258.935 ;
        RECT 3380.500 2258.305 3380.670 2258.475 ;
        RECT 3385.940 2258.305 3386.110 2258.475 ;
        RECT 3380.500 2257.845 3380.670 2258.015 ;
        RECT 3385.940 2257.845 3386.110 2258.015 ;
        RECT 3380.500 2257.385 3380.670 2257.555 ;
        RECT 3385.940 2257.385 3386.110 2257.555 ;
        RECT 3380.500 2256.925 3380.670 2257.095 ;
        RECT 3385.940 2256.925 3386.110 2257.095 ;
        RECT 3380.500 2256.465 3380.670 2256.635 ;
        RECT 3385.940 2256.465 3386.110 2256.635 ;
        RECT 3380.500 2256.005 3380.670 2256.175 ;
        RECT 3385.940 2256.005 3386.110 2256.175 ;
        RECT 3380.500 2255.545 3380.670 2255.715 ;
        RECT 3385.940 2255.545 3386.110 2255.715 ;
        RECT 3380.500 2255.085 3380.670 2255.255 ;
        RECT 3385.940 2255.085 3386.110 2255.255 ;
        RECT 3380.500 2254.625 3380.670 2254.795 ;
        RECT 3385.940 2254.625 3386.110 2254.795 ;
        RECT 3380.500 2254.165 3380.670 2254.335 ;
        RECT 3385.940 2254.165 3386.110 2254.335 ;
        RECT 3380.500 2253.705 3380.670 2253.875 ;
        RECT 3385.940 2253.705 3386.110 2253.875 ;
        RECT 3380.500 2253.245 3380.670 2253.415 ;
        RECT 3385.940 2253.245 3386.110 2253.415 ;
        RECT 3380.500 2252.785 3380.670 2252.955 ;
        RECT 3385.940 2252.785 3386.110 2252.955 ;
        RECT 3380.500 2252.325 3380.670 2252.495 ;
        RECT 3385.940 2252.325 3386.110 2252.495 ;
        RECT 3380.500 2251.865 3380.670 2252.035 ;
        RECT 3385.940 2251.865 3386.110 2252.035 ;
        RECT 3380.500 2251.405 3380.670 2251.575 ;
        RECT 3385.940 2251.405 3386.110 2251.575 ;
        RECT 3380.500 2250.945 3380.670 2251.115 ;
        RECT 3385.940 2250.945 3386.110 2251.115 ;
        RECT 3380.500 2250.485 3380.670 2250.655 ;
        RECT 3385.940 2250.485 3386.110 2250.655 ;
        RECT 3380.500 2250.025 3380.670 2250.195 ;
        RECT 3385.940 2250.025 3386.110 2250.195 ;
        RECT 3380.500 2249.565 3380.670 2249.735 ;
        RECT 3385.940 2249.565 3386.110 2249.735 ;
        RECT 3380.500 2249.105 3380.670 2249.275 ;
        RECT 3385.940 2249.105 3386.110 2249.275 ;
        RECT 3380.500 2248.645 3380.670 2248.815 ;
        RECT 3385.940 2248.645 3386.110 2248.815 ;
        RECT 3380.500 2248.185 3380.670 2248.355 ;
        RECT 3385.940 2248.185 3386.110 2248.355 ;
        RECT 3380.500 2247.725 3380.670 2247.895 ;
        RECT 3385.940 2247.725 3386.110 2247.895 ;
        RECT 3380.500 2247.265 3380.670 2247.435 ;
        RECT 3385.940 2247.265 3386.110 2247.435 ;
        RECT 3380.500 2246.805 3380.670 2246.975 ;
        RECT 3385.940 2246.805 3386.110 2246.975 ;
        RECT 3380.500 2246.345 3380.670 2246.515 ;
        RECT 3385.940 2246.345 3386.110 2246.515 ;
        RECT 3380.500 2245.885 3380.670 2246.055 ;
        RECT 3385.940 2245.885 3386.110 2246.055 ;
        RECT 3380.500 2245.425 3380.670 2245.595 ;
        RECT 3385.940 2245.425 3386.110 2245.595 ;
        RECT 3380.500 2244.965 3380.670 2245.135 ;
        RECT 3385.940 2244.965 3386.110 2245.135 ;
        RECT 3380.500 2244.505 3380.670 2244.675 ;
        RECT 3385.940 2244.505 3386.110 2244.675 ;
        RECT 3380.500 2244.045 3380.670 2244.215 ;
        RECT 3385.940 2244.045 3386.110 2244.215 ;
        RECT 3380.500 2243.585 3380.670 2243.755 ;
        RECT 3385.940 2243.585 3386.110 2243.755 ;
        RECT 3380.500 2243.125 3380.670 2243.295 ;
        RECT 3385.940 2243.125 3386.110 2243.295 ;
        RECT 3380.500 2242.665 3380.670 2242.835 ;
        RECT 3385.940 2242.665 3386.110 2242.835 ;
        RECT 3380.500 2242.205 3380.670 2242.375 ;
        RECT 3385.940 2242.205 3386.110 2242.375 ;
        RECT 3380.500 2241.745 3380.670 2241.915 ;
        RECT 3385.940 2241.745 3386.110 2241.915 ;
        RECT 3380.500 2241.285 3380.670 2241.455 ;
        RECT 3385.940 2241.285 3386.110 2241.455 ;
        RECT 3380.500 2240.825 3380.670 2240.995 ;
        RECT 3385.940 2240.825 3386.110 2240.995 ;
        RECT 3380.500 2240.365 3380.670 2240.535 ;
        RECT 3385.940 2240.365 3386.110 2240.535 ;
        RECT 3380.500 2239.905 3380.670 2240.075 ;
        RECT 3385.940 2239.905 3386.110 2240.075 ;
        RECT 3380.500 2239.445 3380.670 2239.615 ;
        RECT 3385.940 2239.445 3386.110 2239.615 ;
        RECT 3380.500 2238.985 3380.670 2239.155 ;
        RECT 3385.940 2238.985 3386.110 2239.155 ;
        RECT 3380.500 2238.525 3380.670 2238.695 ;
        RECT 3385.940 2238.525 3386.110 2238.695 ;
        RECT 3380.500 2238.065 3380.670 2238.235 ;
        RECT 3385.940 2238.065 3386.110 2238.235 ;
        RECT 3380.500 2237.605 3380.670 2237.775 ;
        RECT 3385.940 2237.605 3386.110 2237.775 ;
        RECT 3380.500 2237.145 3380.670 2237.315 ;
        RECT 3385.940 2237.145 3386.110 2237.315 ;
        RECT 3380.500 2236.685 3380.670 2236.855 ;
        RECT 3385.940 2236.685 3386.110 2236.855 ;
        RECT 3380.500 2236.225 3380.670 2236.395 ;
        RECT 3385.940 2236.225 3386.110 2236.395 ;
        RECT 3380.500 2235.765 3380.670 2235.935 ;
        RECT 3385.940 2235.765 3386.110 2235.935 ;
        RECT 3380.500 2235.305 3380.670 2235.475 ;
        RECT 3385.940 2235.305 3386.110 2235.475 ;
        RECT 3380.500 2234.845 3380.670 2235.015 ;
        RECT 3385.940 2234.845 3386.110 2235.015 ;
        RECT 3380.500 2234.385 3380.670 2234.555 ;
        RECT 3385.940 2234.385 3386.110 2234.555 ;
        RECT 3380.500 2233.925 3380.670 2234.095 ;
        RECT 3385.940 2233.925 3386.110 2234.095 ;
        RECT 3380.500 2233.465 3380.670 2233.635 ;
        RECT 3385.940 2233.465 3386.110 2233.635 ;
        RECT 3380.500 2233.005 3380.670 2233.175 ;
        RECT 3385.940 2233.005 3386.110 2233.175 ;
        RECT 3380.500 2232.545 3380.670 2232.715 ;
        RECT 3385.940 2232.545 3386.110 2232.715 ;
        RECT 3380.500 2232.085 3380.670 2232.255 ;
        RECT 3385.940 2232.085 3386.110 2232.255 ;
        RECT 3380.500 2231.625 3380.670 2231.795 ;
        RECT 3385.940 2231.625 3386.110 2231.795 ;
        RECT 3380.500 2231.165 3380.670 2231.335 ;
        RECT 3385.940 2231.165 3386.110 2231.335 ;
        RECT 3380.500 2230.705 3380.670 2230.875 ;
        RECT 3385.940 2230.705 3386.110 2230.875 ;
        RECT 3380.500 2230.245 3380.670 2230.415 ;
        RECT 3385.940 2230.245 3386.110 2230.415 ;
        RECT 3380.500 2229.785 3380.670 2229.955 ;
        RECT 3385.940 2229.785 3386.110 2229.955 ;
        RECT 3380.500 2229.325 3380.670 2229.495 ;
        RECT 3385.940 2229.325 3386.110 2229.495 ;
        RECT 3380.500 2228.865 3380.670 2229.035 ;
        RECT 3385.940 2228.865 3386.110 2229.035 ;
        RECT 3380.500 2228.405 3380.670 2228.575 ;
        RECT 3385.940 2228.405 3386.110 2228.575 ;
        RECT 3380.500 2227.945 3380.670 2228.115 ;
        RECT 3385.940 2227.945 3386.110 2228.115 ;
        RECT 3380.500 2227.485 3380.670 2227.655 ;
        RECT 3385.940 2227.485 3386.110 2227.655 ;
        RECT 3380.500 2227.025 3380.670 2227.195 ;
        RECT 3385.940 2227.025 3386.110 2227.195 ;
        RECT 3380.500 2226.565 3380.670 2226.735 ;
        RECT 3385.940 2226.565 3386.110 2226.735 ;
        RECT 3380.500 2226.105 3380.670 2226.275 ;
        RECT 3385.940 2226.105 3386.110 2226.275 ;
        RECT 3380.500 2225.645 3380.670 2225.815 ;
        RECT 3385.940 2225.645 3386.110 2225.815 ;
        RECT 3380.500 2225.185 3380.670 2225.355 ;
        RECT 3385.940 2225.185 3386.110 2225.355 ;
        RECT 3380.500 2224.725 3380.670 2224.895 ;
        RECT 3385.940 2224.725 3386.110 2224.895 ;
        RECT 3380.500 2224.265 3380.670 2224.435 ;
        RECT 3385.940 2224.265 3386.110 2224.435 ;
        RECT 3380.500 2223.805 3380.670 2223.975 ;
        RECT 3385.940 2223.805 3386.110 2223.975 ;
        RECT 3380.500 2223.345 3380.670 2223.515 ;
        RECT 3385.940 2223.345 3386.110 2223.515 ;
        RECT 3380.500 2222.885 3380.670 2223.055 ;
        RECT 3385.940 2222.885 3386.110 2223.055 ;
        RECT 3380.500 2222.425 3380.670 2222.595 ;
        RECT 3385.940 2222.425 3386.110 2222.595 ;
        RECT 3380.500 2221.965 3380.670 2222.135 ;
        RECT 3385.940 2221.965 3386.110 2222.135 ;
        RECT 3380.500 2221.505 3380.670 2221.675 ;
        RECT 3385.940 2221.505 3386.110 2221.675 ;
        RECT 3380.500 2221.045 3380.670 2221.215 ;
        RECT 3385.940 2221.045 3386.110 2221.215 ;
        RECT 3380.500 2220.585 3380.670 2220.755 ;
        RECT 3385.940 2220.585 3386.110 2220.755 ;
        RECT 3380.500 2220.125 3380.670 2220.295 ;
        RECT 3385.940 2220.125 3386.110 2220.295 ;
        RECT 3380.500 2219.665 3380.670 2219.835 ;
        RECT 3385.940 2219.665 3386.110 2219.835 ;
        RECT 3380.500 2219.205 3380.670 2219.375 ;
        RECT 3385.940 2219.205 3386.110 2219.375 ;
        RECT 3380.500 2218.745 3380.670 2218.915 ;
        RECT 3385.940 2218.745 3386.110 2218.915 ;
        RECT 3380.500 2218.285 3380.670 2218.455 ;
        RECT 3385.940 2218.285 3386.110 2218.455 ;
        RECT 3380.500 2217.825 3380.670 2217.995 ;
        RECT 3385.940 2217.825 3386.110 2217.995 ;
        RECT 3380.500 2217.365 3380.670 2217.535 ;
        RECT 3385.940 2217.365 3386.110 2217.535 ;
        RECT 3380.500 2216.905 3380.670 2217.075 ;
        RECT 3385.940 2216.905 3386.110 2217.075 ;
        RECT 3380.500 2216.445 3380.670 2216.615 ;
        RECT 3385.940 2216.445 3386.110 2216.615 ;
        RECT 3380.500 2215.985 3380.670 2216.155 ;
        RECT 3385.940 2215.985 3386.110 2216.155 ;
        RECT 3380.500 2215.525 3380.670 2215.695 ;
        RECT 3385.940 2215.525 3386.110 2215.695 ;
        RECT 3380.500 2215.065 3380.670 2215.235 ;
        RECT 3385.940 2215.065 3386.110 2215.235 ;
        RECT 3380.500 2214.605 3380.670 2214.775 ;
        RECT 3385.940 2214.605 3386.110 2214.775 ;
        RECT 3380.500 2214.145 3380.670 2214.315 ;
        RECT 3385.940 2214.145 3386.110 2214.315 ;
        RECT 3380.500 2213.685 3380.670 2213.855 ;
        RECT 3385.940 2213.685 3386.110 2213.855 ;
        RECT 3380.500 2213.225 3380.670 2213.395 ;
        RECT 3385.940 2213.225 3386.110 2213.395 ;
        RECT 3380.500 2212.765 3380.670 2212.935 ;
        RECT 3385.940 2212.765 3386.110 2212.935 ;
        RECT 3380.500 2212.305 3380.670 2212.475 ;
        RECT 3385.940 2212.305 3386.110 2212.475 ;
        RECT 3380.500 2211.845 3380.670 2212.015 ;
        RECT 3385.940 2211.845 3386.110 2212.015 ;
        RECT 3380.500 2211.385 3380.670 2211.555 ;
        RECT 3385.940 2211.385 3386.110 2211.555 ;
        RECT 3380.500 2210.925 3380.670 2211.095 ;
        RECT 3385.940 2210.925 3386.110 2211.095 ;
        RECT 3380.500 2210.465 3380.670 2210.635 ;
        RECT 3385.940 2210.465 3386.110 2210.635 ;
        RECT 3380.500 2210.005 3380.670 2210.175 ;
        RECT 3385.940 2210.005 3386.110 2210.175 ;
        RECT 3380.500 2209.545 3380.670 2209.715 ;
        RECT 3385.940 2209.545 3386.110 2209.715 ;
        RECT 3380.500 2209.085 3380.670 2209.255 ;
        RECT 3385.940 2209.085 3386.110 2209.255 ;
        RECT 3380.500 2208.625 3380.670 2208.795 ;
        RECT 3385.940 2208.625 3386.110 2208.795 ;
        RECT 3380.500 2208.165 3380.670 2208.335 ;
        RECT 3385.940 2208.165 3386.110 2208.335 ;
        RECT 3380.500 2207.705 3380.670 2207.875 ;
        RECT 3385.940 2207.705 3386.110 2207.875 ;
        RECT 3380.500 2207.245 3380.670 2207.415 ;
        RECT 3385.940 2207.245 3386.110 2207.415 ;
        RECT 3380.500 2206.785 3380.670 2206.955 ;
        RECT 3385.940 2206.785 3386.110 2206.955 ;
        RECT 3380.500 2206.325 3380.670 2206.495 ;
        RECT 3385.940 2206.325 3386.110 2206.495 ;
        RECT 3380.500 2205.865 3380.670 2206.035 ;
        RECT 3385.940 2205.865 3386.110 2206.035 ;
        RECT 3380.500 2205.405 3380.670 2205.575 ;
        RECT 3385.940 2205.405 3386.110 2205.575 ;
        RECT 3380.500 2204.945 3380.670 2205.115 ;
        RECT 3385.940 2204.945 3386.110 2205.115 ;
        RECT 3380.500 2204.485 3380.670 2204.655 ;
        RECT 3385.940 2204.485 3386.110 2204.655 ;
        RECT 3380.500 2204.025 3380.670 2204.195 ;
        RECT 3385.940 2204.025 3386.110 2204.195 ;
        RECT 3380.500 2203.565 3380.670 2203.735 ;
        RECT 3385.940 2203.565 3386.110 2203.735 ;
        RECT 3380.500 2203.105 3380.670 2203.275 ;
        RECT 3385.940 2203.105 3386.110 2203.275 ;
        RECT 3380.500 2202.645 3380.670 2202.815 ;
        RECT 3385.940 2202.645 3386.110 2202.815 ;
        RECT 3380.500 2202.185 3380.670 2202.355 ;
        RECT 3385.940 2202.185 3386.110 2202.355 ;
      LAYER li1 ;
        RECT 3380.500 2201.955 3380.670 2202.040 ;
        RECT 3379.955 2201.895 3380.670 2201.955 ;
        RECT 3379.955 2201.725 3380.500 2201.895 ;
      LAYER li1 ;
        RECT 3385.940 2201.725 3386.110 2201.895 ;
      LAYER li1 ;
        RECT 3379.955 2200.370 3380.670 2201.725 ;
      LAYER li1 ;
        RECT 3385.940 2201.265 3386.110 2201.435 ;
        RECT 3385.940 2200.805 3386.110 2200.975 ;
      LAYER li1 ;
        RECT 3379.125 2200.030 3380.670 2200.370 ;
      LAYER li1 ;
        RECT 3385.940 2200.345 3386.110 2200.515 ;
      LAYER li1 ;
        RECT 3379.955 2196.610 3380.670 2200.030 ;
      LAYER li1 ;
        RECT 3385.940 2199.885 3386.110 2200.055 ;
        RECT 3385.940 2199.425 3386.110 2199.595 ;
        RECT 3385.940 2198.965 3386.110 2199.135 ;
        RECT 3385.940 2198.505 3386.110 2198.675 ;
        RECT 3385.940 2198.045 3386.110 2198.215 ;
        RECT 3385.940 2197.585 3386.110 2197.755 ;
        RECT 3385.940 2197.125 3386.110 2197.295 ;
        RECT 3385.940 2196.665 3386.110 2196.835 ;
      LAYER li1 ;
        RECT 3380.500 2196.520 3380.670 2196.610 ;
      LAYER li1 ;
        RECT 3380.500 2196.205 3380.670 2196.375 ;
        RECT 3385.940 2196.205 3386.110 2196.375 ;
      LAYER mcon ;
        RECT 3380.500 2201.265 3380.670 2201.435 ;
        RECT 3380.500 2200.805 3380.670 2200.975 ;
        RECT 3380.500 2200.345 3380.670 2200.515 ;
        RECT 3380.500 2199.885 3380.670 2200.055 ;
        RECT 3380.500 2199.425 3380.670 2199.595 ;
        RECT 3380.500 2198.965 3380.670 2199.135 ;
        RECT 3380.500 2198.505 3380.670 2198.675 ;
        RECT 3380.500 2198.045 3380.670 2198.215 ;
        RECT 3380.500 2197.585 3380.670 2197.755 ;
        RECT 3380.500 2197.125 3380.670 2197.295 ;
        RECT 3380.500 2196.665 3380.670 2196.835 ;
      LAYER met1 ;
        RECT 3380.345 2196.060 3380.825 2268.280 ;
        RECT 3385.785 2196.060 3386.265 2268.280 ;
      LAYER via ;
        RECT 3380.425 2240.475 3380.725 2242.260 ;
        RECT 3385.835 2240.475 3386.135 2242.260 ;
      LAYER met2 ;
        RECT 3380.365 2240.435 3380.795 2242.300 ;
        RECT 3385.790 2240.435 3386.220 2242.300 ;
      LAYER via2 ;
        RECT 3380.425 2240.475 3380.725 2242.260 ;
        RECT 3385.835 2240.475 3386.135 2242.260 ;
      LAYER met3 ;
        RECT 3380.350 2240.440 3387.875 2242.305 ;
    END
    PORT
      LAYER li1 ;
        RECT 3380.500 3638.085 3380.670 3638.255 ;
        RECT 3385.940 3638.085 3386.110 3638.255 ;
        RECT 3380.500 3637.625 3380.670 3637.795 ;
        RECT 3385.940 3637.625 3386.110 3637.795 ;
        RECT 3380.500 3637.165 3380.670 3637.335 ;
        RECT 3385.940 3637.165 3386.110 3637.335 ;
        RECT 3380.500 3636.705 3380.670 3636.875 ;
        RECT 3385.940 3636.705 3386.110 3636.875 ;
        RECT 3380.500 3636.245 3380.670 3636.415 ;
        RECT 3385.940 3636.245 3386.110 3636.415 ;
        RECT 3380.500 3635.785 3380.670 3635.955 ;
        RECT 3385.940 3635.785 3386.110 3635.955 ;
        RECT 3380.500 3635.325 3380.670 3635.495 ;
        RECT 3385.940 3635.325 3386.110 3635.495 ;
        RECT 3380.500 3634.865 3380.670 3635.035 ;
        RECT 3385.940 3634.865 3386.110 3635.035 ;
        RECT 3380.500 3634.405 3380.670 3634.575 ;
        RECT 3385.940 3634.405 3386.110 3634.575 ;
        RECT 3380.500 3633.945 3380.670 3634.115 ;
        RECT 3385.940 3633.945 3386.110 3634.115 ;
        RECT 3380.500 3633.485 3380.670 3633.655 ;
        RECT 3385.940 3633.485 3386.110 3633.655 ;
        RECT 3380.500 3633.025 3380.670 3633.195 ;
        RECT 3385.940 3633.025 3386.110 3633.195 ;
        RECT 3380.500 3632.565 3380.670 3632.735 ;
        RECT 3385.940 3632.565 3386.110 3632.735 ;
        RECT 3380.500 3632.105 3380.670 3632.275 ;
        RECT 3385.940 3632.105 3386.110 3632.275 ;
        RECT 3380.500 3631.645 3380.670 3631.815 ;
        RECT 3385.940 3631.645 3386.110 3631.815 ;
        RECT 3380.500 3631.185 3380.670 3631.355 ;
        RECT 3385.940 3631.185 3386.110 3631.355 ;
        RECT 3380.500 3630.725 3380.670 3630.895 ;
        RECT 3385.940 3630.725 3386.110 3630.895 ;
        RECT 3380.500 3630.265 3380.670 3630.435 ;
        RECT 3385.940 3630.265 3386.110 3630.435 ;
        RECT 3380.500 3629.805 3380.670 3629.975 ;
        RECT 3385.940 3629.805 3386.110 3629.975 ;
        RECT 3380.500 3629.345 3380.670 3629.515 ;
        RECT 3385.940 3629.345 3386.110 3629.515 ;
        RECT 3380.500 3628.885 3380.670 3629.055 ;
        RECT 3385.940 3628.885 3386.110 3629.055 ;
        RECT 3380.500 3628.425 3380.670 3628.595 ;
        RECT 3385.940 3628.425 3386.110 3628.595 ;
        RECT 3380.500 3627.965 3380.670 3628.135 ;
        RECT 3385.940 3627.965 3386.110 3628.135 ;
        RECT 3380.500 3627.505 3380.670 3627.675 ;
        RECT 3385.940 3627.505 3386.110 3627.675 ;
        RECT 3380.500 3627.045 3380.670 3627.215 ;
        RECT 3385.940 3627.045 3386.110 3627.215 ;
        RECT 3380.500 3626.585 3380.670 3626.755 ;
        RECT 3385.940 3626.585 3386.110 3626.755 ;
        RECT 3380.500 3626.125 3380.670 3626.295 ;
        RECT 3385.940 3626.125 3386.110 3626.295 ;
        RECT 3380.500 3625.665 3380.670 3625.835 ;
        RECT 3385.940 3625.665 3386.110 3625.835 ;
        RECT 3380.500 3625.205 3380.670 3625.375 ;
        RECT 3385.940 3625.205 3386.110 3625.375 ;
        RECT 3380.500 3624.745 3380.670 3624.915 ;
        RECT 3385.940 3624.745 3386.110 3624.915 ;
        RECT 3380.500 3624.285 3380.670 3624.455 ;
        RECT 3385.940 3624.285 3386.110 3624.455 ;
        RECT 3380.500 3623.825 3380.670 3623.995 ;
        RECT 3385.940 3623.825 3386.110 3623.995 ;
        RECT 3380.500 3623.365 3380.670 3623.535 ;
        RECT 3385.940 3623.365 3386.110 3623.535 ;
        RECT 3380.500 3622.905 3380.670 3623.075 ;
        RECT 3385.940 3622.905 3386.110 3623.075 ;
        RECT 3380.500 3622.445 3380.670 3622.615 ;
        RECT 3385.940 3622.445 3386.110 3622.615 ;
        RECT 3380.500 3621.985 3380.670 3622.155 ;
        RECT 3385.940 3621.985 3386.110 3622.155 ;
        RECT 3380.500 3621.525 3380.670 3621.695 ;
        RECT 3385.940 3621.525 3386.110 3621.695 ;
        RECT 3380.500 3621.065 3380.670 3621.235 ;
        RECT 3385.940 3621.065 3386.110 3621.235 ;
        RECT 3380.500 3620.605 3380.670 3620.775 ;
        RECT 3385.940 3620.605 3386.110 3620.775 ;
        RECT 3380.500 3620.145 3380.670 3620.315 ;
        RECT 3385.940 3620.145 3386.110 3620.315 ;
        RECT 3380.500 3619.685 3380.670 3619.855 ;
        RECT 3385.940 3619.685 3386.110 3619.855 ;
        RECT 3380.500 3619.225 3380.670 3619.395 ;
        RECT 3385.940 3619.225 3386.110 3619.395 ;
        RECT 3380.500 3618.765 3380.670 3618.935 ;
        RECT 3385.940 3618.765 3386.110 3618.935 ;
        RECT 3380.500 3618.305 3380.670 3618.475 ;
        RECT 3385.940 3618.305 3386.110 3618.475 ;
        RECT 3380.500 3617.845 3380.670 3618.015 ;
        RECT 3385.940 3617.845 3386.110 3618.015 ;
        RECT 3380.500 3617.385 3380.670 3617.555 ;
        RECT 3385.940 3617.385 3386.110 3617.555 ;
        RECT 3380.500 3616.925 3380.670 3617.095 ;
        RECT 3385.940 3616.925 3386.110 3617.095 ;
        RECT 3380.500 3616.465 3380.670 3616.635 ;
        RECT 3385.940 3616.465 3386.110 3616.635 ;
        RECT 3380.500 3616.005 3380.670 3616.175 ;
        RECT 3385.940 3616.005 3386.110 3616.175 ;
        RECT 3380.500 3615.545 3380.670 3615.715 ;
        RECT 3385.940 3615.545 3386.110 3615.715 ;
        RECT 3380.500 3615.085 3380.670 3615.255 ;
        RECT 3385.940 3615.085 3386.110 3615.255 ;
        RECT 3380.500 3614.625 3380.670 3614.795 ;
        RECT 3385.940 3614.625 3386.110 3614.795 ;
        RECT 3380.500 3614.165 3380.670 3614.335 ;
        RECT 3385.940 3614.165 3386.110 3614.335 ;
        RECT 3380.500 3613.705 3380.670 3613.875 ;
        RECT 3385.940 3613.705 3386.110 3613.875 ;
        RECT 3380.500 3613.245 3380.670 3613.415 ;
        RECT 3385.940 3613.245 3386.110 3613.415 ;
        RECT 3380.500 3612.785 3380.670 3612.955 ;
        RECT 3385.940 3612.785 3386.110 3612.955 ;
        RECT 3380.500 3612.325 3380.670 3612.495 ;
        RECT 3385.940 3612.325 3386.110 3612.495 ;
        RECT 3380.500 3611.865 3380.670 3612.035 ;
        RECT 3385.940 3611.865 3386.110 3612.035 ;
        RECT 3380.500 3611.405 3380.670 3611.575 ;
        RECT 3385.940 3611.405 3386.110 3611.575 ;
        RECT 3380.500 3610.945 3380.670 3611.115 ;
        RECT 3385.940 3610.945 3386.110 3611.115 ;
        RECT 3380.500 3610.485 3380.670 3610.655 ;
        RECT 3385.940 3610.485 3386.110 3610.655 ;
        RECT 3380.500 3610.025 3380.670 3610.195 ;
        RECT 3385.940 3610.025 3386.110 3610.195 ;
        RECT 3380.500 3609.565 3380.670 3609.735 ;
        RECT 3385.940 3609.565 3386.110 3609.735 ;
        RECT 3380.500 3609.105 3380.670 3609.275 ;
        RECT 3385.940 3609.105 3386.110 3609.275 ;
        RECT 3380.500 3608.645 3380.670 3608.815 ;
        RECT 3385.940 3608.645 3386.110 3608.815 ;
        RECT 3380.500 3608.185 3380.670 3608.355 ;
        RECT 3385.940 3608.185 3386.110 3608.355 ;
        RECT 3380.500 3607.725 3380.670 3607.895 ;
        RECT 3385.940 3607.725 3386.110 3607.895 ;
        RECT 3380.500 3607.265 3380.670 3607.435 ;
        RECT 3385.940 3607.265 3386.110 3607.435 ;
        RECT 3380.500 3606.805 3380.670 3606.975 ;
        RECT 3385.940 3606.805 3386.110 3606.975 ;
        RECT 3380.500 3606.345 3380.670 3606.515 ;
        RECT 3385.940 3606.345 3386.110 3606.515 ;
        RECT 3380.500 3605.885 3380.670 3606.055 ;
        RECT 3385.940 3605.885 3386.110 3606.055 ;
        RECT 3380.500 3605.425 3380.670 3605.595 ;
        RECT 3385.940 3605.425 3386.110 3605.595 ;
        RECT 3380.500 3604.965 3380.670 3605.135 ;
        RECT 3385.940 3604.965 3386.110 3605.135 ;
        RECT 3380.500 3604.505 3380.670 3604.675 ;
        RECT 3385.940 3604.505 3386.110 3604.675 ;
        RECT 3380.500 3604.045 3380.670 3604.215 ;
        RECT 3385.940 3604.045 3386.110 3604.215 ;
        RECT 3380.500 3603.585 3380.670 3603.755 ;
        RECT 3385.940 3603.585 3386.110 3603.755 ;
        RECT 3380.500 3603.125 3380.670 3603.295 ;
        RECT 3385.940 3603.125 3386.110 3603.295 ;
        RECT 3380.500 3602.665 3380.670 3602.835 ;
        RECT 3385.940 3602.665 3386.110 3602.835 ;
        RECT 3380.500 3602.205 3380.670 3602.375 ;
        RECT 3385.940 3602.205 3386.110 3602.375 ;
      LAYER met1 ;
        RECT 3380.345 3602.060 3380.825 3638.400 ;
        RECT 3385.785 3602.060 3386.265 3638.400 ;
      LAYER via ;
        RECT 3380.465 3622.480 3380.765 3624.265 ;
        RECT 3385.875 3622.480 3386.175 3624.265 ;
      LAYER met2 ;
        RECT 3380.405 3622.440 3380.835 3624.305 ;
        RECT 3385.830 3622.440 3386.260 3624.305 ;
      LAYER via2 ;
        RECT 3380.465 3622.480 3380.765 3624.265 ;
        RECT 3385.875 3622.480 3386.175 3624.265 ;
      LAYER met3 ;
        RECT 3380.390 3622.445 3387.915 3624.310 ;
    END
    PORT
      LAYER li1 ;
        RECT 677.110 217.755 677.450 218.585 ;
        RECT 683.090 217.755 683.430 218.585 ;
        RECT 689.070 217.755 689.410 218.585 ;
        RECT 695.050 217.755 695.390 218.585 ;
        RECT 701.030 217.755 701.370 218.585 ;
        RECT 707.010 217.755 707.350 218.585 ;
        RECT 712.990 217.755 713.330 218.585 ;
        RECT 718.970 217.755 719.310 218.585 ;
        RECT 724.950 217.755 725.290 218.585 ;
        RECT 730.930 217.755 731.270 218.585 ;
        RECT 736.910 217.755 737.250 218.585 ;
        RECT 742.890 217.755 743.230 218.585 ;
        RECT 748.870 217.755 749.210 218.585 ;
        RECT 754.850 217.755 755.190 218.585 ;
        RECT 760.830 217.755 761.170 218.585 ;
        RECT 766.810 217.755 767.150 218.585 ;
        RECT 772.790 217.755 773.130 218.585 ;
        RECT 778.770 217.755 779.110 218.585 ;
        RECT 784.750 217.755 785.090 218.585 ;
        RECT 790.730 217.755 791.070 218.585 ;
        RECT 675.525 217.210 680.870 217.755 ;
        RECT 681.505 217.210 686.850 217.755 ;
        RECT 687.485 217.210 692.830 217.755 ;
        RECT 693.465 217.210 698.810 217.755 ;
        RECT 699.445 217.210 704.790 217.755 ;
        RECT 705.425 217.210 710.770 217.755 ;
        RECT 711.405 217.210 716.750 217.755 ;
        RECT 717.385 217.210 722.730 217.755 ;
        RECT 723.365 217.210 728.710 217.755 ;
        RECT 729.345 217.210 734.690 217.755 ;
        RECT 735.325 217.210 740.670 217.755 ;
        RECT 741.305 217.210 746.650 217.755 ;
        RECT 747.285 217.210 752.630 217.755 ;
        RECT 753.265 217.210 758.610 217.755 ;
        RECT 759.245 217.210 764.590 217.755 ;
        RECT 765.225 217.210 770.570 217.755 ;
        RECT 771.205 217.210 776.550 217.755 ;
        RECT 777.185 217.210 782.530 217.755 ;
        RECT 783.165 217.210 788.510 217.755 ;
        RECT 789.145 217.210 794.490 217.755 ;
      LAYER li1 ;
        RECT 669.145 217.040 669.315 217.210 ;
        RECT 669.605 217.040 669.775 217.210 ;
        RECT 670.065 217.040 670.235 217.210 ;
        RECT 670.525 217.040 670.695 217.210 ;
        RECT 670.985 217.040 671.155 217.210 ;
        RECT 671.445 217.040 671.615 217.210 ;
        RECT 671.905 217.040 672.075 217.210 ;
        RECT 672.365 217.040 672.535 217.210 ;
        RECT 672.825 217.040 672.995 217.210 ;
        RECT 673.285 217.040 673.455 217.210 ;
        RECT 673.745 217.040 673.915 217.210 ;
        RECT 674.205 217.040 674.375 217.210 ;
        RECT 674.665 217.040 674.835 217.210 ;
        RECT 675.125 217.040 675.295 217.210 ;
      LAYER li1 ;
        RECT 675.440 217.040 675.585 217.210 ;
        RECT 675.755 217.040 680.960 217.210 ;
      LAYER li1 ;
        RECT 681.105 217.040 681.275 217.210 ;
      LAYER li1 ;
        RECT 681.420 217.040 681.565 217.210 ;
        RECT 681.735 217.040 686.940 217.210 ;
      LAYER li1 ;
        RECT 687.085 217.040 687.255 217.210 ;
      LAYER li1 ;
        RECT 687.400 217.040 687.545 217.210 ;
        RECT 687.715 217.040 692.920 217.210 ;
      LAYER li1 ;
        RECT 693.065 217.040 693.235 217.210 ;
      LAYER li1 ;
        RECT 693.380 217.040 693.525 217.210 ;
        RECT 693.695 217.040 698.900 217.210 ;
      LAYER li1 ;
        RECT 699.045 217.040 699.215 217.210 ;
      LAYER li1 ;
        RECT 699.360 217.040 699.505 217.210 ;
        RECT 699.675 217.040 704.880 217.210 ;
      LAYER li1 ;
        RECT 705.025 217.040 705.195 217.210 ;
      LAYER li1 ;
        RECT 705.340 217.040 705.485 217.210 ;
        RECT 705.655 217.040 710.860 217.210 ;
      LAYER li1 ;
        RECT 711.005 217.040 711.175 217.210 ;
      LAYER li1 ;
        RECT 711.320 217.040 711.465 217.210 ;
        RECT 711.635 217.040 716.840 217.210 ;
      LAYER li1 ;
        RECT 716.985 217.040 717.155 217.210 ;
      LAYER li1 ;
        RECT 717.300 217.040 717.445 217.210 ;
        RECT 717.615 217.040 722.820 217.210 ;
      LAYER li1 ;
        RECT 722.965 217.040 723.135 217.210 ;
      LAYER li1 ;
        RECT 723.280 217.040 723.425 217.210 ;
        RECT 723.595 217.040 728.800 217.210 ;
      LAYER li1 ;
        RECT 728.945 217.040 729.115 217.210 ;
      LAYER li1 ;
        RECT 729.260 217.040 729.405 217.210 ;
        RECT 729.575 217.040 734.780 217.210 ;
      LAYER li1 ;
        RECT 734.925 217.040 735.095 217.210 ;
      LAYER li1 ;
        RECT 735.240 217.040 735.385 217.210 ;
        RECT 735.555 217.040 740.760 217.210 ;
      LAYER li1 ;
        RECT 740.905 217.040 741.075 217.210 ;
      LAYER li1 ;
        RECT 741.220 217.040 741.365 217.210 ;
        RECT 741.535 217.040 746.740 217.210 ;
      LAYER li1 ;
        RECT 746.885 217.040 747.055 217.210 ;
      LAYER li1 ;
        RECT 747.200 217.040 747.345 217.210 ;
        RECT 747.515 217.040 752.720 217.210 ;
      LAYER li1 ;
        RECT 752.865 217.040 753.035 217.210 ;
      LAYER li1 ;
        RECT 753.180 217.040 753.325 217.210 ;
        RECT 753.495 217.040 758.700 217.210 ;
      LAYER li1 ;
        RECT 758.845 217.040 759.015 217.210 ;
      LAYER li1 ;
        RECT 759.160 217.040 759.305 217.210 ;
        RECT 759.475 217.040 764.680 217.210 ;
      LAYER li1 ;
        RECT 764.825 217.040 764.995 217.210 ;
      LAYER li1 ;
        RECT 765.140 217.040 765.285 217.210 ;
        RECT 765.455 217.040 770.660 217.210 ;
      LAYER li1 ;
        RECT 770.805 217.040 770.975 217.210 ;
      LAYER li1 ;
        RECT 771.120 217.040 771.265 217.210 ;
        RECT 771.435 217.040 776.640 217.210 ;
      LAYER li1 ;
        RECT 776.785 217.040 776.955 217.210 ;
      LAYER li1 ;
        RECT 777.100 217.040 777.245 217.210 ;
        RECT 777.415 217.040 782.620 217.210 ;
      LAYER li1 ;
        RECT 782.765 217.040 782.935 217.210 ;
      LAYER li1 ;
        RECT 783.080 217.040 783.225 217.210 ;
        RECT 783.395 217.040 788.600 217.210 ;
      LAYER li1 ;
        RECT 788.745 217.040 788.915 217.210 ;
      LAYER li1 ;
        RECT 789.060 217.040 789.205 217.210 ;
        RECT 789.375 217.040 794.580 217.210 ;
      LAYER li1 ;
        RECT 794.725 217.040 794.895 217.210 ;
      LAYER li1 ;
        RECT 671.130 212.315 671.470 213.145 ;
        RECT 669.545 211.770 674.890 212.315 ;
      LAYER li1 ;
        RECT 669.145 211.600 669.315 211.770 ;
      LAYER li1 ;
        RECT 669.460 211.600 674.980 211.770 ;
      LAYER li1 ;
        RECT 675.125 211.600 675.295 211.770 ;
        RECT 675.585 211.600 675.755 211.770 ;
        RECT 676.045 211.600 676.215 211.770 ;
        RECT 676.505 211.600 676.675 211.770 ;
        RECT 676.965 211.600 677.135 211.770 ;
        RECT 677.425 211.600 677.595 211.770 ;
        RECT 677.885 211.600 678.055 211.770 ;
        RECT 678.345 211.600 678.515 211.770 ;
        RECT 678.805 211.600 678.975 211.770 ;
        RECT 679.265 211.600 679.435 211.770 ;
        RECT 679.725 211.600 679.895 211.770 ;
        RECT 680.185 211.600 680.355 211.770 ;
        RECT 680.645 211.600 680.815 211.770 ;
        RECT 681.105 211.600 681.275 211.770 ;
        RECT 681.565 211.600 681.735 211.770 ;
        RECT 682.025 211.600 682.195 211.770 ;
        RECT 682.485 211.600 682.655 211.770 ;
        RECT 682.945 211.600 683.115 211.770 ;
        RECT 683.405 211.600 683.575 211.770 ;
        RECT 683.865 211.600 684.035 211.770 ;
        RECT 684.325 211.600 684.495 211.770 ;
        RECT 684.785 211.600 684.955 211.770 ;
        RECT 685.245 211.600 685.415 211.770 ;
        RECT 685.705 211.600 685.875 211.770 ;
        RECT 686.165 211.600 686.335 211.770 ;
        RECT 686.625 211.600 686.795 211.770 ;
        RECT 687.085 211.600 687.255 211.770 ;
        RECT 687.545 211.600 687.715 211.770 ;
        RECT 688.005 211.600 688.175 211.770 ;
        RECT 688.465 211.600 688.635 211.770 ;
        RECT 688.925 211.600 689.095 211.770 ;
        RECT 689.385 211.600 689.555 211.770 ;
        RECT 689.845 211.600 690.015 211.770 ;
        RECT 690.305 211.600 690.475 211.770 ;
        RECT 690.765 211.600 690.935 211.770 ;
        RECT 691.225 211.600 691.395 211.770 ;
        RECT 691.685 211.600 691.855 211.770 ;
        RECT 692.145 211.600 692.315 211.770 ;
        RECT 692.605 211.600 692.775 211.770 ;
        RECT 693.065 211.600 693.235 211.770 ;
        RECT 693.525 211.600 693.695 211.770 ;
        RECT 693.985 211.600 694.155 211.770 ;
        RECT 694.445 211.600 694.615 211.770 ;
        RECT 694.905 211.600 695.075 211.770 ;
        RECT 695.365 211.600 695.535 211.770 ;
        RECT 695.825 211.600 695.995 211.770 ;
        RECT 696.285 211.600 696.455 211.770 ;
        RECT 696.745 211.600 696.915 211.770 ;
        RECT 697.205 211.600 697.375 211.770 ;
        RECT 697.665 211.600 697.835 211.770 ;
        RECT 698.125 211.600 698.295 211.770 ;
        RECT 698.585 211.600 698.755 211.770 ;
        RECT 699.045 211.600 699.215 211.770 ;
        RECT 699.505 211.600 699.675 211.770 ;
        RECT 699.965 211.600 700.135 211.770 ;
        RECT 700.425 211.600 700.595 211.770 ;
        RECT 700.885 211.600 701.055 211.770 ;
        RECT 701.345 211.600 701.515 211.770 ;
        RECT 701.805 211.600 701.975 211.770 ;
        RECT 702.265 211.600 702.435 211.770 ;
        RECT 702.725 211.600 702.895 211.770 ;
        RECT 703.185 211.600 703.355 211.770 ;
        RECT 703.645 211.600 703.815 211.770 ;
        RECT 704.105 211.600 704.275 211.770 ;
        RECT 704.565 211.600 704.735 211.770 ;
        RECT 705.025 211.600 705.195 211.770 ;
        RECT 705.485 211.600 705.655 211.770 ;
        RECT 705.945 211.600 706.115 211.770 ;
        RECT 706.405 211.600 706.575 211.770 ;
        RECT 706.865 211.600 707.035 211.770 ;
        RECT 707.325 211.600 707.495 211.770 ;
        RECT 707.785 211.600 707.955 211.770 ;
        RECT 708.245 211.600 708.415 211.770 ;
        RECT 708.705 211.600 708.875 211.770 ;
        RECT 709.165 211.600 709.335 211.770 ;
        RECT 709.625 211.600 709.795 211.770 ;
        RECT 710.085 211.600 710.255 211.770 ;
        RECT 710.545 211.600 710.715 211.770 ;
        RECT 711.005 211.600 711.175 211.770 ;
        RECT 711.465 211.600 711.635 211.770 ;
        RECT 711.925 211.600 712.095 211.770 ;
        RECT 712.385 211.600 712.555 211.770 ;
        RECT 712.845 211.600 713.015 211.770 ;
        RECT 713.305 211.600 713.475 211.770 ;
        RECT 713.765 211.600 713.935 211.770 ;
        RECT 714.225 211.600 714.395 211.770 ;
        RECT 714.685 211.600 714.855 211.770 ;
        RECT 715.145 211.600 715.315 211.770 ;
        RECT 715.605 211.600 715.775 211.770 ;
        RECT 716.065 211.600 716.235 211.770 ;
        RECT 716.525 211.600 716.695 211.770 ;
        RECT 716.985 211.600 717.155 211.770 ;
        RECT 717.445 211.600 717.615 211.770 ;
        RECT 717.905 211.600 718.075 211.770 ;
        RECT 718.365 211.600 718.535 211.770 ;
        RECT 718.825 211.600 718.995 211.770 ;
        RECT 719.285 211.600 719.455 211.770 ;
        RECT 719.745 211.600 719.915 211.770 ;
        RECT 720.205 211.600 720.375 211.770 ;
        RECT 720.665 211.600 720.835 211.770 ;
        RECT 721.125 211.600 721.295 211.770 ;
        RECT 721.585 211.600 721.755 211.770 ;
        RECT 722.045 211.600 722.215 211.770 ;
        RECT 722.505 211.600 722.675 211.770 ;
        RECT 722.965 211.600 723.135 211.770 ;
        RECT 723.425 211.600 723.595 211.770 ;
        RECT 723.885 211.600 724.055 211.770 ;
        RECT 724.345 211.600 724.515 211.770 ;
        RECT 724.805 211.600 724.975 211.770 ;
        RECT 725.265 211.600 725.435 211.770 ;
        RECT 725.725 211.600 725.895 211.770 ;
        RECT 726.185 211.600 726.355 211.770 ;
        RECT 726.645 211.600 726.815 211.770 ;
        RECT 727.105 211.600 727.275 211.770 ;
        RECT 727.565 211.600 727.735 211.770 ;
        RECT 728.025 211.600 728.195 211.770 ;
        RECT 728.485 211.600 728.655 211.770 ;
        RECT 728.945 211.600 729.115 211.770 ;
        RECT 729.405 211.600 729.575 211.770 ;
        RECT 729.865 211.600 730.035 211.770 ;
        RECT 730.325 211.600 730.495 211.770 ;
        RECT 730.785 211.600 730.955 211.770 ;
        RECT 731.245 211.600 731.415 211.770 ;
        RECT 731.705 211.600 731.875 211.770 ;
        RECT 732.165 211.600 732.335 211.770 ;
        RECT 732.625 211.600 732.795 211.770 ;
        RECT 733.085 211.600 733.255 211.770 ;
        RECT 733.545 211.600 733.715 211.770 ;
        RECT 734.005 211.600 734.175 211.770 ;
        RECT 734.465 211.600 734.635 211.770 ;
        RECT 734.925 211.600 735.095 211.770 ;
        RECT 735.385 211.600 735.555 211.770 ;
        RECT 735.845 211.600 736.015 211.770 ;
        RECT 736.305 211.600 736.475 211.770 ;
        RECT 736.765 211.600 736.935 211.770 ;
        RECT 737.225 211.600 737.395 211.770 ;
        RECT 737.685 211.600 737.855 211.770 ;
        RECT 738.145 211.600 738.315 211.770 ;
        RECT 738.605 211.600 738.775 211.770 ;
        RECT 739.065 211.600 739.235 211.770 ;
        RECT 739.525 211.600 739.695 211.770 ;
        RECT 739.985 211.600 740.155 211.770 ;
        RECT 740.445 211.600 740.615 211.770 ;
        RECT 740.905 211.600 741.075 211.770 ;
        RECT 741.365 211.600 741.535 211.770 ;
        RECT 741.825 211.600 741.995 211.770 ;
        RECT 742.285 211.600 742.455 211.770 ;
        RECT 742.745 211.600 742.915 211.770 ;
        RECT 743.205 211.600 743.375 211.770 ;
        RECT 743.665 211.600 743.835 211.770 ;
        RECT 744.125 211.600 744.295 211.770 ;
        RECT 744.585 211.600 744.755 211.770 ;
        RECT 745.045 211.600 745.215 211.770 ;
        RECT 745.505 211.600 745.675 211.770 ;
        RECT 745.965 211.600 746.135 211.770 ;
        RECT 746.425 211.600 746.595 211.770 ;
        RECT 746.885 211.600 747.055 211.770 ;
        RECT 747.345 211.600 747.515 211.770 ;
        RECT 747.805 211.600 747.975 211.770 ;
        RECT 748.265 211.600 748.435 211.770 ;
        RECT 748.725 211.600 748.895 211.770 ;
        RECT 749.185 211.600 749.355 211.770 ;
        RECT 749.645 211.600 749.815 211.770 ;
        RECT 750.105 211.600 750.275 211.770 ;
        RECT 750.565 211.600 750.735 211.770 ;
        RECT 751.025 211.600 751.195 211.770 ;
        RECT 751.485 211.600 751.655 211.770 ;
        RECT 751.945 211.600 752.115 211.770 ;
        RECT 752.405 211.600 752.575 211.770 ;
        RECT 752.865 211.600 753.035 211.770 ;
        RECT 753.325 211.600 753.495 211.770 ;
        RECT 753.785 211.600 753.955 211.770 ;
        RECT 754.245 211.600 754.415 211.770 ;
        RECT 754.705 211.600 754.875 211.770 ;
        RECT 755.165 211.600 755.335 211.770 ;
        RECT 755.625 211.600 755.795 211.770 ;
        RECT 756.085 211.600 756.255 211.770 ;
        RECT 756.545 211.600 756.715 211.770 ;
        RECT 757.005 211.600 757.175 211.770 ;
        RECT 757.465 211.600 757.635 211.770 ;
        RECT 757.925 211.600 758.095 211.770 ;
        RECT 758.385 211.600 758.555 211.770 ;
        RECT 758.845 211.600 759.015 211.770 ;
        RECT 759.305 211.600 759.475 211.770 ;
        RECT 759.765 211.600 759.935 211.770 ;
        RECT 760.225 211.600 760.395 211.770 ;
        RECT 760.685 211.600 760.855 211.770 ;
        RECT 761.145 211.600 761.315 211.770 ;
        RECT 761.605 211.600 761.775 211.770 ;
        RECT 762.065 211.600 762.235 211.770 ;
        RECT 762.525 211.600 762.695 211.770 ;
        RECT 762.985 211.600 763.155 211.770 ;
        RECT 763.445 211.600 763.615 211.770 ;
        RECT 763.905 211.600 764.075 211.770 ;
        RECT 764.365 211.600 764.535 211.770 ;
        RECT 764.825 211.600 764.995 211.770 ;
        RECT 765.285 211.600 765.455 211.770 ;
        RECT 765.745 211.600 765.915 211.770 ;
        RECT 766.205 211.600 766.375 211.770 ;
        RECT 766.665 211.600 766.835 211.770 ;
        RECT 767.125 211.600 767.295 211.770 ;
        RECT 767.585 211.600 767.755 211.770 ;
        RECT 768.045 211.600 768.215 211.770 ;
        RECT 768.505 211.600 768.675 211.770 ;
        RECT 768.965 211.600 769.135 211.770 ;
        RECT 769.425 211.600 769.595 211.770 ;
        RECT 769.885 211.600 770.055 211.770 ;
        RECT 770.345 211.600 770.515 211.770 ;
        RECT 770.805 211.600 770.975 211.770 ;
        RECT 771.265 211.600 771.435 211.770 ;
        RECT 771.725 211.600 771.895 211.770 ;
        RECT 772.185 211.600 772.355 211.770 ;
        RECT 772.645 211.600 772.815 211.770 ;
        RECT 773.105 211.600 773.275 211.770 ;
        RECT 773.565 211.600 773.735 211.770 ;
        RECT 774.025 211.600 774.195 211.770 ;
        RECT 774.485 211.600 774.655 211.770 ;
        RECT 774.945 211.600 775.115 211.770 ;
        RECT 775.405 211.600 775.575 211.770 ;
        RECT 775.865 211.600 776.035 211.770 ;
        RECT 776.325 211.600 776.495 211.770 ;
        RECT 776.785 211.600 776.955 211.770 ;
        RECT 777.245 211.600 777.415 211.770 ;
        RECT 777.705 211.600 777.875 211.770 ;
        RECT 778.165 211.600 778.335 211.770 ;
        RECT 778.625 211.600 778.795 211.770 ;
        RECT 779.085 211.600 779.255 211.770 ;
        RECT 779.545 211.600 779.715 211.770 ;
        RECT 780.005 211.600 780.175 211.770 ;
        RECT 780.465 211.600 780.635 211.770 ;
        RECT 780.925 211.600 781.095 211.770 ;
        RECT 781.385 211.600 781.555 211.770 ;
        RECT 781.845 211.600 782.015 211.770 ;
        RECT 782.305 211.600 782.475 211.770 ;
        RECT 782.765 211.600 782.935 211.770 ;
        RECT 783.225 211.600 783.395 211.770 ;
        RECT 783.685 211.600 783.855 211.770 ;
        RECT 784.145 211.600 784.315 211.770 ;
        RECT 784.605 211.600 784.775 211.770 ;
        RECT 785.065 211.600 785.235 211.770 ;
        RECT 785.525 211.600 785.695 211.770 ;
        RECT 785.985 211.600 786.155 211.770 ;
        RECT 786.445 211.600 786.615 211.770 ;
        RECT 786.905 211.600 787.075 211.770 ;
        RECT 787.365 211.600 787.535 211.770 ;
        RECT 787.825 211.600 787.995 211.770 ;
        RECT 788.285 211.600 788.455 211.770 ;
        RECT 788.745 211.600 788.915 211.770 ;
        RECT 789.205 211.600 789.375 211.770 ;
        RECT 789.665 211.600 789.835 211.770 ;
        RECT 790.125 211.600 790.295 211.770 ;
        RECT 790.585 211.600 790.755 211.770 ;
        RECT 791.045 211.600 791.215 211.770 ;
        RECT 791.505 211.600 791.675 211.770 ;
        RECT 791.965 211.600 792.135 211.770 ;
        RECT 792.425 211.600 792.595 211.770 ;
        RECT 792.885 211.600 793.055 211.770 ;
        RECT 793.345 211.600 793.515 211.770 ;
        RECT 793.805 211.600 793.975 211.770 ;
        RECT 794.265 211.600 794.435 211.770 ;
        RECT 794.725 211.600 794.895 211.770 ;
      LAYER mcon ;
        RECT 676.045 217.040 676.215 217.210 ;
        RECT 676.505 217.040 676.675 217.210 ;
        RECT 676.965 217.040 677.135 217.210 ;
        RECT 677.425 217.040 677.595 217.210 ;
        RECT 677.885 217.040 678.055 217.210 ;
        RECT 678.345 217.040 678.515 217.210 ;
        RECT 678.805 217.040 678.975 217.210 ;
        RECT 679.265 217.040 679.435 217.210 ;
        RECT 679.725 217.040 679.895 217.210 ;
        RECT 680.185 217.040 680.355 217.210 ;
        RECT 680.645 217.040 680.815 217.210 ;
        RECT 682.025 217.040 682.195 217.210 ;
        RECT 682.485 217.040 682.655 217.210 ;
        RECT 682.945 217.040 683.115 217.210 ;
        RECT 683.405 217.040 683.575 217.210 ;
        RECT 683.865 217.040 684.035 217.210 ;
        RECT 684.325 217.040 684.495 217.210 ;
        RECT 684.785 217.040 684.955 217.210 ;
        RECT 685.245 217.040 685.415 217.210 ;
        RECT 685.705 217.040 685.875 217.210 ;
        RECT 686.165 217.040 686.335 217.210 ;
        RECT 686.625 217.040 686.795 217.210 ;
        RECT 688.005 217.040 688.175 217.210 ;
        RECT 688.465 217.040 688.635 217.210 ;
        RECT 688.925 217.040 689.095 217.210 ;
        RECT 689.385 217.040 689.555 217.210 ;
        RECT 689.845 217.040 690.015 217.210 ;
        RECT 690.305 217.040 690.475 217.210 ;
        RECT 690.765 217.040 690.935 217.210 ;
        RECT 691.225 217.040 691.395 217.210 ;
        RECT 691.685 217.040 691.855 217.210 ;
        RECT 692.145 217.040 692.315 217.210 ;
        RECT 692.605 217.040 692.775 217.210 ;
        RECT 693.985 217.040 694.155 217.210 ;
        RECT 694.445 217.040 694.615 217.210 ;
        RECT 694.905 217.040 695.075 217.210 ;
        RECT 695.365 217.040 695.535 217.210 ;
        RECT 695.825 217.040 695.995 217.210 ;
        RECT 696.285 217.040 696.455 217.210 ;
        RECT 696.745 217.040 696.915 217.210 ;
        RECT 697.205 217.040 697.375 217.210 ;
        RECT 697.665 217.040 697.835 217.210 ;
        RECT 698.125 217.040 698.295 217.210 ;
        RECT 698.585 217.040 698.755 217.210 ;
        RECT 699.965 217.040 700.135 217.210 ;
        RECT 700.425 217.040 700.595 217.210 ;
        RECT 700.885 217.040 701.055 217.210 ;
        RECT 701.345 217.040 701.515 217.210 ;
        RECT 701.805 217.040 701.975 217.210 ;
        RECT 702.265 217.040 702.435 217.210 ;
        RECT 702.725 217.040 702.895 217.210 ;
        RECT 703.185 217.040 703.355 217.210 ;
        RECT 703.645 217.040 703.815 217.210 ;
        RECT 704.105 217.040 704.275 217.210 ;
        RECT 704.565 217.040 704.735 217.210 ;
        RECT 705.945 217.040 706.115 217.210 ;
        RECT 706.405 217.040 706.575 217.210 ;
        RECT 706.865 217.040 707.035 217.210 ;
        RECT 707.325 217.040 707.495 217.210 ;
        RECT 707.785 217.040 707.955 217.210 ;
        RECT 708.245 217.040 708.415 217.210 ;
        RECT 708.705 217.040 708.875 217.210 ;
        RECT 709.165 217.040 709.335 217.210 ;
        RECT 709.625 217.040 709.795 217.210 ;
        RECT 710.085 217.040 710.255 217.210 ;
        RECT 710.545 217.040 710.715 217.210 ;
        RECT 711.925 217.040 712.095 217.210 ;
        RECT 712.385 217.040 712.555 217.210 ;
        RECT 712.845 217.040 713.015 217.210 ;
        RECT 713.305 217.040 713.475 217.210 ;
        RECT 713.765 217.040 713.935 217.210 ;
        RECT 714.225 217.040 714.395 217.210 ;
        RECT 714.685 217.040 714.855 217.210 ;
        RECT 715.145 217.040 715.315 217.210 ;
        RECT 715.605 217.040 715.775 217.210 ;
        RECT 716.065 217.040 716.235 217.210 ;
        RECT 716.525 217.040 716.695 217.210 ;
        RECT 717.905 217.040 718.075 217.210 ;
        RECT 718.365 217.040 718.535 217.210 ;
        RECT 718.825 217.040 718.995 217.210 ;
        RECT 719.285 217.040 719.455 217.210 ;
        RECT 719.745 217.040 719.915 217.210 ;
        RECT 720.205 217.040 720.375 217.210 ;
        RECT 720.665 217.040 720.835 217.210 ;
        RECT 721.125 217.040 721.295 217.210 ;
        RECT 721.585 217.040 721.755 217.210 ;
        RECT 722.045 217.040 722.215 217.210 ;
        RECT 722.505 217.040 722.675 217.210 ;
        RECT 723.885 217.040 724.055 217.210 ;
        RECT 724.345 217.040 724.515 217.210 ;
        RECT 724.805 217.040 724.975 217.210 ;
        RECT 725.265 217.040 725.435 217.210 ;
        RECT 725.725 217.040 725.895 217.210 ;
        RECT 726.185 217.040 726.355 217.210 ;
        RECT 726.645 217.040 726.815 217.210 ;
        RECT 727.105 217.040 727.275 217.210 ;
        RECT 727.565 217.040 727.735 217.210 ;
        RECT 728.025 217.040 728.195 217.210 ;
        RECT 728.485 217.040 728.655 217.210 ;
        RECT 729.865 217.040 730.035 217.210 ;
        RECT 730.325 217.040 730.495 217.210 ;
        RECT 730.785 217.040 730.955 217.210 ;
        RECT 731.245 217.040 731.415 217.210 ;
        RECT 731.705 217.040 731.875 217.210 ;
        RECT 732.165 217.040 732.335 217.210 ;
        RECT 732.625 217.040 732.795 217.210 ;
        RECT 733.085 217.040 733.255 217.210 ;
        RECT 733.545 217.040 733.715 217.210 ;
        RECT 734.005 217.040 734.175 217.210 ;
        RECT 734.465 217.040 734.635 217.210 ;
        RECT 735.845 217.040 736.015 217.210 ;
        RECT 736.305 217.040 736.475 217.210 ;
        RECT 736.765 217.040 736.935 217.210 ;
        RECT 737.225 217.040 737.395 217.210 ;
        RECT 737.685 217.040 737.855 217.210 ;
        RECT 738.145 217.040 738.315 217.210 ;
        RECT 738.605 217.040 738.775 217.210 ;
        RECT 739.065 217.040 739.235 217.210 ;
        RECT 739.525 217.040 739.695 217.210 ;
        RECT 739.985 217.040 740.155 217.210 ;
        RECT 740.445 217.040 740.615 217.210 ;
        RECT 741.825 217.040 741.995 217.210 ;
        RECT 742.285 217.040 742.455 217.210 ;
        RECT 742.745 217.040 742.915 217.210 ;
        RECT 743.205 217.040 743.375 217.210 ;
        RECT 743.665 217.040 743.835 217.210 ;
        RECT 744.125 217.040 744.295 217.210 ;
        RECT 744.585 217.040 744.755 217.210 ;
        RECT 745.045 217.040 745.215 217.210 ;
        RECT 745.505 217.040 745.675 217.210 ;
        RECT 745.965 217.040 746.135 217.210 ;
        RECT 746.425 217.040 746.595 217.210 ;
        RECT 747.805 217.040 747.975 217.210 ;
        RECT 748.265 217.040 748.435 217.210 ;
        RECT 748.725 217.040 748.895 217.210 ;
        RECT 749.185 217.040 749.355 217.210 ;
        RECT 749.645 217.040 749.815 217.210 ;
        RECT 750.105 217.040 750.275 217.210 ;
        RECT 750.565 217.040 750.735 217.210 ;
        RECT 751.025 217.040 751.195 217.210 ;
        RECT 751.485 217.040 751.655 217.210 ;
        RECT 751.945 217.040 752.115 217.210 ;
        RECT 752.405 217.040 752.575 217.210 ;
        RECT 753.785 217.040 753.955 217.210 ;
        RECT 754.245 217.040 754.415 217.210 ;
        RECT 754.705 217.040 754.875 217.210 ;
        RECT 755.165 217.040 755.335 217.210 ;
        RECT 755.625 217.040 755.795 217.210 ;
        RECT 756.085 217.040 756.255 217.210 ;
        RECT 756.545 217.040 756.715 217.210 ;
        RECT 757.005 217.040 757.175 217.210 ;
        RECT 757.465 217.040 757.635 217.210 ;
        RECT 757.925 217.040 758.095 217.210 ;
        RECT 758.385 217.040 758.555 217.210 ;
        RECT 759.765 217.040 759.935 217.210 ;
        RECT 760.225 217.040 760.395 217.210 ;
        RECT 760.685 217.040 760.855 217.210 ;
        RECT 761.145 217.040 761.315 217.210 ;
        RECT 761.605 217.040 761.775 217.210 ;
        RECT 762.065 217.040 762.235 217.210 ;
        RECT 762.525 217.040 762.695 217.210 ;
        RECT 762.985 217.040 763.155 217.210 ;
        RECT 763.445 217.040 763.615 217.210 ;
        RECT 763.905 217.040 764.075 217.210 ;
        RECT 764.365 217.040 764.535 217.210 ;
        RECT 765.745 217.040 765.915 217.210 ;
        RECT 766.205 217.040 766.375 217.210 ;
        RECT 766.665 217.040 766.835 217.210 ;
        RECT 767.125 217.040 767.295 217.210 ;
        RECT 767.585 217.040 767.755 217.210 ;
        RECT 768.045 217.040 768.215 217.210 ;
        RECT 768.505 217.040 768.675 217.210 ;
        RECT 768.965 217.040 769.135 217.210 ;
        RECT 769.425 217.040 769.595 217.210 ;
        RECT 769.885 217.040 770.055 217.210 ;
        RECT 770.345 217.040 770.515 217.210 ;
        RECT 771.725 217.040 771.895 217.210 ;
        RECT 772.185 217.040 772.355 217.210 ;
        RECT 772.645 217.040 772.815 217.210 ;
        RECT 773.105 217.040 773.275 217.210 ;
        RECT 773.565 217.040 773.735 217.210 ;
        RECT 774.025 217.040 774.195 217.210 ;
        RECT 774.485 217.040 774.655 217.210 ;
        RECT 774.945 217.040 775.115 217.210 ;
        RECT 775.405 217.040 775.575 217.210 ;
        RECT 775.865 217.040 776.035 217.210 ;
        RECT 776.325 217.040 776.495 217.210 ;
        RECT 777.705 217.040 777.875 217.210 ;
        RECT 778.165 217.040 778.335 217.210 ;
        RECT 778.625 217.040 778.795 217.210 ;
        RECT 779.085 217.040 779.255 217.210 ;
        RECT 779.545 217.040 779.715 217.210 ;
        RECT 780.005 217.040 780.175 217.210 ;
        RECT 780.465 217.040 780.635 217.210 ;
        RECT 780.925 217.040 781.095 217.210 ;
        RECT 781.385 217.040 781.555 217.210 ;
        RECT 781.845 217.040 782.015 217.210 ;
        RECT 782.305 217.040 782.475 217.210 ;
        RECT 783.685 217.040 783.855 217.210 ;
        RECT 784.145 217.040 784.315 217.210 ;
        RECT 784.605 217.040 784.775 217.210 ;
        RECT 785.065 217.040 785.235 217.210 ;
        RECT 785.525 217.040 785.695 217.210 ;
        RECT 785.985 217.040 786.155 217.210 ;
        RECT 786.445 217.040 786.615 217.210 ;
        RECT 786.905 217.040 787.075 217.210 ;
        RECT 787.365 217.040 787.535 217.210 ;
        RECT 787.825 217.040 787.995 217.210 ;
        RECT 788.285 217.040 788.455 217.210 ;
        RECT 789.665 217.040 789.835 217.210 ;
        RECT 790.125 217.040 790.295 217.210 ;
        RECT 790.585 217.040 790.755 217.210 ;
        RECT 791.045 217.040 791.215 217.210 ;
        RECT 791.505 217.040 791.675 217.210 ;
        RECT 791.965 217.040 792.135 217.210 ;
        RECT 792.425 217.040 792.595 217.210 ;
        RECT 792.885 217.040 793.055 217.210 ;
        RECT 793.345 217.040 793.515 217.210 ;
        RECT 793.805 217.040 793.975 217.210 ;
        RECT 794.265 217.040 794.435 217.210 ;
        RECT 670.065 211.600 670.235 211.770 ;
        RECT 670.525 211.600 670.695 211.770 ;
        RECT 670.985 211.600 671.155 211.770 ;
        RECT 671.445 211.600 671.615 211.770 ;
        RECT 671.905 211.600 672.075 211.770 ;
        RECT 672.365 211.600 672.535 211.770 ;
        RECT 672.825 211.600 672.995 211.770 ;
        RECT 673.285 211.600 673.455 211.770 ;
        RECT 673.745 211.600 673.915 211.770 ;
        RECT 674.205 211.600 674.375 211.770 ;
        RECT 674.665 211.600 674.835 211.770 ;
      LAYER met1 ;
        RECT 669.000 216.885 795.040 217.365 ;
        RECT 669.000 211.445 795.040 211.925 ;
      LAYER via ;
        RECT 736.975 216.985 738.760 217.285 ;
        RECT 736.975 211.575 738.760 211.875 ;
      LAYER met2 ;
        RECT 736.935 216.915 738.800 217.345 ;
        RECT 736.935 211.490 738.800 211.920 ;
      LAYER via2 ;
        RECT 736.975 216.985 738.760 217.285 ;
        RECT 736.975 211.575 738.760 211.875 ;
      LAYER met3 ;
        RECT 736.940 209.835 738.805 217.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 2148.130 217.755 2148.470 218.585 ;
        RECT 2154.110 217.755 2154.450 218.585 ;
        RECT 2160.090 217.755 2160.430 218.585 ;
        RECT 2166.070 217.755 2166.410 218.585 ;
        RECT 2172.050 217.755 2172.390 218.585 ;
        RECT 2178.030 217.755 2178.370 218.585 ;
        RECT 2184.010 217.755 2184.350 218.585 ;
        RECT 2189.990 217.755 2190.330 218.585 ;
        RECT 2195.970 217.755 2196.310 218.585 ;
        RECT 2201.950 217.755 2202.290 218.585 ;
        RECT 2207.930 217.755 2208.270 218.585 ;
        RECT 2213.910 217.755 2214.250 218.585 ;
        RECT 2219.890 217.755 2220.230 218.585 ;
        RECT 2225.870 217.755 2226.210 218.585 ;
        RECT 2231.850 217.755 2232.190 218.585 ;
        RECT 2146.545 217.210 2151.890 217.755 ;
        RECT 2152.525 217.210 2157.870 217.755 ;
        RECT 2158.505 217.210 2163.850 217.755 ;
        RECT 2164.485 217.210 2169.830 217.755 ;
        RECT 2170.465 217.210 2175.810 217.755 ;
        RECT 2176.445 217.210 2181.790 217.755 ;
        RECT 2182.425 217.210 2187.770 217.755 ;
        RECT 2188.405 217.210 2193.750 217.755 ;
        RECT 2194.385 217.210 2199.730 217.755 ;
        RECT 2200.365 217.210 2205.710 217.755 ;
        RECT 2206.345 217.210 2211.690 217.755 ;
        RECT 2212.325 217.210 2217.670 217.755 ;
        RECT 2218.305 217.210 2223.650 217.755 ;
        RECT 2224.285 217.210 2229.630 217.755 ;
        RECT 2230.265 217.210 2235.610 217.755 ;
      LAYER li1 ;
        RECT 2146.145 217.040 2146.315 217.210 ;
      LAYER li1 ;
        RECT 2146.460 217.040 2146.605 217.210 ;
        RECT 2146.775 217.040 2151.980 217.210 ;
      LAYER li1 ;
        RECT 2152.125 217.040 2152.295 217.210 ;
      LAYER li1 ;
        RECT 2152.440 217.040 2152.585 217.210 ;
        RECT 2152.755 217.040 2157.960 217.210 ;
      LAYER li1 ;
        RECT 2158.105 217.040 2158.275 217.210 ;
      LAYER li1 ;
        RECT 2158.420 217.040 2158.565 217.210 ;
        RECT 2158.735 217.040 2163.940 217.210 ;
      LAYER li1 ;
        RECT 2164.085 217.040 2164.255 217.210 ;
      LAYER li1 ;
        RECT 2164.400 217.040 2164.545 217.210 ;
        RECT 2164.715 217.040 2169.920 217.210 ;
      LAYER li1 ;
        RECT 2170.065 217.040 2170.235 217.210 ;
      LAYER li1 ;
        RECT 2170.380 217.040 2170.525 217.210 ;
        RECT 2170.695 217.040 2175.900 217.210 ;
      LAYER li1 ;
        RECT 2176.045 217.040 2176.215 217.210 ;
      LAYER li1 ;
        RECT 2176.360 217.040 2176.505 217.210 ;
        RECT 2176.675 217.040 2181.880 217.210 ;
      LAYER li1 ;
        RECT 2182.025 217.040 2182.195 217.210 ;
      LAYER li1 ;
        RECT 2182.340 217.040 2182.485 217.210 ;
        RECT 2182.655 217.040 2187.860 217.210 ;
      LAYER li1 ;
        RECT 2188.005 217.040 2188.175 217.210 ;
      LAYER li1 ;
        RECT 2188.320 217.040 2188.465 217.210 ;
        RECT 2188.635 217.040 2193.840 217.210 ;
      LAYER li1 ;
        RECT 2193.985 217.040 2194.155 217.210 ;
      LAYER li1 ;
        RECT 2194.300 217.040 2194.445 217.210 ;
        RECT 2194.615 217.040 2199.820 217.210 ;
      LAYER li1 ;
        RECT 2199.965 217.040 2200.135 217.210 ;
      LAYER li1 ;
        RECT 2200.280 217.040 2200.425 217.210 ;
        RECT 2200.595 217.040 2205.800 217.210 ;
      LAYER li1 ;
        RECT 2205.945 217.040 2206.115 217.210 ;
      LAYER li1 ;
        RECT 2206.260 217.040 2206.405 217.210 ;
        RECT 2206.575 217.040 2211.780 217.210 ;
      LAYER li1 ;
        RECT 2211.925 217.040 2212.095 217.210 ;
      LAYER li1 ;
        RECT 2212.240 217.040 2212.385 217.210 ;
        RECT 2212.555 217.040 2217.760 217.210 ;
      LAYER li1 ;
        RECT 2217.905 217.040 2218.075 217.210 ;
      LAYER li1 ;
        RECT 2218.220 217.040 2218.365 217.210 ;
        RECT 2218.535 217.040 2223.740 217.210 ;
      LAYER li1 ;
        RECT 2223.885 217.040 2224.055 217.210 ;
      LAYER li1 ;
        RECT 2224.200 217.040 2224.345 217.210 ;
        RECT 2224.515 217.040 2229.720 217.210 ;
      LAYER li1 ;
        RECT 2229.865 217.040 2230.035 217.210 ;
      LAYER li1 ;
        RECT 2230.180 217.040 2230.325 217.210 ;
        RECT 2230.495 217.040 2235.700 217.210 ;
      LAYER li1 ;
        RECT 2235.845 217.040 2236.015 217.210 ;
        RECT 2236.305 217.040 2236.475 217.210 ;
        RECT 2236.765 217.040 2236.935 217.210 ;
        RECT 2237.225 217.040 2237.395 217.210 ;
        RECT 2237.685 217.040 2237.855 217.210 ;
        RECT 2238.145 217.040 2238.315 217.210 ;
        RECT 2238.605 217.040 2238.775 217.210 ;
        RECT 2239.065 217.040 2239.235 217.210 ;
        RECT 2239.525 217.040 2239.695 217.210 ;
        RECT 2239.985 217.040 2240.155 217.210 ;
        RECT 2240.445 217.040 2240.615 217.210 ;
        RECT 2240.905 217.040 2241.075 217.210 ;
        RECT 2241.365 217.040 2241.535 217.210 ;
        RECT 2241.825 217.040 2241.995 217.210 ;
        RECT 2242.285 217.040 2242.455 217.210 ;
        RECT 2242.745 217.040 2242.915 217.210 ;
        RECT 2243.205 217.040 2243.375 217.210 ;
        RECT 2243.665 217.040 2243.835 217.210 ;
        RECT 2244.125 217.040 2244.295 217.210 ;
        RECT 2244.585 217.040 2244.755 217.210 ;
        RECT 2245.045 217.040 2245.215 217.210 ;
        RECT 2245.505 217.040 2245.675 217.210 ;
        RECT 2245.965 217.040 2246.135 217.210 ;
        RECT 2246.425 217.040 2246.595 217.210 ;
        RECT 2246.885 217.040 2247.055 217.210 ;
        RECT 2247.345 217.040 2247.515 217.210 ;
        RECT 2247.805 217.040 2247.975 217.210 ;
        RECT 2248.265 217.040 2248.435 217.210 ;
        RECT 2248.725 217.040 2248.895 217.210 ;
        RECT 2249.185 217.040 2249.355 217.210 ;
        RECT 2249.645 217.040 2249.815 217.210 ;
        RECT 2250.105 217.040 2250.275 217.210 ;
        RECT 2250.565 217.040 2250.735 217.210 ;
        RECT 2251.025 217.040 2251.195 217.210 ;
        RECT 2251.485 217.040 2251.655 217.210 ;
        RECT 2251.945 217.040 2252.115 217.210 ;
        RECT 2252.405 217.040 2252.575 217.210 ;
        RECT 2252.865 217.040 2253.035 217.210 ;
        RECT 2253.325 217.040 2253.495 217.210 ;
        RECT 2253.785 217.040 2253.955 217.210 ;
        RECT 2254.245 217.040 2254.415 217.210 ;
        RECT 2254.705 217.040 2254.875 217.210 ;
        RECT 2255.165 217.040 2255.335 217.210 ;
        RECT 2255.625 217.040 2255.795 217.210 ;
        RECT 2256.085 217.040 2256.255 217.210 ;
        RECT 2256.545 217.040 2256.715 217.210 ;
        RECT 2257.005 217.040 2257.175 217.210 ;
        RECT 2257.465 217.040 2257.635 217.210 ;
        RECT 2257.925 217.040 2258.095 217.210 ;
        RECT 2258.385 217.040 2258.555 217.210 ;
        RECT 2258.845 217.040 2259.015 217.210 ;
        RECT 2259.305 217.040 2259.475 217.210 ;
        RECT 2259.765 217.040 2259.935 217.210 ;
        RECT 2260.225 217.040 2260.395 217.210 ;
        RECT 2260.685 217.040 2260.855 217.210 ;
        RECT 2261.145 217.040 2261.315 217.210 ;
        RECT 2261.605 217.040 2261.775 217.210 ;
        RECT 2262.065 217.040 2262.235 217.210 ;
        RECT 2262.525 217.040 2262.695 217.210 ;
        RECT 2262.985 217.040 2263.155 217.210 ;
        RECT 2263.445 217.040 2263.615 217.210 ;
        RECT 2263.905 217.040 2264.075 217.210 ;
        RECT 2264.365 217.040 2264.535 217.210 ;
        RECT 2264.825 217.040 2264.995 217.210 ;
        RECT 2265.285 217.040 2265.455 217.210 ;
        RECT 2265.745 217.040 2265.915 217.210 ;
        RECT 2266.205 217.040 2266.375 217.210 ;
        RECT 2266.665 217.040 2266.835 217.210 ;
        RECT 2267.125 217.040 2267.295 217.210 ;
        RECT 2267.585 217.040 2267.755 217.210 ;
        RECT 2268.045 217.040 2268.215 217.210 ;
        RECT 2268.505 217.040 2268.675 217.210 ;
        RECT 2268.965 217.040 2269.135 217.210 ;
        RECT 2269.425 217.040 2269.595 217.210 ;
        RECT 2269.885 217.040 2270.055 217.210 ;
        RECT 2270.345 217.040 2270.515 217.210 ;
        RECT 2270.805 217.040 2270.975 217.210 ;
        RECT 2271.265 217.040 2271.435 217.210 ;
        RECT 2271.725 217.040 2271.895 217.210 ;
      LAYER li1 ;
        RECT 2148.130 212.315 2148.470 213.145 ;
        RECT 2146.545 211.770 2151.890 212.315 ;
      LAYER li1 ;
        RECT 2146.145 211.600 2146.315 211.770 ;
      LAYER li1 ;
        RECT 2146.460 211.600 2151.980 211.770 ;
      LAYER li1 ;
        RECT 2152.125 211.600 2152.295 211.770 ;
        RECT 2152.585 211.600 2152.755 211.770 ;
        RECT 2153.045 211.600 2153.215 211.770 ;
        RECT 2153.505 211.600 2153.675 211.770 ;
        RECT 2153.965 211.600 2154.135 211.770 ;
        RECT 2154.425 211.600 2154.595 211.770 ;
        RECT 2154.885 211.600 2155.055 211.770 ;
        RECT 2155.345 211.600 2155.515 211.770 ;
        RECT 2155.805 211.600 2155.975 211.770 ;
        RECT 2156.265 211.600 2156.435 211.770 ;
        RECT 2156.725 211.600 2156.895 211.770 ;
        RECT 2157.185 211.600 2157.355 211.770 ;
        RECT 2157.645 211.600 2157.815 211.770 ;
        RECT 2158.105 211.600 2158.275 211.770 ;
        RECT 2158.565 211.600 2158.735 211.770 ;
        RECT 2159.025 211.600 2159.195 211.770 ;
        RECT 2159.485 211.600 2159.655 211.770 ;
        RECT 2159.945 211.600 2160.115 211.770 ;
        RECT 2160.405 211.600 2160.575 211.770 ;
        RECT 2160.865 211.600 2161.035 211.770 ;
        RECT 2161.325 211.600 2161.495 211.770 ;
        RECT 2161.785 211.600 2161.955 211.770 ;
        RECT 2162.245 211.600 2162.415 211.770 ;
        RECT 2162.705 211.600 2162.875 211.770 ;
        RECT 2163.165 211.600 2163.335 211.770 ;
        RECT 2163.625 211.600 2163.795 211.770 ;
        RECT 2164.085 211.600 2164.255 211.770 ;
        RECT 2164.545 211.600 2164.715 211.770 ;
        RECT 2165.005 211.600 2165.175 211.770 ;
        RECT 2165.465 211.600 2165.635 211.770 ;
        RECT 2165.925 211.600 2166.095 211.770 ;
        RECT 2166.385 211.600 2166.555 211.770 ;
        RECT 2166.845 211.600 2167.015 211.770 ;
        RECT 2167.305 211.600 2167.475 211.770 ;
        RECT 2167.765 211.600 2167.935 211.770 ;
        RECT 2168.225 211.600 2168.395 211.770 ;
        RECT 2168.685 211.600 2168.855 211.770 ;
        RECT 2169.145 211.600 2169.315 211.770 ;
        RECT 2169.605 211.600 2169.775 211.770 ;
        RECT 2170.065 211.600 2170.235 211.770 ;
        RECT 2170.525 211.600 2170.695 211.770 ;
        RECT 2170.985 211.600 2171.155 211.770 ;
        RECT 2171.445 211.600 2171.615 211.770 ;
        RECT 2171.905 211.600 2172.075 211.770 ;
        RECT 2172.365 211.600 2172.535 211.770 ;
        RECT 2172.825 211.600 2172.995 211.770 ;
        RECT 2173.285 211.600 2173.455 211.770 ;
        RECT 2173.745 211.600 2173.915 211.770 ;
        RECT 2174.205 211.600 2174.375 211.770 ;
        RECT 2174.665 211.600 2174.835 211.770 ;
        RECT 2175.125 211.600 2175.295 211.770 ;
        RECT 2175.585 211.600 2175.755 211.770 ;
        RECT 2176.045 211.600 2176.215 211.770 ;
        RECT 2176.505 211.600 2176.675 211.770 ;
        RECT 2176.965 211.600 2177.135 211.770 ;
        RECT 2177.425 211.600 2177.595 211.770 ;
        RECT 2177.885 211.600 2178.055 211.770 ;
        RECT 2178.345 211.600 2178.515 211.770 ;
        RECT 2178.805 211.600 2178.975 211.770 ;
        RECT 2179.265 211.600 2179.435 211.770 ;
        RECT 2179.725 211.600 2179.895 211.770 ;
        RECT 2180.185 211.600 2180.355 211.770 ;
        RECT 2180.645 211.600 2180.815 211.770 ;
        RECT 2181.105 211.600 2181.275 211.770 ;
        RECT 2181.565 211.600 2181.735 211.770 ;
        RECT 2182.025 211.600 2182.195 211.770 ;
        RECT 2182.485 211.600 2182.655 211.770 ;
        RECT 2182.945 211.600 2183.115 211.770 ;
        RECT 2183.405 211.600 2183.575 211.770 ;
        RECT 2183.865 211.600 2184.035 211.770 ;
        RECT 2184.325 211.600 2184.495 211.770 ;
        RECT 2184.785 211.600 2184.955 211.770 ;
        RECT 2185.245 211.600 2185.415 211.770 ;
        RECT 2185.705 211.600 2185.875 211.770 ;
        RECT 2186.165 211.600 2186.335 211.770 ;
        RECT 2186.625 211.600 2186.795 211.770 ;
        RECT 2187.085 211.600 2187.255 211.770 ;
        RECT 2187.545 211.600 2187.715 211.770 ;
        RECT 2188.005 211.600 2188.175 211.770 ;
        RECT 2188.465 211.600 2188.635 211.770 ;
        RECT 2188.925 211.600 2189.095 211.770 ;
        RECT 2189.385 211.600 2189.555 211.770 ;
        RECT 2189.845 211.600 2190.015 211.770 ;
        RECT 2190.305 211.600 2190.475 211.770 ;
        RECT 2190.765 211.600 2190.935 211.770 ;
        RECT 2191.225 211.600 2191.395 211.770 ;
        RECT 2191.685 211.600 2191.855 211.770 ;
        RECT 2192.145 211.600 2192.315 211.770 ;
        RECT 2192.605 211.600 2192.775 211.770 ;
        RECT 2193.065 211.600 2193.235 211.770 ;
        RECT 2193.525 211.600 2193.695 211.770 ;
        RECT 2193.985 211.600 2194.155 211.770 ;
        RECT 2194.445 211.600 2194.615 211.770 ;
        RECT 2194.905 211.600 2195.075 211.770 ;
        RECT 2195.365 211.600 2195.535 211.770 ;
        RECT 2195.825 211.600 2195.995 211.770 ;
        RECT 2196.285 211.600 2196.455 211.770 ;
        RECT 2196.745 211.600 2196.915 211.770 ;
        RECT 2197.205 211.600 2197.375 211.770 ;
        RECT 2197.665 211.600 2197.835 211.770 ;
        RECT 2198.125 211.600 2198.295 211.770 ;
        RECT 2198.585 211.600 2198.755 211.770 ;
        RECT 2199.045 211.600 2199.215 211.770 ;
        RECT 2199.505 211.600 2199.675 211.770 ;
        RECT 2199.965 211.600 2200.135 211.770 ;
        RECT 2200.425 211.600 2200.595 211.770 ;
        RECT 2200.885 211.600 2201.055 211.770 ;
        RECT 2201.345 211.600 2201.515 211.770 ;
        RECT 2201.805 211.600 2201.975 211.770 ;
        RECT 2202.265 211.600 2202.435 211.770 ;
        RECT 2202.725 211.600 2202.895 211.770 ;
        RECT 2203.185 211.600 2203.355 211.770 ;
        RECT 2203.645 211.600 2203.815 211.770 ;
        RECT 2204.105 211.600 2204.275 211.770 ;
        RECT 2204.565 211.600 2204.735 211.770 ;
        RECT 2205.025 211.600 2205.195 211.770 ;
        RECT 2205.485 211.600 2205.655 211.770 ;
        RECT 2205.945 211.600 2206.115 211.770 ;
        RECT 2206.405 211.600 2206.575 211.770 ;
        RECT 2206.865 211.600 2207.035 211.770 ;
        RECT 2207.325 211.600 2207.495 211.770 ;
        RECT 2207.785 211.600 2207.955 211.770 ;
        RECT 2208.245 211.600 2208.415 211.770 ;
        RECT 2208.705 211.600 2208.875 211.770 ;
        RECT 2209.165 211.600 2209.335 211.770 ;
        RECT 2209.625 211.600 2209.795 211.770 ;
        RECT 2210.085 211.600 2210.255 211.770 ;
        RECT 2210.545 211.600 2210.715 211.770 ;
        RECT 2211.005 211.600 2211.175 211.770 ;
        RECT 2211.465 211.600 2211.635 211.770 ;
        RECT 2211.925 211.600 2212.095 211.770 ;
        RECT 2212.385 211.600 2212.555 211.770 ;
        RECT 2212.845 211.600 2213.015 211.770 ;
        RECT 2213.305 211.600 2213.475 211.770 ;
        RECT 2213.765 211.600 2213.935 211.770 ;
        RECT 2214.225 211.600 2214.395 211.770 ;
        RECT 2214.685 211.600 2214.855 211.770 ;
        RECT 2215.145 211.600 2215.315 211.770 ;
        RECT 2215.605 211.600 2215.775 211.770 ;
        RECT 2216.065 211.600 2216.235 211.770 ;
        RECT 2216.525 211.600 2216.695 211.770 ;
        RECT 2216.985 211.600 2217.155 211.770 ;
        RECT 2217.445 211.600 2217.615 211.770 ;
        RECT 2217.905 211.600 2218.075 211.770 ;
        RECT 2218.365 211.600 2218.535 211.770 ;
        RECT 2218.825 211.600 2218.995 211.770 ;
        RECT 2219.285 211.600 2219.455 211.770 ;
        RECT 2219.745 211.600 2219.915 211.770 ;
        RECT 2220.205 211.600 2220.375 211.770 ;
        RECT 2220.665 211.600 2220.835 211.770 ;
        RECT 2221.125 211.600 2221.295 211.770 ;
        RECT 2221.585 211.600 2221.755 211.770 ;
        RECT 2222.045 211.600 2222.215 211.770 ;
        RECT 2222.505 211.600 2222.675 211.770 ;
        RECT 2222.965 211.600 2223.135 211.770 ;
        RECT 2223.425 211.600 2223.595 211.770 ;
        RECT 2223.885 211.600 2224.055 211.770 ;
        RECT 2224.345 211.600 2224.515 211.770 ;
        RECT 2224.805 211.600 2224.975 211.770 ;
        RECT 2225.265 211.600 2225.435 211.770 ;
        RECT 2225.725 211.600 2225.895 211.770 ;
        RECT 2226.185 211.600 2226.355 211.770 ;
        RECT 2226.645 211.600 2226.815 211.770 ;
        RECT 2227.105 211.600 2227.275 211.770 ;
        RECT 2227.565 211.600 2227.735 211.770 ;
        RECT 2228.025 211.600 2228.195 211.770 ;
        RECT 2228.485 211.600 2228.655 211.770 ;
        RECT 2228.945 211.600 2229.115 211.770 ;
        RECT 2229.405 211.600 2229.575 211.770 ;
        RECT 2229.865 211.600 2230.035 211.770 ;
        RECT 2230.325 211.600 2230.495 211.770 ;
        RECT 2230.785 211.600 2230.955 211.770 ;
        RECT 2231.245 211.600 2231.415 211.770 ;
        RECT 2231.705 211.600 2231.875 211.770 ;
        RECT 2232.165 211.600 2232.335 211.770 ;
        RECT 2232.625 211.600 2232.795 211.770 ;
        RECT 2233.085 211.600 2233.255 211.770 ;
        RECT 2233.545 211.600 2233.715 211.770 ;
        RECT 2234.005 211.600 2234.175 211.770 ;
        RECT 2234.465 211.600 2234.635 211.770 ;
        RECT 2234.925 211.600 2235.095 211.770 ;
        RECT 2235.385 211.600 2235.555 211.770 ;
        RECT 2235.845 211.600 2236.015 211.770 ;
        RECT 2236.305 211.600 2236.475 211.770 ;
        RECT 2236.765 211.600 2236.935 211.770 ;
        RECT 2237.225 211.600 2237.395 211.770 ;
        RECT 2237.685 211.600 2237.855 211.770 ;
        RECT 2238.145 211.600 2238.315 211.770 ;
        RECT 2238.605 211.600 2238.775 211.770 ;
        RECT 2239.065 211.600 2239.235 211.770 ;
        RECT 2239.525 211.600 2239.695 211.770 ;
        RECT 2239.985 211.600 2240.155 211.770 ;
        RECT 2240.445 211.600 2240.615 211.770 ;
        RECT 2240.905 211.600 2241.075 211.770 ;
        RECT 2241.365 211.600 2241.535 211.770 ;
        RECT 2241.825 211.600 2241.995 211.770 ;
        RECT 2242.285 211.600 2242.455 211.770 ;
        RECT 2242.745 211.600 2242.915 211.770 ;
        RECT 2243.205 211.600 2243.375 211.770 ;
        RECT 2243.665 211.600 2243.835 211.770 ;
        RECT 2244.125 211.600 2244.295 211.770 ;
        RECT 2244.585 211.600 2244.755 211.770 ;
        RECT 2245.045 211.600 2245.215 211.770 ;
        RECT 2245.505 211.600 2245.675 211.770 ;
        RECT 2245.965 211.600 2246.135 211.770 ;
        RECT 2246.425 211.600 2246.595 211.770 ;
        RECT 2246.885 211.600 2247.055 211.770 ;
        RECT 2247.345 211.600 2247.515 211.770 ;
        RECT 2247.805 211.600 2247.975 211.770 ;
        RECT 2248.265 211.600 2248.435 211.770 ;
        RECT 2248.725 211.600 2248.895 211.770 ;
        RECT 2249.185 211.600 2249.355 211.770 ;
        RECT 2249.645 211.600 2249.815 211.770 ;
        RECT 2250.105 211.600 2250.275 211.770 ;
        RECT 2250.565 211.600 2250.735 211.770 ;
        RECT 2251.025 211.600 2251.195 211.770 ;
        RECT 2251.485 211.600 2251.655 211.770 ;
        RECT 2251.945 211.600 2252.115 211.770 ;
        RECT 2252.405 211.600 2252.575 211.770 ;
        RECT 2252.865 211.600 2253.035 211.770 ;
        RECT 2253.325 211.600 2253.495 211.770 ;
        RECT 2253.785 211.600 2253.955 211.770 ;
        RECT 2254.245 211.600 2254.415 211.770 ;
        RECT 2254.705 211.600 2254.875 211.770 ;
        RECT 2255.165 211.600 2255.335 211.770 ;
        RECT 2255.625 211.600 2255.795 211.770 ;
        RECT 2256.085 211.600 2256.255 211.770 ;
        RECT 2256.545 211.600 2256.715 211.770 ;
        RECT 2257.005 211.600 2257.175 211.770 ;
        RECT 2257.465 211.600 2257.635 211.770 ;
        RECT 2257.925 211.600 2258.095 211.770 ;
        RECT 2258.385 211.600 2258.555 211.770 ;
        RECT 2258.845 211.600 2259.015 211.770 ;
        RECT 2259.305 211.600 2259.475 211.770 ;
        RECT 2259.765 211.600 2259.935 211.770 ;
        RECT 2260.225 211.600 2260.395 211.770 ;
        RECT 2260.685 211.600 2260.855 211.770 ;
        RECT 2261.145 211.600 2261.315 211.770 ;
        RECT 2261.605 211.600 2261.775 211.770 ;
        RECT 2262.065 211.600 2262.235 211.770 ;
        RECT 2262.525 211.600 2262.695 211.770 ;
        RECT 2262.985 211.600 2263.155 211.770 ;
        RECT 2263.445 211.600 2263.615 211.770 ;
        RECT 2263.905 211.600 2264.075 211.770 ;
        RECT 2264.365 211.600 2264.535 211.770 ;
        RECT 2264.825 211.600 2264.995 211.770 ;
        RECT 2265.285 211.600 2265.455 211.770 ;
        RECT 2265.745 211.600 2265.915 211.770 ;
        RECT 2266.205 211.600 2266.375 211.770 ;
        RECT 2266.665 211.600 2266.835 211.770 ;
        RECT 2267.125 211.600 2267.295 211.770 ;
        RECT 2267.585 211.600 2267.755 211.770 ;
        RECT 2268.045 211.600 2268.215 211.770 ;
        RECT 2268.505 211.600 2268.675 211.770 ;
        RECT 2268.965 211.600 2269.135 211.770 ;
        RECT 2269.425 211.600 2269.595 211.770 ;
        RECT 2269.885 211.600 2270.055 211.770 ;
        RECT 2270.345 211.600 2270.515 211.770 ;
        RECT 2270.805 211.600 2270.975 211.770 ;
        RECT 2271.265 211.600 2271.435 211.770 ;
        RECT 2271.725 211.600 2271.895 211.770 ;
      LAYER mcon ;
        RECT 2147.065 217.040 2147.235 217.210 ;
        RECT 2147.525 217.040 2147.695 217.210 ;
        RECT 2147.985 217.040 2148.155 217.210 ;
        RECT 2148.445 217.040 2148.615 217.210 ;
        RECT 2148.905 217.040 2149.075 217.210 ;
        RECT 2149.365 217.040 2149.535 217.210 ;
        RECT 2149.825 217.040 2149.995 217.210 ;
        RECT 2150.285 217.040 2150.455 217.210 ;
        RECT 2150.745 217.040 2150.915 217.210 ;
        RECT 2151.205 217.040 2151.375 217.210 ;
        RECT 2151.665 217.040 2151.835 217.210 ;
        RECT 2153.045 217.040 2153.215 217.210 ;
        RECT 2153.505 217.040 2153.675 217.210 ;
        RECT 2153.965 217.040 2154.135 217.210 ;
        RECT 2154.425 217.040 2154.595 217.210 ;
        RECT 2154.885 217.040 2155.055 217.210 ;
        RECT 2155.345 217.040 2155.515 217.210 ;
        RECT 2155.805 217.040 2155.975 217.210 ;
        RECT 2156.265 217.040 2156.435 217.210 ;
        RECT 2156.725 217.040 2156.895 217.210 ;
        RECT 2157.185 217.040 2157.355 217.210 ;
        RECT 2157.645 217.040 2157.815 217.210 ;
        RECT 2159.025 217.040 2159.195 217.210 ;
        RECT 2159.485 217.040 2159.655 217.210 ;
        RECT 2159.945 217.040 2160.115 217.210 ;
        RECT 2160.405 217.040 2160.575 217.210 ;
        RECT 2160.865 217.040 2161.035 217.210 ;
        RECT 2161.325 217.040 2161.495 217.210 ;
        RECT 2161.785 217.040 2161.955 217.210 ;
        RECT 2162.245 217.040 2162.415 217.210 ;
        RECT 2162.705 217.040 2162.875 217.210 ;
        RECT 2163.165 217.040 2163.335 217.210 ;
        RECT 2163.625 217.040 2163.795 217.210 ;
        RECT 2165.005 217.040 2165.175 217.210 ;
        RECT 2165.465 217.040 2165.635 217.210 ;
        RECT 2165.925 217.040 2166.095 217.210 ;
        RECT 2166.385 217.040 2166.555 217.210 ;
        RECT 2166.845 217.040 2167.015 217.210 ;
        RECT 2167.305 217.040 2167.475 217.210 ;
        RECT 2167.765 217.040 2167.935 217.210 ;
        RECT 2168.225 217.040 2168.395 217.210 ;
        RECT 2168.685 217.040 2168.855 217.210 ;
        RECT 2169.145 217.040 2169.315 217.210 ;
        RECT 2169.605 217.040 2169.775 217.210 ;
        RECT 2170.985 217.040 2171.155 217.210 ;
        RECT 2171.445 217.040 2171.615 217.210 ;
        RECT 2171.905 217.040 2172.075 217.210 ;
        RECT 2172.365 217.040 2172.535 217.210 ;
        RECT 2172.825 217.040 2172.995 217.210 ;
        RECT 2173.285 217.040 2173.455 217.210 ;
        RECT 2173.745 217.040 2173.915 217.210 ;
        RECT 2174.205 217.040 2174.375 217.210 ;
        RECT 2174.665 217.040 2174.835 217.210 ;
        RECT 2175.125 217.040 2175.295 217.210 ;
        RECT 2175.585 217.040 2175.755 217.210 ;
        RECT 2176.965 217.040 2177.135 217.210 ;
        RECT 2177.425 217.040 2177.595 217.210 ;
        RECT 2177.885 217.040 2178.055 217.210 ;
        RECT 2178.345 217.040 2178.515 217.210 ;
        RECT 2178.805 217.040 2178.975 217.210 ;
        RECT 2179.265 217.040 2179.435 217.210 ;
        RECT 2179.725 217.040 2179.895 217.210 ;
        RECT 2180.185 217.040 2180.355 217.210 ;
        RECT 2180.645 217.040 2180.815 217.210 ;
        RECT 2181.105 217.040 2181.275 217.210 ;
        RECT 2181.565 217.040 2181.735 217.210 ;
        RECT 2182.945 217.040 2183.115 217.210 ;
        RECT 2183.405 217.040 2183.575 217.210 ;
        RECT 2183.865 217.040 2184.035 217.210 ;
        RECT 2184.325 217.040 2184.495 217.210 ;
        RECT 2184.785 217.040 2184.955 217.210 ;
        RECT 2185.245 217.040 2185.415 217.210 ;
        RECT 2185.705 217.040 2185.875 217.210 ;
        RECT 2186.165 217.040 2186.335 217.210 ;
        RECT 2186.625 217.040 2186.795 217.210 ;
        RECT 2187.085 217.040 2187.255 217.210 ;
        RECT 2187.545 217.040 2187.715 217.210 ;
        RECT 2188.925 217.040 2189.095 217.210 ;
        RECT 2189.385 217.040 2189.555 217.210 ;
        RECT 2189.845 217.040 2190.015 217.210 ;
        RECT 2190.305 217.040 2190.475 217.210 ;
        RECT 2190.765 217.040 2190.935 217.210 ;
        RECT 2191.225 217.040 2191.395 217.210 ;
        RECT 2191.685 217.040 2191.855 217.210 ;
        RECT 2192.145 217.040 2192.315 217.210 ;
        RECT 2192.605 217.040 2192.775 217.210 ;
        RECT 2193.065 217.040 2193.235 217.210 ;
        RECT 2193.525 217.040 2193.695 217.210 ;
        RECT 2194.905 217.040 2195.075 217.210 ;
        RECT 2195.365 217.040 2195.535 217.210 ;
        RECT 2195.825 217.040 2195.995 217.210 ;
        RECT 2196.285 217.040 2196.455 217.210 ;
        RECT 2196.745 217.040 2196.915 217.210 ;
        RECT 2197.205 217.040 2197.375 217.210 ;
        RECT 2197.665 217.040 2197.835 217.210 ;
        RECT 2198.125 217.040 2198.295 217.210 ;
        RECT 2198.585 217.040 2198.755 217.210 ;
        RECT 2199.045 217.040 2199.215 217.210 ;
        RECT 2199.505 217.040 2199.675 217.210 ;
        RECT 2200.885 217.040 2201.055 217.210 ;
        RECT 2201.345 217.040 2201.515 217.210 ;
        RECT 2201.805 217.040 2201.975 217.210 ;
        RECT 2202.265 217.040 2202.435 217.210 ;
        RECT 2202.725 217.040 2202.895 217.210 ;
        RECT 2203.185 217.040 2203.355 217.210 ;
        RECT 2203.645 217.040 2203.815 217.210 ;
        RECT 2204.105 217.040 2204.275 217.210 ;
        RECT 2204.565 217.040 2204.735 217.210 ;
        RECT 2205.025 217.040 2205.195 217.210 ;
        RECT 2205.485 217.040 2205.655 217.210 ;
        RECT 2206.865 217.040 2207.035 217.210 ;
        RECT 2207.325 217.040 2207.495 217.210 ;
        RECT 2207.785 217.040 2207.955 217.210 ;
        RECT 2208.245 217.040 2208.415 217.210 ;
        RECT 2208.705 217.040 2208.875 217.210 ;
        RECT 2209.165 217.040 2209.335 217.210 ;
        RECT 2209.625 217.040 2209.795 217.210 ;
        RECT 2210.085 217.040 2210.255 217.210 ;
        RECT 2210.545 217.040 2210.715 217.210 ;
        RECT 2211.005 217.040 2211.175 217.210 ;
        RECT 2211.465 217.040 2211.635 217.210 ;
        RECT 2212.845 217.040 2213.015 217.210 ;
        RECT 2213.305 217.040 2213.475 217.210 ;
        RECT 2213.765 217.040 2213.935 217.210 ;
        RECT 2214.225 217.040 2214.395 217.210 ;
        RECT 2214.685 217.040 2214.855 217.210 ;
        RECT 2215.145 217.040 2215.315 217.210 ;
        RECT 2215.605 217.040 2215.775 217.210 ;
        RECT 2216.065 217.040 2216.235 217.210 ;
        RECT 2216.525 217.040 2216.695 217.210 ;
        RECT 2216.985 217.040 2217.155 217.210 ;
        RECT 2217.445 217.040 2217.615 217.210 ;
        RECT 2218.825 217.040 2218.995 217.210 ;
        RECT 2219.285 217.040 2219.455 217.210 ;
        RECT 2219.745 217.040 2219.915 217.210 ;
        RECT 2220.205 217.040 2220.375 217.210 ;
        RECT 2220.665 217.040 2220.835 217.210 ;
        RECT 2221.125 217.040 2221.295 217.210 ;
        RECT 2221.585 217.040 2221.755 217.210 ;
        RECT 2222.045 217.040 2222.215 217.210 ;
        RECT 2222.505 217.040 2222.675 217.210 ;
        RECT 2222.965 217.040 2223.135 217.210 ;
        RECT 2223.425 217.040 2223.595 217.210 ;
        RECT 2224.805 217.040 2224.975 217.210 ;
        RECT 2225.265 217.040 2225.435 217.210 ;
        RECT 2225.725 217.040 2225.895 217.210 ;
        RECT 2226.185 217.040 2226.355 217.210 ;
        RECT 2226.645 217.040 2226.815 217.210 ;
        RECT 2227.105 217.040 2227.275 217.210 ;
        RECT 2227.565 217.040 2227.735 217.210 ;
        RECT 2228.025 217.040 2228.195 217.210 ;
        RECT 2228.485 217.040 2228.655 217.210 ;
        RECT 2228.945 217.040 2229.115 217.210 ;
        RECT 2229.405 217.040 2229.575 217.210 ;
        RECT 2230.785 217.040 2230.955 217.210 ;
        RECT 2231.245 217.040 2231.415 217.210 ;
        RECT 2231.705 217.040 2231.875 217.210 ;
        RECT 2232.165 217.040 2232.335 217.210 ;
        RECT 2232.625 217.040 2232.795 217.210 ;
        RECT 2233.085 217.040 2233.255 217.210 ;
        RECT 2233.545 217.040 2233.715 217.210 ;
        RECT 2234.005 217.040 2234.175 217.210 ;
        RECT 2234.465 217.040 2234.635 217.210 ;
        RECT 2234.925 217.040 2235.095 217.210 ;
        RECT 2235.385 217.040 2235.555 217.210 ;
        RECT 2147.065 211.600 2147.235 211.770 ;
        RECT 2147.525 211.600 2147.695 211.770 ;
        RECT 2147.985 211.600 2148.155 211.770 ;
        RECT 2148.445 211.600 2148.615 211.770 ;
        RECT 2148.905 211.600 2149.075 211.770 ;
        RECT 2149.365 211.600 2149.535 211.770 ;
        RECT 2149.825 211.600 2149.995 211.770 ;
        RECT 2150.285 211.600 2150.455 211.770 ;
        RECT 2150.745 211.600 2150.915 211.770 ;
        RECT 2151.205 211.600 2151.375 211.770 ;
        RECT 2151.665 211.600 2151.835 211.770 ;
      LAYER met1 ;
        RECT 2146.000 216.885 2272.040 217.365 ;
        RECT 2146.000 211.445 2272.040 211.925 ;
      LAYER via ;
        RECT 2208.130 216.950 2209.915 217.250 ;
        RECT 2208.130 211.540 2209.915 211.840 ;
      LAYER met2 ;
        RECT 2208.090 216.880 2209.955 217.310 ;
        RECT 2208.090 211.455 2209.955 211.885 ;
      LAYER via2 ;
        RECT 2208.130 216.950 2209.915 217.250 ;
        RECT 2208.130 211.540 2209.915 211.840 ;
      LAYER met3 ;
        RECT 2208.095 209.800 2209.960 217.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.995 1762.750 202.165 1762.920 ;
        RECT 207.435 1762.750 207.605 1762.920 ;
      LAYER li1 ;
        RECT 207.435 1762.520 207.605 1762.605 ;
        RECT 207.435 1762.460 208.150 1762.520 ;
      LAYER li1 ;
        RECT 201.995 1762.290 202.165 1762.460 ;
      LAYER li1 ;
        RECT 207.605 1762.290 208.150 1762.460 ;
      LAYER li1 ;
        RECT 201.995 1761.830 202.165 1762.000 ;
        RECT 201.995 1761.370 202.165 1761.540 ;
        RECT 201.995 1760.910 202.165 1761.080 ;
      LAYER li1 ;
        RECT 207.435 1760.935 208.150 1762.290 ;
      LAYER li1 ;
        RECT 201.995 1760.450 202.165 1760.620 ;
      LAYER li1 ;
        RECT 207.435 1760.595 208.980 1760.935 ;
      LAYER li1 ;
        RECT 201.995 1759.990 202.165 1760.160 ;
        RECT 201.995 1759.530 202.165 1759.700 ;
        RECT 201.995 1759.070 202.165 1759.240 ;
        RECT 201.995 1758.610 202.165 1758.780 ;
        RECT 201.995 1758.150 202.165 1758.320 ;
        RECT 201.995 1757.690 202.165 1757.860 ;
        RECT 201.995 1757.230 202.165 1757.400 ;
      LAYER li1 ;
        RECT 207.435 1757.175 208.150 1760.595 ;
        RECT 207.435 1757.085 207.605 1757.175 ;
      LAYER li1 ;
        RECT 201.995 1756.770 202.165 1756.940 ;
        RECT 207.435 1756.770 207.605 1756.940 ;
      LAYER li1 ;
        RECT 207.435 1756.540 207.605 1756.625 ;
        RECT 207.435 1756.480 208.150 1756.540 ;
      LAYER li1 ;
        RECT 201.995 1756.310 202.165 1756.480 ;
      LAYER li1 ;
        RECT 207.605 1756.310 208.150 1756.480 ;
      LAYER li1 ;
        RECT 201.995 1755.850 202.165 1756.020 ;
        RECT 201.995 1755.390 202.165 1755.560 ;
        RECT 201.995 1754.930 202.165 1755.100 ;
      LAYER li1 ;
        RECT 207.435 1754.955 208.150 1756.310 ;
      LAYER li1 ;
        RECT 201.995 1754.470 202.165 1754.640 ;
      LAYER li1 ;
        RECT 207.435 1754.615 208.980 1754.955 ;
      LAYER li1 ;
        RECT 201.995 1754.010 202.165 1754.180 ;
        RECT 201.995 1753.550 202.165 1753.720 ;
        RECT 201.995 1753.090 202.165 1753.260 ;
        RECT 201.995 1752.630 202.165 1752.800 ;
        RECT 201.995 1752.170 202.165 1752.340 ;
        RECT 201.995 1751.710 202.165 1751.880 ;
        RECT 201.995 1751.250 202.165 1751.420 ;
      LAYER li1 ;
        RECT 207.435 1751.195 208.150 1754.615 ;
        RECT 207.435 1751.105 207.605 1751.195 ;
      LAYER li1 ;
        RECT 201.995 1750.790 202.165 1750.960 ;
        RECT 207.435 1750.790 207.605 1750.960 ;
        RECT 201.995 1750.330 202.165 1750.500 ;
        RECT 207.435 1750.330 207.605 1750.500 ;
        RECT 201.995 1749.870 202.165 1750.040 ;
        RECT 207.435 1749.870 207.605 1750.040 ;
        RECT 201.995 1749.410 202.165 1749.580 ;
        RECT 207.435 1749.410 207.605 1749.580 ;
        RECT 201.995 1748.950 202.165 1749.120 ;
        RECT 207.435 1748.950 207.605 1749.120 ;
        RECT 201.995 1748.490 202.165 1748.660 ;
        RECT 207.435 1748.490 207.605 1748.660 ;
        RECT 201.995 1748.030 202.165 1748.200 ;
        RECT 207.435 1748.030 207.605 1748.200 ;
        RECT 201.995 1747.570 202.165 1747.740 ;
        RECT 207.435 1747.570 207.605 1747.740 ;
        RECT 201.995 1747.110 202.165 1747.280 ;
        RECT 207.435 1747.110 207.605 1747.280 ;
        RECT 201.995 1746.650 202.165 1746.820 ;
        RECT 207.435 1746.650 207.605 1746.820 ;
        RECT 201.995 1746.190 202.165 1746.360 ;
        RECT 207.435 1746.190 207.605 1746.360 ;
        RECT 201.995 1745.730 202.165 1745.900 ;
        RECT 207.435 1745.730 207.605 1745.900 ;
        RECT 201.995 1745.270 202.165 1745.440 ;
        RECT 207.435 1745.270 207.605 1745.440 ;
        RECT 201.995 1744.810 202.165 1744.980 ;
        RECT 207.435 1744.810 207.605 1744.980 ;
      LAYER li1 ;
        RECT 207.435 1744.580 207.605 1744.665 ;
        RECT 207.435 1744.520 208.150 1744.580 ;
      LAYER li1 ;
        RECT 201.995 1744.350 202.165 1744.520 ;
      LAYER li1 ;
        RECT 207.605 1744.350 208.150 1744.520 ;
      LAYER li1 ;
        RECT 201.995 1743.890 202.165 1744.060 ;
        RECT 201.995 1743.430 202.165 1743.600 ;
        RECT 201.995 1742.970 202.165 1743.140 ;
      LAYER li1 ;
        RECT 207.435 1742.995 208.150 1744.350 ;
      LAYER li1 ;
        RECT 201.995 1742.510 202.165 1742.680 ;
      LAYER li1 ;
        RECT 207.435 1742.655 208.980 1742.995 ;
      LAYER li1 ;
        RECT 201.995 1742.050 202.165 1742.220 ;
        RECT 201.995 1741.590 202.165 1741.760 ;
        RECT 201.995 1741.130 202.165 1741.300 ;
        RECT 201.995 1740.670 202.165 1740.840 ;
        RECT 201.995 1740.210 202.165 1740.380 ;
        RECT 201.995 1739.750 202.165 1739.920 ;
        RECT 201.995 1739.290 202.165 1739.460 ;
      LAYER li1 ;
        RECT 207.435 1739.235 208.150 1742.655 ;
        RECT 207.435 1739.145 207.605 1739.235 ;
      LAYER li1 ;
        RECT 201.995 1738.830 202.165 1739.000 ;
        RECT 207.435 1738.830 207.605 1739.000 ;
      LAYER li1 ;
        RECT 207.435 1738.600 207.605 1738.685 ;
        RECT 207.435 1738.540 208.150 1738.600 ;
      LAYER li1 ;
        RECT 201.995 1738.370 202.165 1738.540 ;
      LAYER li1 ;
        RECT 207.605 1738.370 208.150 1738.540 ;
      LAYER li1 ;
        RECT 201.995 1737.910 202.165 1738.080 ;
        RECT 201.995 1737.450 202.165 1737.620 ;
        RECT 201.995 1736.990 202.165 1737.160 ;
      LAYER li1 ;
        RECT 207.435 1737.015 208.150 1738.370 ;
      LAYER li1 ;
        RECT 201.995 1736.530 202.165 1736.700 ;
      LAYER li1 ;
        RECT 207.435 1736.675 208.980 1737.015 ;
      LAYER li1 ;
        RECT 201.995 1736.070 202.165 1736.240 ;
        RECT 201.995 1735.610 202.165 1735.780 ;
        RECT 201.995 1735.150 202.165 1735.320 ;
        RECT 201.995 1734.690 202.165 1734.860 ;
        RECT 201.995 1734.230 202.165 1734.400 ;
        RECT 201.995 1733.770 202.165 1733.940 ;
        RECT 201.995 1733.310 202.165 1733.480 ;
      LAYER li1 ;
        RECT 207.435 1733.255 208.150 1736.675 ;
        RECT 207.435 1733.165 207.605 1733.255 ;
      LAYER li1 ;
        RECT 201.995 1732.850 202.165 1733.020 ;
        RECT 207.435 1732.850 207.605 1733.020 ;
      LAYER li1 ;
        RECT 207.435 1732.620 207.605 1732.705 ;
        RECT 207.435 1732.560 208.150 1732.620 ;
      LAYER li1 ;
        RECT 201.995 1732.390 202.165 1732.560 ;
      LAYER li1 ;
        RECT 207.605 1732.390 208.150 1732.560 ;
      LAYER li1 ;
        RECT 201.995 1731.930 202.165 1732.100 ;
        RECT 201.995 1731.470 202.165 1731.640 ;
        RECT 201.995 1731.010 202.165 1731.180 ;
      LAYER li1 ;
        RECT 207.435 1731.035 208.150 1732.390 ;
      LAYER li1 ;
        RECT 201.995 1730.550 202.165 1730.720 ;
      LAYER li1 ;
        RECT 207.435 1730.695 208.980 1731.035 ;
      LAYER li1 ;
        RECT 201.995 1730.090 202.165 1730.260 ;
        RECT 201.995 1729.630 202.165 1729.800 ;
        RECT 201.995 1729.170 202.165 1729.340 ;
        RECT 201.995 1728.710 202.165 1728.880 ;
        RECT 201.995 1728.250 202.165 1728.420 ;
        RECT 201.995 1727.790 202.165 1727.960 ;
        RECT 201.995 1727.330 202.165 1727.500 ;
      LAYER li1 ;
        RECT 207.435 1727.275 208.150 1730.695 ;
        RECT 207.435 1727.185 207.605 1727.275 ;
      LAYER li1 ;
        RECT 201.995 1726.870 202.165 1727.040 ;
        RECT 207.435 1726.870 207.605 1727.040 ;
      LAYER li1 ;
        RECT 207.435 1726.640 207.605 1726.725 ;
        RECT 207.435 1726.580 208.150 1726.640 ;
      LAYER li1 ;
        RECT 201.995 1726.410 202.165 1726.580 ;
      LAYER li1 ;
        RECT 207.605 1726.410 208.150 1726.580 ;
      LAYER li1 ;
        RECT 201.995 1725.950 202.165 1726.120 ;
        RECT 201.995 1725.490 202.165 1725.660 ;
        RECT 201.995 1725.030 202.165 1725.200 ;
      LAYER li1 ;
        RECT 207.435 1725.055 208.150 1726.410 ;
      LAYER li1 ;
        RECT 201.995 1724.570 202.165 1724.740 ;
      LAYER li1 ;
        RECT 207.435 1724.715 208.980 1725.055 ;
      LAYER li1 ;
        RECT 201.995 1724.110 202.165 1724.280 ;
        RECT 201.995 1723.650 202.165 1723.820 ;
        RECT 201.995 1723.190 202.165 1723.360 ;
        RECT 201.995 1722.730 202.165 1722.900 ;
        RECT 201.995 1722.270 202.165 1722.440 ;
        RECT 201.995 1721.810 202.165 1721.980 ;
        RECT 201.995 1721.350 202.165 1721.520 ;
      LAYER li1 ;
        RECT 207.435 1721.295 208.150 1724.715 ;
        RECT 207.435 1721.205 207.605 1721.295 ;
      LAYER li1 ;
        RECT 201.995 1720.890 202.165 1721.060 ;
        RECT 207.435 1720.890 207.605 1721.060 ;
      LAYER li1 ;
        RECT 207.435 1720.660 207.605 1720.745 ;
        RECT 207.435 1720.600 208.150 1720.660 ;
      LAYER li1 ;
        RECT 201.995 1720.430 202.165 1720.600 ;
      LAYER li1 ;
        RECT 207.605 1720.430 208.150 1720.600 ;
      LAYER li1 ;
        RECT 201.995 1719.970 202.165 1720.140 ;
        RECT 201.995 1719.510 202.165 1719.680 ;
        RECT 201.995 1719.050 202.165 1719.220 ;
      LAYER li1 ;
        RECT 207.435 1719.075 208.150 1720.430 ;
      LAYER li1 ;
        RECT 201.995 1718.590 202.165 1718.760 ;
      LAYER li1 ;
        RECT 207.435 1718.735 208.980 1719.075 ;
      LAYER li1 ;
        RECT 201.995 1718.130 202.165 1718.300 ;
        RECT 201.995 1717.670 202.165 1717.840 ;
        RECT 201.995 1717.210 202.165 1717.380 ;
        RECT 201.995 1716.750 202.165 1716.920 ;
        RECT 201.995 1716.290 202.165 1716.460 ;
        RECT 201.995 1715.830 202.165 1716.000 ;
        RECT 201.995 1715.370 202.165 1715.540 ;
      LAYER li1 ;
        RECT 207.435 1715.315 208.150 1718.735 ;
        RECT 207.435 1715.225 207.605 1715.315 ;
      LAYER li1 ;
        RECT 201.995 1714.910 202.165 1715.080 ;
        RECT 207.435 1714.910 207.605 1715.080 ;
      LAYER li1 ;
        RECT 207.435 1714.680 207.605 1714.765 ;
        RECT 207.435 1714.620 208.150 1714.680 ;
      LAYER li1 ;
        RECT 201.995 1714.450 202.165 1714.620 ;
      LAYER li1 ;
        RECT 207.605 1714.450 208.150 1714.620 ;
      LAYER li1 ;
        RECT 201.995 1713.990 202.165 1714.160 ;
        RECT 201.995 1713.530 202.165 1713.700 ;
        RECT 201.995 1713.070 202.165 1713.240 ;
      LAYER li1 ;
        RECT 207.435 1713.095 208.150 1714.450 ;
      LAYER li1 ;
        RECT 201.995 1712.610 202.165 1712.780 ;
      LAYER li1 ;
        RECT 207.435 1712.755 208.980 1713.095 ;
      LAYER li1 ;
        RECT 201.995 1712.150 202.165 1712.320 ;
        RECT 201.995 1711.690 202.165 1711.860 ;
        RECT 201.995 1711.230 202.165 1711.400 ;
        RECT 201.995 1710.770 202.165 1710.940 ;
        RECT 201.995 1710.310 202.165 1710.480 ;
        RECT 201.995 1709.850 202.165 1710.020 ;
        RECT 201.995 1709.390 202.165 1709.560 ;
      LAYER li1 ;
        RECT 207.435 1709.335 208.150 1712.755 ;
        RECT 207.435 1709.245 207.605 1709.335 ;
      LAYER li1 ;
        RECT 201.995 1708.930 202.165 1709.100 ;
        RECT 207.435 1708.930 207.605 1709.100 ;
      LAYER li1 ;
        RECT 207.435 1708.700 207.605 1708.785 ;
        RECT 207.435 1708.640 208.150 1708.700 ;
      LAYER li1 ;
        RECT 201.995 1708.470 202.165 1708.640 ;
      LAYER li1 ;
        RECT 207.605 1708.470 208.150 1708.640 ;
      LAYER li1 ;
        RECT 201.995 1708.010 202.165 1708.180 ;
        RECT 201.995 1707.550 202.165 1707.720 ;
        RECT 201.995 1707.090 202.165 1707.260 ;
      LAYER li1 ;
        RECT 207.435 1707.115 208.150 1708.470 ;
      LAYER li1 ;
        RECT 201.995 1706.630 202.165 1706.800 ;
      LAYER li1 ;
        RECT 207.435 1706.775 208.980 1707.115 ;
      LAYER li1 ;
        RECT 201.995 1706.170 202.165 1706.340 ;
        RECT 201.995 1705.710 202.165 1705.880 ;
        RECT 201.995 1705.250 202.165 1705.420 ;
        RECT 201.995 1704.790 202.165 1704.960 ;
        RECT 201.995 1704.330 202.165 1704.500 ;
        RECT 201.995 1703.870 202.165 1704.040 ;
        RECT 201.995 1703.410 202.165 1703.580 ;
      LAYER li1 ;
        RECT 207.435 1703.355 208.150 1706.775 ;
        RECT 207.435 1703.265 207.605 1703.355 ;
      LAYER li1 ;
        RECT 201.995 1702.950 202.165 1703.120 ;
        RECT 207.435 1702.950 207.605 1703.120 ;
      LAYER li1 ;
        RECT 207.435 1702.720 207.605 1702.805 ;
        RECT 207.435 1702.660 208.150 1702.720 ;
      LAYER li1 ;
        RECT 201.995 1702.490 202.165 1702.660 ;
      LAYER li1 ;
        RECT 207.605 1702.490 208.150 1702.660 ;
      LAYER li1 ;
        RECT 201.995 1702.030 202.165 1702.200 ;
        RECT 201.995 1701.570 202.165 1701.740 ;
        RECT 201.995 1701.110 202.165 1701.280 ;
      LAYER li1 ;
        RECT 207.435 1701.135 208.150 1702.490 ;
      LAYER li1 ;
        RECT 201.995 1700.650 202.165 1700.820 ;
      LAYER li1 ;
        RECT 207.435 1700.795 208.980 1701.135 ;
      LAYER li1 ;
        RECT 201.995 1700.190 202.165 1700.360 ;
        RECT 201.995 1699.730 202.165 1699.900 ;
        RECT 201.995 1699.270 202.165 1699.440 ;
        RECT 201.995 1698.810 202.165 1698.980 ;
        RECT 201.995 1698.350 202.165 1698.520 ;
        RECT 201.995 1697.890 202.165 1698.060 ;
        RECT 201.995 1697.430 202.165 1697.600 ;
      LAYER li1 ;
        RECT 207.435 1697.375 208.150 1700.795 ;
        RECT 207.435 1697.285 207.605 1697.375 ;
      LAYER li1 ;
        RECT 201.995 1696.970 202.165 1697.140 ;
        RECT 207.435 1696.970 207.605 1697.140 ;
      LAYER li1 ;
        RECT 207.435 1696.740 207.605 1696.825 ;
        RECT 207.435 1696.680 208.150 1696.740 ;
      LAYER li1 ;
        RECT 201.995 1696.510 202.165 1696.680 ;
      LAYER li1 ;
        RECT 207.605 1696.510 208.150 1696.680 ;
      LAYER li1 ;
        RECT 201.995 1696.050 202.165 1696.220 ;
        RECT 201.995 1695.590 202.165 1695.760 ;
        RECT 201.995 1695.130 202.165 1695.300 ;
      LAYER li1 ;
        RECT 207.435 1695.155 208.150 1696.510 ;
      LAYER li1 ;
        RECT 201.995 1694.670 202.165 1694.840 ;
      LAYER li1 ;
        RECT 207.435 1694.815 208.980 1695.155 ;
      LAYER li1 ;
        RECT 201.995 1694.210 202.165 1694.380 ;
        RECT 201.995 1693.750 202.165 1693.920 ;
        RECT 201.995 1693.290 202.165 1693.460 ;
        RECT 201.995 1692.830 202.165 1693.000 ;
        RECT 201.995 1692.370 202.165 1692.540 ;
        RECT 201.995 1691.910 202.165 1692.080 ;
        RECT 201.995 1691.450 202.165 1691.620 ;
      LAYER li1 ;
        RECT 207.435 1691.395 208.150 1694.815 ;
        RECT 207.435 1691.305 207.605 1691.395 ;
      LAYER li1 ;
        RECT 201.995 1690.990 202.165 1691.160 ;
        RECT 207.435 1690.990 207.605 1691.160 ;
      LAYER li1 ;
        RECT 207.435 1690.760 207.605 1690.845 ;
        RECT 207.435 1690.700 208.150 1690.760 ;
      LAYER li1 ;
        RECT 201.995 1690.530 202.165 1690.700 ;
      LAYER li1 ;
        RECT 207.605 1690.530 208.150 1690.700 ;
      LAYER li1 ;
        RECT 201.995 1690.070 202.165 1690.240 ;
        RECT 201.995 1689.610 202.165 1689.780 ;
        RECT 201.995 1689.150 202.165 1689.320 ;
      LAYER li1 ;
        RECT 207.435 1689.175 208.150 1690.530 ;
      LAYER li1 ;
        RECT 201.995 1688.690 202.165 1688.860 ;
      LAYER li1 ;
        RECT 207.435 1688.835 208.980 1689.175 ;
      LAYER li1 ;
        RECT 201.995 1688.230 202.165 1688.400 ;
        RECT 201.995 1687.770 202.165 1687.940 ;
        RECT 201.995 1687.310 202.165 1687.480 ;
        RECT 201.995 1686.850 202.165 1687.020 ;
        RECT 201.995 1686.390 202.165 1686.560 ;
        RECT 201.995 1685.930 202.165 1686.100 ;
        RECT 201.995 1685.470 202.165 1685.640 ;
      LAYER li1 ;
        RECT 207.435 1685.415 208.150 1688.835 ;
        RECT 207.435 1685.325 207.605 1685.415 ;
      LAYER li1 ;
        RECT 201.995 1685.010 202.165 1685.180 ;
        RECT 207.435 1685.010 207.605 1685.180 ;
      LAYER li1 ;
        RECT 207.435 1684.780 207.605 1684.865 ;
        RECT 207.435 1684.720 208.150 1684.780 ;
      LAYER li1 ;
        RECT 201.995 1684.550 202.165 1684.720 ;
      LAYER li1 ;
        RECT 207.605 1684.550 208.150 1684.720 ;
      LAYER li1 ;
        RECT 201.995 1684.090 202.165 1684.260 ;
        RECT 201.995 1683.630 202.165 1683.800 ;
        RECT 201.995 1683.170 202.165 1683.340 ;
      LAYER li1 ;
        RECT 207.435 1683.195 208.150 1684.550 ;
      LAYER li1 ;
        RECT 201.995 1682.710 202.165 1682.880 ;
      LAYER li1 ;
        RECT 207.435 1682.855 208.980 1683.195 ;
      LAYER li1 ;
        RECT 201.995 1682.250 202.165 1682.420 ;
        RECT 201.995 1681.790 202.165 1681.960 ;
        RECT 201.995 1681.330 202.165 1681.500 ;
        RECT 201.995 1680.870 202.165 1681.040 ;
        RECT 201.995 1680.410 202.165 1680.580 ;
        RECT 201.995 1679.950 202.165 1680.120 ;
        RECT 201.995 1679.490 202.165 1679.660 ;
      LAYER li1 ;
        RECT 207.435 1679.435 208.150 1682.855 ;
        RECT 207.435 1679.345 207.605 1679.435 ;
      LAYER li1 ;
        RECT 201.995 1679.030 202.165 1679.200 ;
        RECT 207.435 1679.030 207.605 1679.200 ;
      LAYER li1 ;
        RECT 207.435 1678.800 207.605 1678.885 ;
        RECT 207.435 1678.740 208.150 1678.800 ;
      LAYER li1 ;
        RECT 201.995 1678.570 202.165 1678.740 ;
      LAYER li1 ;
        RECT 207.605 1678.570 208.150 1678.740 ;
      LAYER li1 ;
        RECT 201.995 1678.110 202.165 1678.280 ;
        RECT 201.995 1677.650 202.165 1677.820 ;
        RECT 201.995 1677.190 202.165 1677.360 ;
      LAYER li1 ;
        RECT 207.435 1677.215 208.150 1678.570 ;
      LAYER li1 ;
        RECT 201.995 1676.730 202.165 1676.900 ;
      LAYER li1 ;
        RECT 207.435 1676.875 208.980 1677.215 ;
      LAYER li1 ;
        RECT 201.995 1676.270 202.165 1676.440 ;
        RECT 201.995 1675.810 202.165 1675.980 ;
        RECT 201.995 1675.350 202.165 1675.520 ;
        RECT 201.995 1674.890 202.165 1675.060 ;
        RECT 201.995 1674.430 202.165 1674.600 ;
        RECT 201.995 1673.970 202.165 1674.140 ;
        RECT 201.995 1673.510 202.165 1673.680 ;
      LAYER li1 ;
        RECT 207.435 1673.455 208.150 1676.875 ;
        RECT 207.435 1673.365 207.605 1673.455 ;
      LAYER li1 ;
        RECT 201.995 1673.050 202.165 1673.220 ;
        RECT 207.435 1673.050 207.605 1673.220 ;
      LAYER mcon ;
        RECT 207.435 1761.830 207.605 1762.000 ;
        RECT 207.435 1761.370 207.605 1761.540 ;
        RECT 207.435 1760.910 207.605 1761.080 ;
        RECT 207.435 1760.450 207.605 1760.620 ;
        RECT 207.435 1759.990 207.605 1760.160 ;
        RECT 207.435 1759.530 207.605 1759.700 ;
        RECT 207.435 1759.070 207.605 1759.240 ;
        RECT 207.435 1758.610 207.605 1758.780 ;
        RECT 207.435 1758.150 207.605 1758.320 ;
        RECT 207.435 1757.690 207.605 1757.860 ;
        RECT 207.435 1757.230 207.605 1757.400 ;
        RECT 207.435 1755.850 207.605 1756.020 ;
        RECT 207.435 1755.390 207.605 1755.560 ;
        RECT 207.435 1754.930 207.605 1755.100 ;
        RECT 207.435 1754.470 207.605 1754.640 ;
        RECT 207.435 1754.010 207.605 1754.180 ;
        RECT 207.435 1753.550 207.605 1753.720 ;
        RECT 207.435 1753.090 207.605 1753.260 ;
        RECT 207.435 1752.630 207.605 1752.800 ;
        RECT 207.435 1752.170 207.605 1752.340 ;
        RECT 207.435 1751.710 207.605 1751.880 ;
        RECT 207.435 1751.250 207.605 1751.420 ;
        RECT 207.435 1743.890 207.605 1744.060 ;
        RECT 207.435 1743.430 207.605 1743.600 ;
        RECT 207.435 1742.970 207.605 1743.140 ;
        RECT 207.435 1742.510 207.605 1742.680 ;
        RECT 207.435 1742.050 207.605 1742.220 ;
        RECT 207.435 1741.590 207.605 1741.760 ;
        RECT 207.435 1741.130 207.605 1741.300 ;
        RECT 207.435 1740.670 207.605 1740.840 ;
        RECT 207.435 1740.210 207.605 1740.380 ;
        RECT 207.435 1739.750 207.605 1739.920 ;
        RECT 207.435 1739.290 207.605 1739.460 ;
        RECT 207.435 1737.910 207.605 1738.080 ;
        RECT 207.435 1737.450 207.605 1737.620 ;
        RECT 207.435 1736.990 207.605 1737.160 ;
        RECT 207.435 1736.530 207.605 1736.700 ;
        RECT 207.435 1736.070 207.605 1736.240 ;
        RECT 207.435 1735.610 207.605 1735.780 ;
        RECT 207.435 1735.150 207.605 1735.320 ;
        RECT 207.435 1734.690 207.605 1734.860 ;
        RECT 207.435 1734.230 207.605 1734.400 ;
        RECT 207.435 1733.770 207.605 1733.940 ;
        RECT 207.435 1733.310 207.605 1733.480 ;
        RECT 207.435 1731.930 207.605 1732.100 ;
        RECT 207.435 1731.470 207.605 1731.640 ;
        RECT 207.435 1731.010 207.605 1731.180 ;
        RECT 207.435 1730.550 207.605 1730.720 ;
        RECT 207.435 1730.090 207.605 1730.260 ;
        RECT 207.435 1729.630 207.605 1729.800 ;
        RECT 207.435 1729.170 207.605 1729.340 ;
        RECT 207.435 1728.710 207.605 1728.880 ;
        RECT 207.435 1728.250 207.605 1728.420 ;
        RECT 207.435 1727.790 207.605 1727.960 ;
        RECT 207.435 1727.330 207.605 1727.500 ;
        RECT 207.435 1725.950 207.605 1726.120 ;
        RECT 207.435 1725.490 207.605 1725.660 ;
        RECT 207.435 1725.030 207.605 1725.200 ;
        RECT 207.435 1724.570 207.605 1724.740 ;
        RECT 207.435 1724.110 207.605 1724.280 ;
        RECT 207.435 1723.650 207.605 1723.820 ;
        RECT 207.435 1723.190 207.605 1723.360 ;
        RECT 207.435 1722.730 207.605 1722.900 ;
        RECT 207.435 1722.270 207.605 1722.440 ;
        RECT 207.435 1721.810 207.605 1721.980 ;
        RECT 207.435 1721.350 207.605 1721.520 ;
        RECT 207.435 1719.970 207.605 1720.140 ;
        RECT 207.435 1719.510 207.605 1719.680 ;
        RECT 207.435 1719.050 207.605 1719.220 ;
        RECT 207.435 1718.590 207.605 1718.760 ;
        RECT 207.435 1718.130 207.605 1718.300 ;
        RECT 207.435 1717.670 207.605 1717.840 ;
        RECT 207.435 1717.210 207.605 1717.380 ;
        RECT 207.435 1716.750 207.605 1716.920 ;
        RECT 207.435 1716.290 207.605 1716.460 ;
        RECT 207.435 1715.830 207.605 1716.000 ;
        RECT 207.435 1715.370 207.605 1715.540 ;
        RECT 207.435 1713.990 207.605 1714.160 ;
        RECT 207.435 1713.530 207.605 1713.700 ;
        RECT 207.435 1713.070 207.605 1713.240 ;
        RECT 207.435 1712.610 207.605 1712.780 ;
        RECT 207.435 1712.150 207.605 1712.320 ;
        RECT 207.435 1711.690 207.605 1711.860 ;
        RECT 207.435 1711.230 207.605 1711.400 ;
        RECT 207.435 1710.770 207.605 1710.940 ;
        RECT 207.435 1710.310 207.605 1710.480 ;
        RECT 207.435 1709.850 207.605 1710.020 ;
        RECT 207.435 1709.390 207.605 1709.560 ;
        RECT 207.435 1708.010 207.605 1708.180 ;
        RECT 207.435 1707.550 207.605 1707.720 ;
        RECT 207.435 1707.090 207.605 1707.260 ;
        RECT 207.435 1706.630 207.605 1706.800 ;
        RECT 207.435 1706.170 207.605 1706.340 ;
        RECT 207.435 1705.710 207.605 1705.880 ;
        RECT 207.435 1705.250 207.605 1705.420 ;
        RECT 207.435 1704.790 207.605 1704.960 ;
        RECT 207.435 1704.330 207.605 1704.500 ;
        RECT 207.435 1703.870 207.605 1704.040 ;
        RECT 207.435 1703.410 207.605 1703.580 ;
        RECT 207.435 1702.030 207.605 1702.200 ;
        RECT 207.435 1701.570 207.605 1701.740 ;
        RECT 207.435 1701.110 207.605 1701.280 ;
        RECT 207.435 1700.650 207.605 1700.820 ;
        RECT 207.435 1700.190 207.605 1700.360 ;
        RECT 207.435 1699.730 207.605 1699.900 ;
        RECT 207.435 1699.270 207.605 1699.440 ;
        RECT 207.435 1698.810 207.605 1698.980 ;
        RECT 207.435 1698.350 207.605 1698.520 ;
        RECT 207.435 1697.890 207.605 1698.060 ;
        RECT 207.435 1697.430 207.605 1697.600 ;
        RECT 207.435 1696.050 207.605 1696.220 ;
        RECT 207.435 1695.590 207.605 1695.760 ;
        RECT 207.435 1695.130 207.605 1695.300 ;
        RECT 207.435 1694.670 207.605 1694.840 ;
        RECT 207.435 1694.210 207.605 1694.380 ;
        RECT 207.435 1693.750 207.605 1693.920 ;
        RECT 207.435 1693.290 207.605 1693.460 ;
        RECT 207.435 1692.830 207.605 1693.000 ;
        RECT 207.435 1692.370 207.605 1692.540 ;
        RECT 207.435 1691.910 207.605 1692.080 ;
        RECT 207.435 1691.450 207.605 1691.620 ;
        RECT 207.435 1690.070 207.605 1690.240 ;
        RECT 207.435 1689.610 207.605 1689.780 ;
        RECT 207.435 1689.150 207.605 1689.320 ;
        RECT 207.435 1688.690 207.605 1688.860 ;
        RECT 207.435 1688.230 207.605 1688.400 ;
        RECT 207.435 1687.770 207.605 1687.940 ;
        RECT 207.435 1687.310 207.605 1687.480 ;
        RECT 207.435 1686.850 207.605 1687.020 ;
        RECT 207.435 1686.390 207.605 1686.560 ;
        RECT 207.435 1685.930 207.605 1686.100 ;
        RECT 207.435 1685.470 207.605 1685.640 ;
        RECT 207.435 1684.090 207.605 1684.260 ;
        RECT 207.435 1683.630 207.605 1683.800 ;
        RECT 207.435 1683.170 207.605 1683.340 ;
        RECT 207.435 1682.710 207.605 1682.880 ;
        RECT 207.435 1682.250 207.605 1682.420 ;
        RECT 207.435 1681.790 207.605 1681.960 ;
        RECT 207.435 1681.330 207.605 1681.500 ;
        RECT 207.435 1680.870 207.605 1681.040 ;
        RECT 207.435 1680.410 207.605 1680.580 ;
        RECT 207.435 1679.950 207.605 1680.120 ;
        RECT 207.435 1679.490 207.605 1679.660 ;
        RECT 207.435 1678.110 207.605 1678.280 ;
        RECT 207.435 1677.650 207.605 1677.820 ;
        RECT 207.435 1677.190 207.605 1677.360 ;
        RECT 207.435 1676.730 207.605 1676.900 ;
        RECT 207.435 1676.270 207.605 1676.440 ;
        RECT 207.435 1675.810 207.605 1675.980 ;
        RECT 207.435 1675.350 207.605 1675.520 ;
        RECT 207.435 1674.890 207.605 1675.060 ;
        RECT 207.435 1674.430 207.605 1674.600 ;
        RECT 207.435 1673.970 207.605 1674.140 ;
        RECT 207.435 1673.510 207.605 1673.680 ;
      LAYER met1 ;
        RECT 201.840 1672.905 202.320 1763.065 ;
        RECT 207.280 1672.905 207.760 1763.065 ;
      LAYER via ;
        RECT 201.950 1734.795 202.250 1736.580 ;
        RECT 207.360 1734.795 207.660 1736.580 ;
      LAYER met2 ;
        RECT 201.865 1734.755 202.295 1736.620 ;
        RECT 207.290 1734.755 207.720 1736.620 ;
      LAYER via2 ;
        RECT 201.950 1734.795 202.250 1736.580 ;
        RECT 207.360 1734.795 207.660 1736.580 ;
      LAYER met3 ;
        RECT 200.210 1734.750 207.735 1736.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.885 3050.655 202.055 3050.825 ;
        RECT 207.325 3050.655 207.495 3050.825 ;
        RECT 201.885 3050.195 202.055 3050.365 ;
        RECT 207.325 3050.195 207.495 3050.365 ;
        RECT 201.885 3049.735 202.055 3049.905 ;
        RECT 207.325 3049.735 207.495 3049.905 ;
        RECT 201.885 3049.275 202.055 3049.445 ;
        RECT 207.325 3049.275 207.495 3049.445 ;
        RECT 201.885 3048.815 202.055 3048.985 ;
        RECT 207.325 3048.815 207.495 3048.985 ;
        RECT 201.885 3048.355 202.055 3048.525 ;
        RECT 207.325 3048.355 207.495 3048.525 ;
        RECT 201.885 3047.895 202.055 3048.065 ;
        RECT 207.325 3047.895 207.495 3048.065 ;
        RECT 201.885 3047.435 202.055 3047.605 ;
        RECT 207.325 3047.435 207.495 3047.605 ;
        RECT 201.885 3046.975 202.055 3047.145 ;
        RECT 207.325 3046.975 207.495 3047.145 ;
        RECT 201.885 3046.515 202.055 3046.685 ;
        RECT 207.325 3046.515 207.495 3046.685 ;
        RECT 201.885 3046.055 202.055 3046.225 ;
        RECT 207.325 3046.055 207.495 3046.225 ;
        RECT 201.885 3045.595 202.055 3045.765 ;
        RECT 207.325 3045.595 207.495 3045.765 ;
        RECT 201.885 3045.135 202.055 3045.305 ;
        RECT 207.325 3045.135 207.495 3045.305 ;
        RECT 201.885 3044.675 202.055 3044.845 ;
        RECT 207.325 3044.675 207.495 3044.845 ;
        RECT 201.885 3044.215 202.055 3044.385 ;
        RECT 207.325 3044.215 207.495 3044.385 ;
        RECT 201.885 3043.755 202.055 3043.925 ;
        RECT 207.325 3043.755 207.495 3043.925 ;
        RECT 201.885 3043.295 202.055 3043.465 ;
        RECT 207.325 3043.295 207.495 3043.465 ;
        RECT 201.885 3042.835 202.055 3043.005 ;
        RECT 207.325 3042.835 207.495 3043.005 ;
        RECT 201.885 3042.375 202.055 3042.545 ;
        RECT 207.325 3042.375 207.495 3042.545 ;
        RECT 201.885 3041.915 202.055 3042.085 ;
        RECT 207.325 3041.915 207.495 3042.085 ;
        RECT 201.885 3041.455 202.055 3041.625 ;
        RECT 207.325 3041.455 207.495 3041.625 ;
        RECT 201.885 3040.995 202.055 3041.165 ;
        RECT 207.325 3040.995 207.495 3041.165 ;
        RECT 201.885 3040.535 202.055 3040.705 ;
        RECT 207.325 3040.535 207.495 3040.705 ;
        RECT 201.885 3040.075 202.055 3040.245 ;
        RECT 207.325 3040.075 207.495 3040.245 ;
        RECT 201.885 3039.615 202.055 3039.785 ;
        RECT 207.325 3039.615 207.495 3039.785 ;
        RECT 201.885 3039.155 202.055 3039.325 ;
        RECT 207.325 3039.155 207.495 3039.325 ;
        RECT 201.885 3038.695 202.055 3038.865 ;
        RECT 207.325 3038.695 207.495 3038.865 ;
        RECT 201.885 3038.235 202.055 3038.405 ;
        RECT 207.325 3038.235 207.495 3038.405 ;
        RECT 201.885 3037.775 202.055 3037.945 ;
        RECT 207.325 3037.775 207.495 3037.945 ;
        RECT 201.885 3037.315 202.055 3037.485 ;
        RECT 207.325 3037.315 207.495 3037.485 ;
        RECT 201.885 3036.855 202.055 3037.025 ;
        RECT 207.325 3036.855 207.495 3037.025 ;
        RECT 201.885 3036.395 202.055 3036.565 ;
        RECT 207.325 3036.395 207.495 3036.565 ;
        RECT 201.885 3035.935 202.055 3036.105 ;
        RECT 207.325 3035.935 207.495 3036.105 ;
        RECT 201.885 3035.475 202.055 3035.645 ;
        RECT 207.325 3035.475 207.495 3035.645 ;
        RECT 201.885 3035.015 202.055 3035.185 ;
        RECT 207.325 3035.015 207.495 3035.185 ;
        RECT 201.885 3034.555 202.055 3034.725 ;
        RECT 207.325 3034.555 207.495 3034.725 ;
        RECT 201.885 3034.095 202.055 3034.265 ;
        RECT 207.325 3034.095 207.495 3034.265 ;
        RECT 201.885 3033.635 202.055 3033.805 ;
        RECT 207.325 3033.635 207.495 3033.805 ;
        RECT 201.885 3033.175 202.055 3033.345 ;
        RECT 207.325 3033.175 207.495 3033.345 ;
        RECT 201.885 3032.715 202.055 3032.885 ;
        RECT 207.325 3032.715 207.495 3032.885 ;
        RECT 201.885 3032.255 202.055 3032.425 ;
        RECT 207.325 3032.255 207.495 3032.425 ;
        RECT 201.885 3031.795 202.055 3031.965 ;
        RECT 207.325 3031.795 207.495 3031.965 ;
        RECT 201.885 3031.335 202.055 3031.505 ;
        RECT 207.325 3031.335 207.495 3031.505 ;
        RECT 201.885 3030.875 202.055 3031.045 ;
        RECT 207.325 3030.875 207.495 3031.045 ;
        RECT 201.885 3030.415 202.055 3030.585 ;
        RECT 207.325 3030.415 207.495 3030.585 ;
        RECT 201.885 3029.955 202.055 3030.125 ;
        RECT 207.325 3029.955 207.495 3030.125 ;
        RECT 201.885 3029.495 202.055 3029.665 ;
        RECT 207.325 3029.495 207.495 3029.665 ;
        RECT 201.885 3029.035 202.055 3029.205 ;
        RECT 207.325 3029.035 207.495 3029.205 ;
        RECT 201.885 3028.575 202.055 3028.745 ;
        RECT 207.325 3028.575 207.495 3028.745 ;
        RECT 201.885 3028.115 202.055 3028.285 ;
        RECT 207.325 3028.115 207.495 3028.285 ;
        RECT 201.885 3027.655 202.055 3027.825 ;
        RECT 207.325 3027.655 207.495 3027.825 ;
        RECT 201.885 3027.195 202.055 3027.365 ;
        RECT 207.325 3027.195 207.495 3027.365 ;
        RECT 201.885 3026.735 202.055 3026.905 ;
        RECT 207.325 3026.735 207.495 3026.905 ;
        RECT 201.885 3026.275 202.055 3026.445 ;
        RECT 207.325 3026.275 207.495 3026.445 ;
        RECT 201.885 3025.815 202.055 3025.985 ;
        RECT 207.325 3025.815 207.495 3025.985 ;
        RECT 201.885 3025.355 202.055 3025.525 ;
        RECT 207.325 3025.355 207.495 3025.525 ;
        RECT 201.885 3024.895 202.055 3025.065 ;
        RECT 207.325 3024.895 207.495 3025.065 ;
        RECT 201.885 3024.435 202.055 3024.605 ;
        RECT 207.325 3024.435 207.495 3024.605 ;
        RECT 201.885 3023.975 202.055 3024.145 ;
        RECT 207.325 3023.975 207.495 3024.145 ;
        RECT 201.885 3023.515 202.055 3023.685 ;
        RECT 207.325 3023.515 207.495 3023.685 ;
        RECT 201.885 3023.055 202.055 3023.225 ;
        RECT 207.325 3023.055 207.495 3023.225 ;
        RECT 201.885 3022.595 202.055 3022.765 ;
        RECT 207.325 3022.595 207.495 3022.765 ;
        RECT 201.885 3022.135 202.055 3022.305 ;
        RECT 207.325 3022.135 207.495 3022.305 ;
        RECT 201.885 3021.675 202.055 3021.845 ;
        RECT 207.325 3021.675 207.495 3021.845 ;
        RECT 201.885 3021.215 202.055 3021.385 ;
        RECT 207.325 3021.215 207.495 3021.385 ;
        RECT 201.885 3020.755 202.055 3020.925 ;
        RECT 207.325 3020.755 207.495 3020.925 ;
        RECT 201.885 3020.295 202.055 3020.465 ;
        RECT 207.325 3020.295 207.495 3020.465 ;
        RECT 201.885 3019.835 202.055 3020.005 ;
        RECT 207.325 3019.835 207.495 3020.005 ;
        RECT 201.885 3019.375 202.055 3019.545 ;
        RECT 207.325 3019.375 207.495 3019.545 ;
        RECT 201.885 3018.915 202.055 3019.085 ;
        RECT 207.325 3018.915 207.495 3019.085 ;
        RECT 201.885 3018.455 202.055 3018.625 ;
        RECT 207.325 3018.455 207.495 3018.625 ;
        RECT 201.885 3017.995 202.055 3018.165 ;
        RECT 207.325 3017.995 207.495 3018.165 ;
        RECT 201.885 3017.535 202.055 3017.705 ;
        RECT 207.325 3017.535 207.495 3017.705 ;
        RECT 201.885 3017.075 202.055 3017.245 ;
        RECT 207.325 3017.075 207.495 3017.245 ;
        RECT 201.885 3016.615 202.055 3016.785 ;
        RECT 207.325 3016.615 207.495 3016.785 ;
        RECT 201.885 3016.155 202.055 3016.325 ;
        RECT 207.325 3016.155 207.495 3016.325 ;
        RECT 201.885 3015.695 202.055 3015.865 ;
        RECT 207.325 3015.695 207.495 3015.865 ;
        RECT 201.885 3015.235 202.055 3015.405 ;
        RECT 207.325 3015.235 207.495 3015.405 ;
        RECT 201.885 3014.775 202.055 3014.945 ;
        RECT 207.325 3014.775 207.495 3014.945 ;
        RECT 201.885 3014.315 202.055 3014.485 ;
        RECT 207.325 3014.315 207.495 3014.485 ;
        RECT 201.885 3013.855 202.055 3014.025 ;
        RECT 207.325 3013.855 207.495 3014.025 ;
        RECT 201.885 3013.395 202.055 3013.565 ;
        RECT 207.325 3013.395 207.495 3013.565 ;
        RECT 201.885 3012.935 202.055 3013.105 ;
        RECT 207.325 3012.935 207.495 3013.105 ;
        RECT 201.885 3012.475 202.055 3012.645 ;
        RECT 207.325 3012.475 207.495 3012.645 ;
        RECT 201.885 3012.015 202.055 3012.185 ;
        RECT 207.325 3012.015 207.495 3012.185 ;
        RECT 201.885 3011.555 202.055 3011.725 ;
        RECT 207.325 3011.555 207.495 3011.725 ;
        RECT 201.885 3011.095 202.055 3011.265 ;
        RECT 207.325 3011.095 207.495 3011.265 ;
        RECT 201.885 3010.635 202.055 3010.805 ;
        RECT 207.325 3010.635 207.495 3010.805 ;
        RECT 201.885 3010.175 202.055 3010.345 ;
        RECT 207.325 3010.175 207.495 3010.345 ;
        RECT 201.885 3009.715 202.055 3009.885 ;
        RECT 207.325 3009.715 207.495 3009.885 ;
        RECT 201.885 3009.255 202.055 3009.425 ;
        RECT 207.325 3009.255 207.495 3009.425 ;
        RECT 201.885 3008.795 202.055 3008.965 ;
        RECT 207.325 3008.795 207.495 3008.965 ;
        RECT 201.885 3008.335 202.055 3008.505 ;
        RECT 207.325 3008.335 207.495 3008.505 ;
        RECT 201.885 3007.875 202.055 3008.045 ;
        RECT 207.325 3007.875 207.495 3008.045 ;
        RECT 201.885 3007.415 202.055 3007.585 ;
        RECT 207.325 3007.415 207.495 3007.585 ;
        RECT 201.885 3006.955 202.055 3007.125 ;
        RECT 207.325 3006.955 207.495 3007.125 ;
        RECT 201.885 3006.495 202.055 3006.665 ;
        RECT 207.325 3006.495 207.495 3006.665 ;
        RECT 201.885 3006.035 202.055 3006.205 ;
        RECT 207.325 3006.035 207.495 3006.205 ;
        RECT 201.885 3005.575 202.055 3005.745 ;
        RECT 207.325 3005.575 207.495 3005.745 ;
        RECT 201.885 3005.115 202.055 3005.285 ;
        RECT 207.325 3005.115 207.495 3005.285 ;
        RECT 201.885 3004.655 202.055 3004.825 ;
        RECT 207.325 3004.655 207.495 3004.825 ;
        RECT 201.885 3004.195 202.055 3004.365 ;
        RECT 207.325 3004.195 207.495 3004.365 ;
        RECT 201.885 3003.735 202.055 3003.905 ;
        RECT 207.325 3003.735 207.495 3003.905 ;
        RECT 201.885 3003.275 202.055 3003.445 ;
        RECT 207.325 3003.275 207.495 3003.445 ;
        RECT 201.885 3002.815 202.055 3002.985 ;
        RECT 207.325 3002.815 207.495 3002.985 ;
        RECT 201.885 3002.355 202.055 3002.525 ;
        RECT 207.325 3002.355 207.495 3002.525 ;
        RECT 201.885 3001.895 202.055 3002.065 ;
        RECT 207.325 3001.895 207.495 3002.065 ;
        RECT 201.885 3001.435 202.055 3001.605 ;
        RECT 207.325 3001.435 207.495 3001.605 ;
        RECT 201.885 3000.975 202.055 3001.145 ;
        RECT 207.325 3000.975 207.495 3001.145 ;
        RECT 201.885 3000.515 202.055 3000.685 ;
        RECT 207.325 3000.515 207.495 3000.685 ;
        RECT 201.885 3000.055 202.055 3000.225 ;
        RECT 207.325 3000.055 207.495 3000.225 ;
        RECT 201.885 2999.595 202.055 2999.765 ;
        RECT 207.325 2999.595 207.495 2999.765 ;
        RECT 201.885 2999.135 202.055 2999.305 ;
        RECT 207.325 2999.135 207.495 2999.305 ;
        RECT 201.885 2998.675 202.055 2998.845 ;
        RECT 207.325 2998.675 207.495 2998.845 ;
        RECT 201.885 2998.215 202.055 2998.385 ;
        RECT 207.325 2998.215 207.495 2998.385 ;
        RECT 201.885 2997.755 202.055 2997.925 ;
        RECT 207.325 2997.755 207.495 2997.925 ;
        RECT 201.885 2997.295 202.055 2997.465 ;
        RECT 207.325 2997.295 207.495 2997.465 ;
        RECT 201.885 2996.835 202.055 2997.005 ;
        RECT 207.325 2996.835 207.495 2997.005 ;
        RECT 201.885 2996.375 202.055 2996.545 ;
        RECT 207.325 2996.375 207.495 2996.545 ;
        RECT 201.885 2995.915 202.055 2996.085 ;
        RECT 207.325 2995.915 207.495 2996.085 ;
        RECT 201.885 2995.455 202.055 2995.625 ;
        RECT 207.325 2995.455 207.495 2995.625 ;
        RECT 201.885 2994.995 202.055 2995.165 ;
        RECT 207.325 2994.995 207.495 2995.165 ;
        RECT 201.885 2994.535 202.055 2994.705 ;
        RECT 207.325 2994.535 207.495 2994.705 ;
        RECT 201.885 2994.075 202.055 2994.245 ;
        RECT 207.325 2994.075 207.495 2994.245 ;
        RECT 201.885 2993.615 202.055 2993.785 ;
        RECT 207.325 2993.615 207.495 2993.785 ;
        RECT 201.885 2993.155 202.055 2993.325 ;
        RECT 207.325 2993.155 207.495 2993.325 ;
        RECT 201.885 2992.695 202.055 2992.865 ;
        RECT 207.325 2992.695 207.495 2992.865 ;
        RECT 201.885 2992.235 202.055 2992.405 ;
        RECT 207.325 2992.235 207.495 2992.405 ;
        RECT 201.885 2991.775 202.055 2991.945 ;
        RECT 207.325 2991.775 207.495 2991.945 ;
        RECT 201.885 2991.315 202.055 2991.485 ;
        RECT 207.325 2991.315 207.495 2991.485 ;
        RECT 201.885 2990.855 202.055 2991.025 ;
        RECT 207.325 2990.855 207.495 2991.025 ;
      LAYER li1 ;
        RECT 207.325 2990.625 207.495 2990.710 ;
        RECT 207.325 2990.565 208.040 2990.625 ;
      LAYER li1 ;
        RECT 201.885 2990.395 202.055 2990.565 ;
      LAYER li1 ;
        RECT 207.495 2990.395 208.040 2990.565 ;
      LAYER li1 ;
        RECT 201.885 2989.935 202.055 2990.105 ;
        RECT 201.885 2989.475 202.055 2989.645 ;
        RECT 201.885 2989.015 202.055 2989.185 ;
      LAYER li1 ;
        RECT 207.325 2989.040 208.040 2990.395 ;
      LAYER li1 ;
        RECT 201.885 2988.555 202.055 2988.725 ;
      LAYER li1 ;
        RECT 207.325 2988.700 208.870 2989.040 ;
      LAYER li1 ;
        RECT 201.885 2988.095 202.055 2988.265 ;
        RECT 201.885 2987.635 202.055 2987.805 ;
        RECT 201.885 2987.175 202.055 2987.345 ;
        RECT 201.885 2986.715 202.055 2986.885 ;
        RECT 201.885 2986.255 202.055 2986.425 ;
        RECT 201.885 2985.795 202.055 2985.965 ;
        RECT 201.885 2985.335 202.055 2985.505 ;
      LAYER li1 ;
        RECT 207.325 2985.280 208.040 2988.700 ;
        RECT 207.325 2985.190 207.495 2985.280 ;
      LAYER li1 ;
        RECT 201.885 2984.875 202.055 2985.045 ;
        RECT 207.325 2984.875 207.495 2985.045 ;
      LAYER mcon ;
        RECT 207.325 2989.935 207.495 2990.105 ;
        RECT 207.325 2989.475 207.495 2989.645 ;
        RECT 207.325 2989.015 207.495 2989.185 ;
        RECT 207.325 2988.555 207.495 2988.725 ;
        RECT 207.325 2988.095 207.495 2988.265 ;
        RECT 207.325 2987.635 207.495 2987.805 ;
        RECT 207.325 2987.175 207.495 2987.345 ;
        RECT 207.325 2986.715 207.495 2986.885 ;
        RECT 207.325 2986.255 207.495 2986.425 ;
        RECT 207.325 2985.795 207.495 2985.965 ;
        RECT 207.325 2985.335 207.495 2985.505 ;
      LAYER met1 ;
        RECT 201.730 2984.730 202.210 3050.970 ;
        RECT 207.170 2984.730 207.650 3050.970 ;
      LAYER via ;
        RECT 201.855 3023.050 202.155 3024.835 ;
        RECT 207.265 3023.050 207.565 3024.835 ;
      LAYER met2 ;
        RECT 201.770 3023.010 202.200 3024.875 ;
        RECT 207.195 3023.010 207.625 3024.875 ;
      LAYER via2 ;
        RECT 201.855 3023.050 202.155 3024.835 ;
        RECT 207.265 3023.050 207.565 3024.835 ;
      LAYER met3 ;
        RECT 200.115 3023.005 207.640 3024.870 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.760 4456.885 201.930 4457.055 ;
        RECT 207.200 4456.885 207.370 4457.055 ;
        RECT 201.760 4456.425 201.930 4456.595 ;
        RECT 207.200 4456.425 207.370 4456.595 ;
        RECT 201.760 4455.965 201.930 4456.135 ;
        RECT 207.200 4455.965 207.370 4456.135 ;
        RECT 201.760 4455.505 201.930 4455.675 ;
        RECT 207.200 4455.505 207.370 4455.675 ;
        RECT 201.760 4455.045 201.930 4455.215 ;
        RECT 207.200 4455.045 207.370 4455.215 ;
        RECT 201.760 4454.585 201.930 4454.755 ;
        RECT 207.200 4454.585 207.370 4454.755 ;
        RECT 201.760 4454.125 201.930 4454.295 ;
        RECT 207.200 4454.125 207.370 4454.295 ;
        RECT 201.760 4453.665 201.930 4453.835 ;
        RECT 207.200 4453.665 207.370 4453.835 ;
        RECT 201.760 4453.205 201.930 4453.375 ;
        RECT 207.200 4453.205 207.370 4453.375 ;
        RECT 201.760 4452.745 201.930 4452.915 ;
        RECT 207.200 4452.745 207.370 4452.915 ;
        RECT 201.760 4452.285 201.930 4452.455 ;
        RECT 207.200 4452.285 207.370 4452.455 ;
        RECT 201.760 4451.825 201.930 4451.995 ;
        RECT 207.200 4451.825 207.370 4451.995 ;
        RECT 201.760 4451.365 201.930 4451.535 ;
        RECT 207.200 4451.365 207.370 4451.535 ;
        RECT 201.760 4450.905 201.930 4451.075 ;
        RECT 207.200 4450.905 207.370 4451.075 ;
        RECT 201.760 4450.445 201.930 4450.615 ;
        RECT 207.200 4450.445 207.370 4450.615 ;
        RECT 201.760 4449.985 201.930 4450.155 ;
        RECT 207.200 4449.985 207.370 4450.155 ;
        RECT 201.760 4449.525 201.930 4449.695 ;
        RECT 207.200 4449.525 207.370 4449.695 ;
        RECT 201.760 4449.065 201.930 4449.235 ;
        RECT 207.200 4449.065 207.370 4449.235 ;
        RECT 201.760 4448.605 201.930 4448.775 ;
        RECT 207.200 4448.605 207.370 4448.775 ;
        RECT 201.760 4448.145 201.930 4448.315 ;
        RECT 207.200 4448.145 207.370 4448.315 ;
        RECT 201.760 4447.685 201.930 4447.855 ;
        RECT 207.200 4447.685 207.370 4447.855 ;
        RECT 201.760 4447.225 201.930 4447.395 ;
        RECT 207.200 4447.225 207.370 4447.395 ;
        RECT 201.760 4446.765 201.930 4446.935 ;
        RECT 207.200 4446.765 207.370 4446.935 ;
        RECT 201.760 4446.305 201.930 4446.475 ;
        RECT 207.200 4446.305 207.370 4446.475 ;
        RECT 201.760 4445.845 201.930 4446.015 ;
        RECT 207.200 4445.845 207.370 4446.015 ;
        RECT 201.760 4445.385 201.930 4445.555 ;
        RECT 207.200 4445.385 207.370 4445.555 ;
        RECT 201.760 4444.925 201.930 4445.095 ;
        RECT 207.200 4444.925 207.370 4445.095 ;
        RECT 201.760 4444.465 201.930 4444.635 ;
        RECT 207.200 4444.465 207.370 4444.635 ;
        RECT 201.760 4444.005 201.930 4444.175 ;
        RECT 207.200 4444.005 207.370 4444.175 ;
        RECT 201.760 4443.545 201.930 4443.715 ;
        RECT 207.200 4443.545 207.370 4443.715 ;
        RECT 201.760 4443.085 201.930 4443.255 ;
        RECT 207.200 4443.085 207.370 4443.255 ;
        RECT 201.760 4442.625 201.930 4442.795 ;
        RECT 207.200 4442.625 207.370 4442.795 ;
        RECT 201.760 4442.165 201.930 4442.335 ;
        RECT 207.200 4442.165 207.370 4442.335 ;
        RECT 201.760 4441.705 201.930 4441.875 ;
        RECT 207.200 4441.705 207.370 4441.875 ;
        RECT 201.760 4441.245 201.930 4441.415 ;
        RECT 207.200 4441.245 207.370 4441.415 ;
        RECT 201.760 4440.785 201.930 4440.955 ;
        RECT 207.200 4440.785 207.370 4440.955 ;
        RECT 201.760 4440.325 201.930 4440.495 ;
        RECT 207.200 4440.325 207.370 4440.495 ;
        RECT 201.760 4439.865 201.930 4440.035 ;
        RECT 207.200 4439.865 207.370 4440.035 ;
        RECT 201.760 4439.405 201.930 4439.575 ;
        RECT 207.200 4439.405 207.370 4439.575 ;
        RECT 201.760 4438.945 201.930 4439.115 ;
        RECT 207.200 4438.945 207.370 4439.115 ;
        RECT 201.760 4438.485 201.930 4438.655 ;
        RECT 207.200 4438.485 207.370 4438.655 ;
        RECT 201.760 4438.025 201.930 4438.195 ;
        RECT 207.200 4438.025 207.370 4438.195 ;
        RECT 201.760 4437.565 201.930 4437.735 ;
        RECT 207.200 4437.565 207.370 4437.735 ;
        RECT 201.760 4437.105 201.930 4437.275 ;
        RECT 207.200 4437.105 207.370 4437.275 ;
        RECT 201.760 4436.645 201.930 4436.815 ;
        RECT 207.200 4436.645 207.370 4436.815 ;
        RECT 201.760 4436.185 201.930 4436.355 ;
        RECT 207.200 4436.185 207.370 4436.355 ;
        RECT 201.760 4435.725 201.930 4435.895 ;
        RECT 207.200 4435.725 207.370 4435.895 ;
        RECT 201.760 4435.265 201.930 4435.435 ;
        RECT 207.200 4435.265 207.370 4435.435 ;
        RECT 201.760 4434.805 201.930 4434.975 ;
        RECT 207.200 4434.805 207.370 4434.975 ;
        RECT 201.760 4434.345 201.930 4434.515 ;
        RECT 207.200 4434.345 207.370 4434.515 ;
        RECT 201.760 4433.885 201.930 4434.055 ;
        RECT 207.200 4433.885 207.370 4434.055 ;
        RECT 201.760 4433.425 201.930 4433.595 ;
        RECT 207.200 4433.425 207.370 4433.595 ;
        RECT 201.760 4432.965 201.930 4433.135 ;
        RECT 207.200 4432.965 207.370 4433.135 ;
        RECT 201.760 4432.505 201.930 4432.675 ;
        RECT 207.200 4432.505 207.370 4432.675 ;
        RECT 201.760 4432.045 201.930 4432.215 ;
        RECT 207.200 4432.045 207.370 4432.215 ;
        RECT 201.760 4431.585 201.930 4431.755 ;
        RECT 207.200 4431.585 207.370 4431.755 ;
        RECT 201.760 4431.125 201.930 4431.295 ;
        RECT 207.200 4431.125 207.370 4431.295 ;
        RECT 201.760 4430.665 201.930 4430.835 ;
        RECT 207.200 4430.665 207.370 4430.835 ;
        RECT 201.760 4430.205 201.930 4430.375 ;
        RECT 207.200 4430.205 207.370 4430.375 ;
        RECT 201.760 4429.745 201.930 4429.915 ;
        RECT 207.200 4429.745 207.370 4429.915 ;
        RECT 201.760 4429.285 201.930 4429.455 ;
        RECT 207.200 4429.285 207.370 4429.455 ;
        RECT 201.760 4428.825 201.930 4428.995 ;
        RECT 207.200 4428.825 207.370 4428.995 ;
        RECT 201.760 4428.365 201.930 4428.535 ;
        RECT 207.200 4428.365 207.370 4428.535 ;
        RECT 201.760 4427.905 201.930 4428.075 ;
        RECT 207.200 4427.905 207.370 4428.075 ;
        RECT 201.760 4427.445 201.930 4427.615 ;
        RECT 207.200 4427.445 207.370 4427.615 ;
        RECT 201.760 4426.985 201.930 4427.155 ;
        RECT 207.200 4426.985 207.370 4427.155 ;
      LAYER met1 ;
        RECT 201.605 4426.840 202.085 4457.200 ;
        RECT 207.045 4426.840 207.525 4457.200 ;
      LAYER via ;
        RECT 201.700 4446.920 202.000 4448.705 ;
        RECT 207.110 4446.920 207.410 4448.705 ;
      LAYER met2 ;
        RECT 201.615 4446.880 202.045 4448.745 ;
        RECT 207.040 4446.880 207.470 4448.745 ;
      LAYER via2 ;
        RECT 201.700 4446.920 202.000 4448.705 ;
        RECT 207.110 4446.920 207.410 4448.705 ;
      LAYER met3 ;
        RECT 199.960 4446.875 207.485 4448.740 ;
    END
  END vssd
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 2082.975 4984.895 2083.145 4985.065 ;
        RECT 2083.435 4984.895 2083.605 4985.065 ;
        RECT 2083.895 4984.895 2084.065 4985.065 ;
        RECT 2084.355 4984.895 2084.525 4985.065 ;
        RECT 2084.815 4984.895 2084.985 4985.065 ;
        RECT 2085.275 4984.895 2085.445 4985.065 ;
        RECT 2085.735 4984.895 2085.905 4985.065 ;
        RECT 2086.195 4984.895 2086.365 4985.065 ;
        RECT 2086.655 4984.895 2086.825 4985.065 ;
        RECT 2087.115 4984.895 2087.285 4985.065 ;
        RECT 2087.575 4984.895 2087.745 4985.065 ;
        RECT 2088.035 4984.895 2088.205 4985.065 ;
        RECT 2088.495 4984.895 2088.665 4985.065 ;
        RECT 2088.955 4984.895 2089.125 4985.065 ;
      LAYER li1 ;
        RECT 2084.970 4980.060 2085.320 4981.310 ;
        RECT 2083.380 4979.625 2088.725 4980.060 ;
      LAYER li1 ;
        RECT 2082.975 4979.455 2083.145 4979.625 ;
      LAYER li1 ;
        RECT 2083.290 4979.455 2088.810 4979.625 ;
      LAYER li1 ;
        RECT 2088.955 4979.455 2089.125 4979.625 ;
      LAYER mcon ;
        RECT 2083.435 4979.455 2083.605 4979.625 ;
        RECT 2083.895 4979.455 2084.065 4979.625 ;
        RECT 2084.355 4979.455 2084.525 4979.625 ;
        RECT 2084.815 4979.455 2084.985 4979.625 ;
        RECT 2085.275 4979.455 2085.445 4979.625 ;
        RECT 2085.735 4979.455 2085.905 4979.625 ;
        RECT 2086.195 4979.455 2086.365 4979.625 ;
        RECT 2086.655 4979.455 2086.825 4979.625 ;
        RECT 2087.115 4979.455 2087.285 4979.625 ;
        RECT 2087.575 4979.455 2087.745 4979.625 ;
        RECT 2088.035 4979.455 2088.205 4979.625 ;
      LAYER met1 ;
        RECT 2082.830 4984.740 2092.990 4985.220 ;
        RECT 2082.830 4979.300 2092.990 4979.780 ;
      LAYER via ;
        RECT 2091.115 4984.830 2092.900 4985.130 ;
        RECT 2091.115 4979.390 2092.900 4979.690 ;
      LAYER met2 ;
        RECT 2091.075 4984.760 2092.940 4985.190 ;
        RECT 2091.075 4979.320 2092.940 4979.750 ;
      LAYER via2 ;
        RECT 2091.115 4984.830 2092.900 4985.130 ;
        RECT 2091.115 4979.390 2092.900 4979.690 ;
      LAYER met3 ;
        RECT 2091.080 4979.320 2092.930 4989.575 ;
    END
    PORT
      LAYER li1 ;
        RECT 834.795 4983.270 834.965 4983.440 ;
        RECT 835.255 4983.270 835.425 4983.440 ;
        RECT 835.715 4983.270 835.885 4983.440 ;
        RECT 836.175 4983.270 836.345 4983.440 ;
        RECT 836.635 4983.270 836.805 4983.440 ;
        RECT 837.095 4983.270 837.265 4983.440 ;
        RECT 837.555 4983.270 837.725 4983.440 ;
        RECT 838.015 4983.270 838.185 4983.440 ;
        RECT 838.475 4983.270 838.645 4983.440 ;
        RECT 838.935 4983.270 839.105 4983.440 ;
        RECT 839.395 4983.270 839.565 4983.440 ;
        RECT 839.855 4983.270 840.025 4983.440 ;
        RECT 840.315 4983.270 840.485 4983.440 ;
        RECT 840.775 4983.270 840.945 4983.440 ;
        RECT 841.235 4983.270 841.405 4983.440 ;
        RECT 841.695 4983.270 841.865 4983.440 ;
        RECT 842.155 4983.270 842.325 4983.440 ;
        RECT 842.615 4983.270 842.785 4983.440 ;
        RECT 843.075 4983.270 843.245 4983.440 ;
        RECT 843.535 4983.270 843.705 4983.440 ;
        RECT 843.995 4983.270 844.165 4983.440 ;
        RECT 844.455 4983.270 844.625 4983.440 ;
        RECT 844.915 4983.270 845.085 4983.440 ;
        RECT 845.375 4983.270 845.545 4983.440 ;
        RECT 845.835 4983.270 846.005 4983.440 ;
        RECT 846.295 4983.270 846.465 4983.440 ;
        RECT 846.755 4983.270 846.925 4983.440 ;
        RECT 847.215 4983.270 847.385 4983.440 ;
        RECT 847.675 4983.270 847.845 4983.440 ;
        RECT 848.135 4983.270 848.305 4983.440 ;
        RECT 848.595 4983.270 848.765 4983.440 ;
        RECT 849.055 4983.270 849.225 4983.440 ;
        RECT 849.515 4983.270 849.685 4983.440 ;
        RECT 849.975 4983.270 850.145 4983.440 ;
        RECT 850.435 4983.270 850.605 4983.440 ;
        RECT 850.895 4983.270 851.065 4983.440 ;
        RECT 851.355 4983.270 851.525 4983.440 ;
        RECT 851.815 4983.270 851.985 4983.440 ;
        RECT 852.275 4983.270 852.445 4983.440 ;
        RECT 852.735 4983.270 852.905 4983.440 ;
      LAYER li1 ;
        RECT 836.790 4978.435 837.140 4979.685 ;
        RECT 842.770 4978.435 843.120 4979.685 ;
        RECT 848.750 4978.435 849.100 4979.685 ;
        RECT 835.200 4978.000 840.545 4978.435 ;
        RECT 841.180 4978.000 846.525 4978.435 ;
        RECT 847.160 4978.000 852.505 4978.435 ;
      LAYER li1 ;
        RECT 834.795 4977.830 834.965 4978.000 ;
      LAYER li1 ;
        RECT 835.110 4977.830 840.630 4978.000 ;
      LAYER li1 ;
        RECT 840.775 4977.830 840.945 4978.000 ;
      LAYER li1 ;
        RECT 841.090 4977.830 846.610 4978.000 ;
      LAYER li1 ;
        RECT 846.755 4977.830 846.925 4978.000 ;
      LAYER li1 ;
        RECT 847.070 4977.830 852.590 4978.000 ;
      LAYER li1 ;
        RECT 852.735 4977.830 852.905 4978.000 ;
      LAYER mcon ;
        RECT 835.255 4977.830 835.425 4978.000 ;
        RECT 835.715 4977.830 835.885 4978.000 ;
        RECT 836.175 4977.830 836.345 4978.000 ;
        RECT 836.635 4977.830 836.805 4978.000 ;
        RECT 837.095 4977.830 837.265 4978.000 ;
        RECT 837.555 4977.830 837.725 4978.000 ;
        RECT 838.015 4977.830 838.185 4978.000 ;
        RECT 838.475 4977.830 838.645 4978.000 ;
        RECT 838.935 4977.830 839.105 4978.000 ;
        RECT 839.395 4977.830 839.565 4978.000 ;
        RECT 839.855 4977.830 840.025 4978.000 ;
        RECT 841.235 4977.830 841.405 4978.000 ;
        RECT 841.695 4977.830 841.865 4978.000 ;
        RECT 842.155 4977.830 842.325 4978.000 ;
        RECT 842.615 4977.830 842.785 4978.000 ;
        RECT 843.075 4977.830 843.245 4978.000 ;
        RECT 843.535 4977.830 843.705 4978.000 ;
        RECT 843.995 4977.830 844.165 4978.000 ;
        RECT 844.455 4977.830 844.625 4978.000 ;
        RECT 844.915 4977.830 845.085 4978.000 ;
        RECT 845.375 4977.830 845.545 4978.000 ;
        RECT 845.835 4977.830 846.005 4978.000 ;
        RECT 847.215 4977.830 847.385 4978.000 ;
        RECT 847.675 4977.830 847.845 4978.000 ;
        RECT 848.135 4977.830 848.305 4978.000 ;
        RECT 848.595 4977.830 848.765 4978.000 ;
        RECT 849.055 4977.830 849.225 4978.000 ;
        RECT 849.515 4977.830 849.685 4978.000 ;
        RECT 849.975 4977.830 850.145 4978.000 ;
        RECT 850.435 4977.830 850.605 4978.000 ;
        RECT 850.895 4977.830 851.065 4978.000 ;
        RECT 851.355 4977.830 851.525 4978.000 ;
        RECT 851.815 4977.830 851.985 4978.000 ;
      LAYER met1 ;
        RECT 834.650 4983.115 853.050 4983.595 ;
        RECT 834.650 4977.675 853.050 4978.155 ;
      LAYER via ;
        RECT 848.930 4983.185 850.715 4983.485 ;
        RECT 848.930 4977.745 850.715 4978.045 ;
      LAYER met2 ;
        RECT 848.890 4983.115 850.755 4983.545 ;
        RECT 848.890 4977.675 850.755 4978.105 ;
      LAYER via2 ;
        RECT 848.930 4983.185 850.715 4983.485 ;
        RECT 848.930 4977.745 850.715 4978.045 ;
      LAYER met3 ;
        RECT 848.895 4977.675 850.745 4987.930 ;
    END
    PORT
      LAYER li1 ;
        RECT 3309.980 4984.485 3310.150 4984.655 ;
        RECT 3310.440 4984.485 3310.610 4984.655 ;
        RECT 3310.900 4984.485 3311.070 4984.655 ;
        RECT 3311.360 4984.485 3311.530 4984.655 ;
        RECT 3311.820 4984.485 3311.990 4984.655 ;
        RECT 3312.280 4984.485 3312.450 4984.655 ;
        RECT 3312.740 4984.485 3312.910 4984.655 ;
        RECT 3313.200 4984.485 3313.370 4984.655 ;
        RECT 3313.660 4984.485 3313.830 4984.655 ;
        RECT 3314.120 4984.485 3314.290 4984.655 ;
        RECT 3314.580 4984.485 3314.750 4984.655 ;
        RECT 3315.040 4984.485 3315.210 4984.655 ;
        RECT 3315.500 4984.485 3315.670 4984.655 ;
        RECT 3315.960 4984.485 3316.130 4984.655 ;
        RECT 3316.420 4984.485 3316.590 4984.655 ;
        RECT 3316.880 4984.485 3317.050 4984.655 ;
        RECT 3317.340 4984.485 3317.510 4984.655 ;
        RECT 3317.800 4984.485 3317.970 4984.655 ;
        RECT 3318.260 4984.485 3318.430 4984.655 ;
        RECT 3318.720 4984.485 3318.890 4984.655 ;
        RECT 3319.180 4984.485 3319.350 4984.655 ;
        RECT 3319.640 4984.485 3319.810 4984.655 ;
        RECT 3320.100 4984.485 3320.270 4984.655 ;
        RECT 3320.560 4984.485 3320.730 4984.655 ;
        RECT 3321.020 4984.485 3321.190 4984.655 ;
        RECT 3321.480 4984.485 3321.650 4984.655 ;
        RECT 3321.940 4984.485 3322.110 4984.655 ;
        RECT 3322.400 4984.485 3322.570 4984.655 ;
        RECT 3322.860 4984.485 3323.030 4984.655 ;
        RECT 3323.320 4984.485 3323.490 4984.655 ;
        RECT 3323.780 4984.485 3323.950 4984.655 ;
        RECT 3324.240 4984.485 3324.410 4984.655 ;
        RECT 3324.700 4984.485 3324.870 4984.655 ;
        RECT 3325.160 4984.485 3325.330 4984.655 ;
        RECT 3325.620 4984.485 3325.790 4984.655 ;
        RECT 3326.080 4984.485 3326.250 4984.655 ;
        RECT 3326.540 4984.485 3326.710 4984.655 ;
        RECT 3327.000 4984.485 3327.170 4984.655 ;
        RECT 3327.460 4984.485 3327.630 4984.655 ;
        RECT 3327.920 4984.485 3328.090 4984.655 ;
        RECT 3328.380 4984.485 3328.550 4984.655 ;
        RECT 3328.840 4984.485 3329.010 4984.655 ;
        RECT 3329.300 4984.485 3329.470 4984.655 ;
        RECT 3329.760 4984.485 3329.930 4984.655 ;
        RECT 3330.220 4984.485 3330.390 4984.655 ;
        RECT 3330.680 4984.485 3330.850 4984.655 ;
        RECT 3331.140 4984.485 3331.310 4984.655 ;
        RECT 3331.600 4984.485 3331.770 4984.655 ;
        RECT 3332.060 4984.485 3332.230 4984.655 ;
        RECT 3332.520 4984.485 3332.690 4984.655 ;
        RECT 3332.980 4984.485 3333.150 4984.655 ;
        RECT 3333.440 4984.485 3333.610 4984.655 ;
        RECT 3333.900 4984.485 3334.070 4984.655 ;
      LAYER li1 ;
        RECT 3311.975 4979.650 3312.325 4980.900 ;
        RECT 3317.955 4979.650 3318.305 4980.900 ;
        RECT 3323.935 4979.650 3324.285 4980.900 ;
        RECT 3329.915 4979.650 3330.265 4980.900 ;
        RECT 3310.385 4979.215 3315.730 4979.650 ;
        RECT 3316.365 4979.215 3321.710 4979.650 ;
        RECT 3322.345 4979.215 3327.690 4979.650 ;
        RECT 3328.325 4979.215 3333.670 4979.650 ;
      LAYER li1 ;
        RECT 3309.980 4979.045 3310.150 4979.215 ;
      LAYER li1 ;
        RECT 3310.295 4979.045 3315.815 4979.215 ;
      LAYER li1 ;
        RECT 3315.960 4979.045 3316.130 4979.215 ;
      LAYER li1 ;
        RECT 3316.275 4979.045 3321.795 4979.215 ;
      LAYER li1 ;
        RECT 3321.940 4979.045 3322.110 4979.215 ;
      LAYER li1 ;
        RECT 3322.255 4979.045 3327.775 4979.215 ;
      LAYER li1 ;
        RECT 3327.920 4979.045 3328.090 4979.215 ;
      LAYER li1 ;
        RECT 3328.235 4979.045 3333.755 4979.215 ;
      LAYER li1 ;
        RECT 3333.900 4979.045 3334.070 4979.215 ;
      LAYER mcon ;
        RECT 3310.440 4979.045 3310.610 4979.215 ;
        RECT 3310.900 4979.045 3311.070 4979.215 ;
        RECT 3311.360 4979.045 3311.530 4979.215 ;
        RECT 3311.820 4979.045 3311.990 4979.215 ;
        RECT 3312.280 4979.045 3312.450 4979.215 ;
        RECT 3312.740 4979.045 3312.910 4979.215 ;
        RECT 3313.200 4979.045 3313.370 4979.215 ;
        RECT 3313.660 4979.045 3313.830 4979.215 ;
        RECT 3314.120 4979.045 3314.290 4979.215 ;
        RECT 3314.580 4979.045 3314.750 4979.215 ;
        RECT 3315.040 4979.045 3315.210 4979.215 ;
        RECT 3316.420 4979.045 3316.590 4979.215 ;
        RECT 3316.880 4979.045 3317.050 4979.215 ;
        RECT 3317.340 4979.045 3317.510 4979.215 ;
        RECT 3317.800 4979.045 3317.970 4979.215 ;
        RECT 3318.260 4979.045 3318.430 4979.215 ;
        RECT 3318.720 4979.045 3318.890 4979.215 ;
        RECT 3319.180 4979.045 3319.350 4979.215 ;
        RECT 3319.640 4979.045 3319.810 4979.215 ;
        RECT 3320.100 4979.045 3320.270 4979.215 ;
        RECT 3320.560 4979.045 3320.730 4979.215 ;
        RECT 3321.020 4979.045 3321.190 4979.215 ;
        RECT 3322.400 4979.045 3322.570 4979.215 ;
        RECT 3322.860 4979.045 3323.030 4979.215 ;
        RECT 3323.320 4979.045 3323.490 4979.215 ;
        RECT 3323.780 4979.045 3323.950 4979.215 ;
        RECT 3324.240 4979.045 3324.410 4979.215 ;
        RECT 3324.700 4979.045 3324.870 4979.215 ;
        RECT 3325.160 4979.045 3325.330 4979.215 ;
        RECT 3325.620 4979.045 3325.790 4979.215 ;
        RECT 3326.080 4979.045 3326.250 4979.215 ;
        RECT 3326.540 4979.045 3326.710 4979.215 ;
        RECT 3327.000 4979.045 3327.170 4979.215 ;
        RECT 3328.380 4979.045 3328.550 4979.215 ;
        RECT 3328.840 4979.045 3329.010 4979.215 ;
        RECT 3329.300 4979.045 3329.470 4979.215 ;
        RECT 3329.760 4979.045 3329.930 4979.215 ;
        RECT 3330.220 4979.045 3330.390 4979.215 ;
        RECT 3330.680 4979.045 3330.850 4979.215 ;
        RECT 3331.140 4979.045 3331.310 4979.215 ;
        RECT 3331.600 4979.045 3331.770 4979.215 ;
        RECT 3332.060 4979.045 3332.230 4979.215 ;
        RECT 3332.520 4979.045 3332.690 4979.215 ;
        RECT 3332.980 4979.045 3333.150 4979.215 ;
      LAYER met1 ;
        RECT 3309.835 4984.330 3334.215 4984.810 ;
        RECT 3309.835 4978.890 3334.215 4979.370 ;
      LAYER via ;
        RECT 3324.165 4984.420 3325.950 4984.720 ;
        RECT 3324.165 4978.980 3325.950 4979.280 ;
      LAYER met2 ;
        RECT 3324.125 4984.350 3325.990 4984.780 ;
        RECT 3324.125 4978.910 3325.990 4979.340 ;
      LAYER via2 ;
        RECT 3324.165 4984.420 3325.950 4984.720 ;
        RECT 3324.165 4978.980 3325.950 4979.280 ;
      LAYER met3 ;
        RECT 3324.130 4978.910 3325.980 4989.165 ;
    END
    PORT
      LAYER li1 ;
        RECT 3377.780 2267.965 3377.950 2268.135 ;
        RECT 3383.220 2267.965 3383.390 2268.135 ;
      LAYER li1 ;
        RECT 3377.780 2267.735 3377.950 2267.820 ;
        RECT 3377.780 2264.330 3378.385 2267.735 ;
      LAYER li1 ;
        RECT 3383.220 2267.505 3383.390 2267.675 ;
        RECT 3383.220 2267.045 3383.390 2267.215 ;
        RECT 3383.220 2266.585 3383.390 2266.755 ;
        RECT 3383.220 2266.125 3383.390 2266.295 ;
        RECT 3383.220 2265.665 3383.390 2265.835 ;
        RECT 3383.220 2265.205 3383.390 2265.375 ;
        RECT 3383.220 2264.745 3383.390 2264.915 ;
      LAYER li1 ;
        RECT 3377.780 2263.980 3379.635 2264.330 ;
      LAYER li1 ;
        RECT 3383.220 2264.285 3383.390 2264.455 ;
      LAYER li1 ;
        RECT 3377.780 2262.390 3378.385 2263.980 ;
      LAYER li1 ;
        RECT 3383.220 2263.825 3383.390 2263.995 ;
        RECT 3383.220 2263.365 3383.390 2263.535 ;
        RECT 3383.220 2262.905 3383.390 2263.075 ;
        RECT 3383.220 2262.445 3383.390 2262.615 ;
      LAYER li1 ;
        RECT 3377.780 2262.300 3377.950 2262.390 ;
      LAYER li1 ;
        RECT 3377.780 2261.985 3377.950 2262.155 ;
        RECT 3383.220 2261.985 3383.390 2262.155 ;
      LAYER li1 ;
        RECT 3377.780 2261.755 3377.950 2261.840 ;
        RECT 3377.780 2258.350 3378.385 2261.755 ;
      LAYER li1 ;
        RECT 3383.220 2261.525 3383.390 2261.695 ;
        RECT 3383.220 2261.065 3383.390 2261.235 ;
        RECT 3383.220 2260.605 3383.390 2260.775 ;
        RECT 3383.220 2260.145 3383.390 2260.315 ;
        RECT 3383.220 2259.685 3383.390 2259.855 ;
        RECT 3383.220 2259.225 3383.390 2259.395 ;
        RECT 3383.220 2258.765 3383.390 2258.935 ;
      LAYER li1 ;
        RECT 3377.780 2258.000 3379.635 2258.350 ;
      LAYER li1 ;
        RECT 3383.220 2258.305 3383.390 2258.475 ;
      LAYER li1 ;
        RECT 3377.780 2256.410 3378.385 2258.000 ;
      LAYER li1 ;
        RECT 3383.220 2257.845 3383.390 2258.015 ;
        RECT 3383.220 2257.385 3383.390 2257.555 ;
        RECT 3383.220 2256.925 3383.390 2257.095 ;
        RECT 3383.220 2256.465 3383.390 2256.635 ;
      LAYER li1 ;
        RECT 3377.780 2256.320 3377.950 2256.410 ;
      LAYER li1 ;
        RECT 3377.780 2256.005 3377.950 2256.175 ;
        RECT 3383.220 2256.005 3383.390 2256.175 ;
      LAYER li1 ;
        RECT 3377.780 2255.775 3377.950 2255.860 ;
        RECT 3377.780 2252.370 3378.385 2255.775 ;
      LAYER li1 ;
        RECT 3383.220 2255.545 3383.390 2255.715 ;
        RECT 3383.220 2255.085 3383.390 2255.255 ;
        RECT 3383.220 2254.625 3383.390 2254.795 ;
        RECT 3383.220 2254.165 3383.390 2254.335 ;
        RECT 3383.220 2253.705 3383.390 2253.875 ;
        RECT 3383.220 2253.245 3383.390 2253.415 ;
        RECT 3383.220 2252.785 3383.390 2252.955 ;
      LAYER li1 ;
        RECT 3377.780 2252.020 3379.635 2252.370 ;
      LAYER li1 ;
        RECT 3383.220 2252.325 3383.390 2252.495 ;
      LAYER li1 ;
        RECT 3377.780 2250.430 3378.385 2252.020 ;
      LAYER li1 ;
        RECT 3383.220 2251.865 3383.390 2252.035 ;
        RECT 3383.220 2251.405 3383.390 2251.575 ;
        RECT 3383.220 2250.945 3383.390 2251.115 ;
        RECT 3383.220 2250.485 3383.390 2250.655 ;
      LAYER li1 ;
        RECT 3377.780 2250.340 3377.950 2250.430 ;
      LAYER li1 ;
        RECT 3377.780 2250.025 3377.950 2250.195 ;
        RECT 3383.220 2250.025 3383.390 2250.195 ;
      LAYER li1 ;
        RECT 3377.780 2249.795 3377.950 2249.880 ;
        RECT 3377.780 2246.390 3378.385 2249.795 ;
      LAYER li1 ;
        RECT 3383.220 2249.565 3383.390 2249.735 ;
        RECT 3383.220 2249.105 3383.390 2249.275 ;
        RECT 3383.220 2248.645 3383.390 2248.815 ;
        RECT 3383.220 2248.185 3383.390 2248.355 ;
        RECT 3383.220 2247.725 3383.390 2247.895 ;
        RECT 3383.220 2247.265 3383.390 2247.435 ;
        RECT 3383.220 2246.805 3383.390 2246.975 ;
      LAYER li1 ;
        RECT 3377.780 2246.040 3379.635 2246.390 ;
      LAYER li1 ;
        RECT 3383.220 2246.345 3383.390 2246.515 ;
      LAYER li1 ;
        RECT 3377.780 2244.450 3378.385 2246.040 ;
      LAYER li1 ;
        RECT 3383.220 2245.885 3383.390 2246.055 ;
        RECT 3383.220 2245.425 3383.390 2245.595 ;
        RECT 3383.220 2244.965 3383.390 2245.135 ;
        RECT 3383.220 2244.505 3383.390 2244.675 ;
      LAYER li1 ;
        RECT 3377.780 2244.360 3377.950 2244.450 ;
      LAYER li1 ;
        RECT 3377.780 2244.045 3377.950 2244.215 ;
        RECT 3383.220 2244.045 3383.390 2244.215 ;
      LAYER li1 ;
        RECT 3377.780 2243.815 3377.950 2243.900 ;
        RECT 3377.780 2240.410 3378.385 2243.815 ;
      LAYER li1 ;
        RECT 3383.220 2243.585 3383.390 2243.755 ;
        RECT 3383.220 2243.125 3383.390 2243.295 ;
        RECT 3383.220 2242.665 3383.390 2242.835 ;
        RECT 3383.220 2242.205 3383.390 2242.375 ;
        RECT 3383.220 2241.745 3383.390 2241.915 ;
        RECT 3383.220 2241.285 3383.390 2241.455 ;
        RECT 3383.220 2240.825 3383.390 2240.995 ;
      LAYER li1 ;
        RECT 3377.780 2240.060 3379.635 2240.410 ;
      LAYER li1 ;
        RECT 3383.220 2240.365 3383.390 2240.535 ;
      LAYER li1 ;
        RECT 3377.780 2238.470 3378.385 2240.060 ;
      LAYER li1 ;
        RECT 3383.220 2239.905 3383.390 2240.075 ;
        RECT 3383.220 2239.445 3383.390 2239.615 ;
        RECT 3383.220 2238.985 3383.390 2239.155 ;
        RECT 3383.220 2238.525 3383.390 2238.695 ;
      LAYER li1 ;
        RECT 3377.780 2238.380 3377.950 2238.470 ;
      LAYER li1 ;
        RECT 3377.780 2238.065 3377.950 2238.235 ;
        RECT 3383.220 2238.065 3383.390 2238.235 ;
      LAYER li1 ;
        RECT 3377.780 2237.835 3377.950 2237.920 ;
        RECT 3377.780 2234.430 3378.385 2237.835 ;
      LAYER li1 ;
        RECT 3383.220 2237.605 3383.390 2237.775 ;
        RECT 3383.220 2237.145 3383.390 2237.315 ;
        RECT 3383.220 2236.685 3383.390 2236.855 ;
        RECT 3383.220 2236.225 3383.390 2236.395 ;
        RECT 3383.220 2235.765 3383.390 2235.935 ;
        RECT 3383.220 2235.305 3383.390 2235.475 ;
        RECT 3383.220 2234.845 3383.390 2235.015 ;
      LAYER li1 ;
        RECT 3377.780 2234.080 3379.635 2234.430 ;
      LAYER li1 ;
        RECT 3383.220 2234.385 3383.390 2234.555 ;
      LAYER li1 ;
        RECT 3377.780 2232.490 3378.385 2234.080 ;
      LAYER li1 ;
        RECT 3383.220 2233.925 3383.390 2234.095 ;
        RECT 3383.220 2233.465 3383.390 2233.635 ;
        RECT 3383.220 2233.005 3383.390 2233.175 ;
        RECT 3383.220 2232.545 3383.390 2232.715 ;
      LAYER li1 ;
        RECT 3377.780 2232.400 3377.950 2232.490 ;
      LAYER li1 ;
        RECT 3377.780 2232.085 3377.950 2232.255 ;
        RECT 3383.220 2232.085 3383.390 2232.255 ;
      LAYER li1 ;
        RECT 3377.780 2231.855 3377.950 2231.940 ;
        RECT 3377.780 2228.450 3378.385 2231.855 ;
      LAYER li1 ;
        RECT 3383.220 2231.625 3383.390 2231.795 ;
        RECT 3383.220 2231.165 3383.390 2231.335 ;
        RECT 3383.220 2230.705 3383.390 2230.875 ;
        RECT 3383.220 2230.245 3383.390 2230.415 ;
        RECT 3383.220 2229.785 3383.390 2229.955 ;
        RECT 3383.220 2229.325 3383.390 2229.495 ;
        RECT 3383.220 2228.865 3383.390 2229.035 ;
      LAYER li1 ;
        RECT 3377.780 2228.100 3379.635 2228.450 ;
      LAYER li1 ;
        RECT 3383.220 2228.405 3383.390 2228.575 ;
      LAYER li1 ;
        RECT 3377.780 2226.510 3378.385 2228.100 ;
      LAYER li1 ;
        RECT 3383.220 2227.945 3383.390 2228.115 ;
        RECT 3383.220 2227.485 3383.390 2227.655 ;
        RECT 3383.220 2227.025 3383.390 2227.195 ;
        RECT 3383.220 2226.565 3383.390 2226.735 ;
      LAYER li1 ;
        RECT 3377.780 2226.420 3377.950 2226.510 ;
      LAYER li1 ;
        RECT 3377.780 2226.105 3377.950 2226.275 ;
        RECT 3383.220 2226.105 3383.390 2226.275 ;
      LAYER li1 ;
        RECT 3377.780 2225.875 3377.950 2225.960 ;
        RECT 3377.780 2222.470 3378.385 2225.875 ;
      LAYER li1 ;
        RECT 3383.220 2225.645 3383.390 2225.815 ;
        RECT 3383.220 2225.185 3383.390 2225.355 ;
        RECT 3383.220 2224.725 3383.390 2224.895 ;
        RECT 3383.220 2224.265 3383.390 2224.435 ;
        RECT 3383.220 2223.805 3383.390 2223.975 ;
        RECT 3383.220 2223.345 3383.390 2223.515 ;
        RECT 3383.220 2222.885 3383.390 2223.055 ;
      LAYER li1 ;
        RECT 3377.780 2222.120 3379.635 2222.470 ;
      LAYER li1 ;
        RECT 3383.220 2222.425 3383.390 2222.595 ;
      LAYER li1 ;
        RECT 3377.780 2220.530 3378.385 2222.120 ;
      LAYER li1 ;
        RECT 3383.220 2221.965 3383.390 2222.135 ;
        RECT 3383.220 2221.505 3383.390 2221.675 ;
        RECT 3383.220 2221.045 3383.390 2221.215 ;
        RECT 3383.220 2220.585 3383.390 2220.755 ;
      LAYER li1 ;
        RECT 3377.780 2220.440 3377.950 2220.530 ;
      LAYER li1 ;
        RECT 3377.780 2220.125 3377.950 2220.295 ;
        RECT 3383.220 2220.125 3383.390 2220.295 ;
      LAYER li1 ;
        RECT 3377.780 2219.895 3377.950 2219.980 ;
        RECT 3377.780 2216.490 3378.385 2219.895 ;
      LAYER li1 ;
        RECT 3383.220 2219.665 3383.390 2219.835 ;
        RECT 3383.220 2219.205 3383.390 2219.375 ;
        RECT 3383.220 2218.745 3383.390 2218.915 ;
        RECT 3383.220 2218.285 3383.390 2218.455 ;
        RECT 3383.220 2217.825 3383.390 2217.995 ;
        RECT 3383.220 2217.365 3383.390 2217.535 ;
        RECT 3383.220 2216.905 3383.390 2217.075 ;
      LAYER li1 ;
        RECT 3377.780 2216.140 3379.635 2216.490 ;
      LAYER li1 ;
        RECT 3383.220 2216.445 3383.390 2216.615 ;
      LAYER li1 ;
        RECT 3377.780 2214.550 3378.385 2216.140 ;
      LAYER li1 ;
        RECT 3383.220 2215.985 3383.390 2216.155 ;
        RECT 3383.220 2215.525 3383.390 2215.695 ;
        RECT 3383.220 2215.065 3383.390 2215.235 ;
        RECT 3383.220 2214.605 3383.390 2214.775 ;
      LAYER li1 ;
        RECT 3377.780 2214.460 3377.950 2214.550 ;
      LAYER li1 ;
        RECT 3377.780 2214.145 3377.950 2214.315 ;
        RECT 3383.220 2214.145 3383.390 2214.315 ;
      LAYER li1 ;
        RECT 3377.780 2213.915 3377.950 2214.000 ;
        RECT 3377.780 2210.510 3378.385 2213.915 ;
      LAYER li1 ;
        RECT 3383.220 2213.685 3383.390 2213.855 ;
        RECT 3383.220 2213.225 3383.390 2213.395 ;
        RECT 3383.220 2212.765 3383.390 2212.935 ;
        RECT 3383.220 2212.305 3383.390 2212.475 ;
        RECT 3383.220 2211.845 3383.390 2212.015 ;
        RECT 3383.220 2211.385 3383.390 2211.555 ;
        RECT 3383.220 2210.925 3383.390 2211.095 ;
      LAYER li1 ;
        RECT 3377.780 2210.160 3379.635 2210.510 ;
      LAYER li1 ;
        RECT 3383.220 2210.465 3383.390 2210.635 ;
      LAYER li1 ;
        RECT 3377.780 2208.570 3378.385 2210.160 ;
      LAYER li1 ;
        RECT 3383.220 2210.005 3383.390 2210.175 ;
        RECT 3383.220 2209.545 3383.390 2209.715 ;
        RECT 3383.220 2209.085 3383.390 2209.255 ;
        RECT 3383.220 2208.625 3383.390 2208.795 ;
      LAYER li1 ;
        RECT 3377.780 2208.480 3377.950 2208.570 ;
      LAYER li1 ;
        RECT 3377.780 2208.165 3377.950 2208.335 ;
        RECT 3383.220 2208.165 3383.390 2208.335 ;
      LAYER li1 ;
        RECT 3377.780 2207.935 3377.950 2208.020 ;
        RECT 3377.780 2204.530 3378.385 2207.935 ;
      LAYER li1 ;
        RECT 3383.220 2207.705 3383.390 2207.875 ;
        RECT 3383.220 2207.245 3383.390 2207.415 ;
        RECT 3383.220 2206.785 3383.390 2206.955 ;
        RECT 3383.220 2206.325 3383.390 2206.495 ;
        RECT 3383.220 2205.865 3383.390 2206.035 ;
        RECT 3383.220 2205.405 3383.390 2205.575 ;
        RECT 3383.220 2204.945 3383.390 2205.115 ;
      LAYER li1 ;
        RECT 3377.780 2204.180 3379.635 2204.530 ;
      LAYER li1 ;
        RECT 3383.220 2204.485 3383.390 2204.655 ;
      LAYER li1 ;
        RECT 3377.780 2202.590 3378.385 2204.180 ;
      LAYER li1 ;
        RECT 3383.220 2204.025 3383.390 2204.195 ;
        RECT 3383.220 2203.565 3383.390 2203.735 ;
        RECT 3383.220 2203.105 3383.390 2203.275 ;
        RECT 3383.220 2202.645 3383.390 2202.815 ;
      LAYER li1 ;
        RECT 3377.780 2202.500 3377.950 2202.590 ;
      LAYER li1 ;
        RECT 3377.780 2202.185 3377.950 2202.355 ;
        RECT 3383.220 2202.185 3383.390 2202.355 ;
      LAYER li1 ;
        RECT 3377.780 2201.955 3377.950 2202.040 ;
        RECT 3377.780 2198.550 3378.385 2201.955 ;
      LAYER li1 ;
        RECT 3383.220 2201.725 3383.390 2201.895 ;
        RECT 3383.220 2201.265 3383.390 2201.435 ;
        RECT 3383.220 2200.805 3383.390 2200.975 ;
        RECT 3383.220 2200.345 3383.390 2200.515 ;
        RECT 3383.220 2199.885 3383.390 2200.055 ;
        RECT 3383.220 2199.425 3383.390 2199.595 ;
        RECT 3383.220 2198.965 3383.390 2199.135 ;
      LAYER li1 ;
        RECT 3377.780 2198.200 3379.635 2198.550 ;
      LAYER li1 ;
        RECT 3383.220 2198.505 3383.390 2198.675 ;
      LAYER li1 ;
        RECT 3377.780 2196.610 3378.385 2198.200 ;
      LAYER li1 ;
        RECT 3383.220 2198.045 3383.390 2198.215 ;
        RECT 3383.220 2197.585 3383.390 2197.755 ;
        RECT 3383.220 2197.125 3383.390 2197.295 ;
        RECT 3383.220 2196.665 3383.390 2196.835 ;
      LAYER li1 ;
        RECT 3377.780 2196.520 3377.950 2196.610 ;
      LAYER li1 ;
        RECT 3377.780 2196.205 3377.950 2196.375 ;
        RECT 3383.220 2196.205 3383.390 2196.375 ;
      LAYER mcon ;
        RECT 3377.780 2267.045 3377.950 2267.215 ;
        RECT 3377.780 2266.585 3377.950 2266.755 ;
        RECT 3377.780 2266.125 3377.950 2266.295 ;
        RECT 3377.780 2265.665 3377.950 2265.835 ;
        RECT 3377.780 2265.205 3377.950 2265.375 ;
        RECT 3377.780 2264.745 3377.950 2264.915 ;
        RECT 3377.780 2264.285 3377.950 2264.455 ;
        RECT 3377.780 2263.825 3377.950 2263.995 ;
        RECT 3377.780 2263.365 3377.950 2263.535 ;
        RECT 3377.780 2262.905 3377.950 2263.075 ;
        RECT 3377.780 2262.445 3377.950 2262.615 ;
        RECT 3377.780 2261.065 3377.950 2261.235 ;
        RECT 3377.780 2260.605 3377.950 2260.775 ;
        RECT 3377.780 2260.145 3377.950 2260.315 ;
        RECT 3377.780 2259.685 3377.950 2259.855 ;
        RECT 3377.780 2259.225 3377.950 2259.395 ;
        RECT 3377.780 2258.765 3377.950 2258.935 ;
        RECT 3377.780 2258.305 3377.950 2258.475 ;
        RECT 3377.780 2257.845 3377.950 2258.015 ;
        RECT 3377.780 2257.385 3377.950 2257.555 ;
        RECT 3377.780 2256.925 3377.950 2257.095 ;
        RECT 3377.780 2256.465 3377.950 2256.635 ;
        RECT 3377.780 2255.085 3377.950 2255.255 ;
        RECT 3377.780 2254.625 3377.950 2254.795 ;
        RECT 3377.780 2254.165 3377.950 2254.335 ;
        RECT 3377.780 2253.705 3377.950 2253.875 ;
        RECT 3377.780 2253.245 3377.950 2253.415 ;
        RECT 3377.780 2252.785 3377.950 2252.955 ;
        RECT 3377.780 2252.325 3377.950 2252.495 ;
        RECT 3377.780 2251.865 3377.950 2252.035 ;
        RECT 3377.780 2251.405 3377.950 2251.575 ;
        RECT 3377.780 2250.945 3377.950 2251.115 ;
        RECT 3377.780 2250.485 3377.950 2250.655 ;
        RECT 3377.780 2249.105 3377.950 2249.275 ;
        RECT 3377.780 2248.645 3377.950 2248.815 ;
        RECT 3377.780 2248.185 3377.950 2248.355 ;
        RECT 3377.780 2247.725 3377.950 2247.895 ;
        RECT 3377.780 2247.265 3377.950 2247.435 ;
        RECT 3377.780 2246.805 3377.950 2246.975 ;
        RECT 3377.780 2246.345 3377.950 2246.515 ;
        RECT 3377.780 2245.885 3377.950 2246.055 ;
        RECT 3377.780 2245.425 3377.950 2245.595 ;
        RECT 3377.780 2244.965 3377.950 2245.135 ;
        RECT 3377.780 2244.505 3377.950 2244.675 ;
        RECT 3377.780 2243.125 3377.950 2243.295 ;
        RECT 3377.780 2242.665 3377.950 2242.835 ;
        RECT 3377.780 2242.205 3377.950 2242.375 ;
        RECT 3377.780 2241.745 3377.950 2241.915 ;
        RECT 3377.780 2241.285 3377.950 2241.455 ;
        RECT 3377.780 2240.825 3377.950 2240.995 ;
        RECT 3377.780 2240.365 3377.950 2240.535 ;
        RECT 3377.780 2239.905 3377.950 2240.075 ;
        RECT 3377.780 2239.445 3377.950 2239.615 ;
        RECT 3377.780 2238.985 3377.950 2239.155 ;
        RECT 3377.780 2238.525 3377.950 2238.695 ;
        RECT 3377.780 2237.145 3377.950 2237.315 ;
        RECT 3377.780 2236.685 3377.950 2236.855 ;
        RECT 3377.780 2236.225 3377.950 2236.395 ;
        RECT 3377.780 2235.765 3377.950 2235.935 ;
        RECT 3377.780 2235.305 3377.950 2235.475 ;
        RECT 3377.780 2234.845 3377.950 2235.015 ;
        RECT 3377.780 2234.385 3377.950 2234.555 ;
        RECT 3377.780 2233.925 3377.950 2234.095 ;
        RECT 3377.780 2233.465 3377.950 2233.635 ;
        RECT 3377.780 2233.005 3377.950 2233.175 ;
        RECT 3377.780 2232.545 3377.950 2232.715 ;
        RECT 3377.780 2231.165 3377.950 2231.335 ;
        RECT 3377.780 2230.705 3377.950 2230.875 ;
        RECT 3377.780 2230.245 3377.950 2230.415 ;
        RECT 3377.780 2229.785 3377.950 2229.955 ;
        RECT 3377.780 2229.325 3377.950 2229.495 ;
        RECT 3377.780 2228.865 3377.950 2229.035 ;
        RECT 3377.780 2228.405 3377.950 2228.575 ;
        RECT 3377.780 2227.945 3377.950 2228.115 ;
        RECT 3377.780 2227.485 3377.950 2227.655 ;
        RECT 3377.780 2227.025 3377.950 2227.195 ;
        RECT 3377.780 2226.565 3377.950 2226.735 ;
        RECT 3377.780 2225.185 3377.950 2225.355 ;
        RECT 3377.780 2224.725 3377.950 2224.895 ;
        RECT 3377.780 2224.265 3377.950 2224.435 ;
        RECT 3377.780 2223.805 3377.950 2223.975 ;
        RECT 3377.780 2223.345 3377.950 2223.515 ;
        RECT 3377.780 2222.885 3377.950 2223.055 ;
        RECT 3377.780 2222.425 3377.950 2222.595 ;
        RECT 3377.780 2221.965 3377.950 2222.135 ;
        RECT 3377.780 2221.505 3377.950 2221.675 ;
        RECT 3377.780 2221.045 3377.950 2221.215 ;
        RECT 3377.780 2220.585 3377.950 2220.755 ;
        RECT 3377.780 2219.205 3377.950 2219.375 ;
        RECT 3377.780 2218.745 3377.950 2218.915 ;
        RECT 3377.780 2218.285 3377.950 2218.455 ;
        RECT 3377.780 2217.825 3377.950 2217.995 ;
        RECT 3377.780 2217.365 3377.950 2217.535 ;
        RECT 3377.780 2216.905 3377.950 2217.075 ;
        RECT 3377.780 2216.445 3377.950 2216.615 ;
        RECT 3377.780 2215.985 3377.950 2216.155 ;
        RECT 3377.780 2215.525 3377.950 2215.695 ;
        RECT 3377.780 2215.065 3377.950 2215.235 ;
        RECT 3377.780 2214.605 3377.950 2214.775 ;
        RECT 3377.780 2213.225 3377.950 2213.395 ;
        RECT 3377.780 2212.765 3377.950 2212.935 ;
        RECT 3377.780 2212.305 3377.950 2212.475 ;
        RECT 3377.780 2211.845 3377.950 2212.015 ;
        RECT 3377.780 2211.385 3377.950 2211.555 ;
        RECT 3377.780 2210.925 3377.950 2211.095 ;
        RECT 3377.780 2210.465 3377.950 2210.635 ;
        RECT 3377.780 2210.005 3377.950 2210.175 ;
        RECT 3377.780 2209.545 3377.950 2209.715 ;
        RECT 3377.780 2209.085 3377.950 2209.255 ;
        RECT 3377.780 2208.625 3377.950 2208.795 ;
        RECT 3377.780 2207.245 3377.950 2207.415 ;
        RECT 3377.780 2206.785 3377.950 2206.955 ;
        RECT 3377.780 2206.325 3377.950 2206.495 ;
        RECT 3377.780 2205.865 3377.950 2206.035 ;
        RECT 3377.780 2205.405 3377.950 2205.575 ;
        RECT 3377.780 2204.945 3377.950 2205.115 ;
        RECT 3377.780 2204.485 3377.950 2204.655 ;
        RECT 3377.780 2204.025 3377.950 2204.195 ;
        RECT 3377.780 2203.565 3377.950 2203.735 ;
        RECT 3377.780 2203.105 3377.950 2203.275 ;
        RECT 3377.780 2202.645 3377.950 2202.815 ;
        RECT 3377.780 2201.265 3377.950 2201.435 ;
        RECT 3377.780 2200.805 3377.950 2200.975 ;
        RECT 3377.780 2200.345 3377.950 2200.515 ;
        RECT 3377.780 2199.885 3377.950 2200.055 ;
        RECT 3377.780 2199.425 3377.950 2199.595 ;
        RECT 3377.780 2198.965 3377.950 2199.135 ;
        RECT 3377.780 2198.505 3377.950 2198.675 ;
        RECT 3377.780 2198.045 3377.950 2198.215 ;
        RECT 3377.780 2197.585 3377.950 2197.755 ;
        RECT 3377.780 2197.125 3377.950 2197.295 ;
        RECT 3377.780 2196.665 3377.950 2196.835 ;
      LAYER met1 ;
        RECT 3377.625 2196.060 3378.105 2268.280 ;
        RECT 3383.065 2196.060 3383.545 2268.280 ;
      LAYER via ;
        RECT 3377.690 2234.495 3377.990 2236.280 ;
        RECT 3383.130 2234.495 3383.430 2236.280 ;
      LAYER met2 ;
        RECT 3377.620 2234.455 3378.050 2236.320 ;
        RECT 3383.060 2234.455 3383.490 2236.320 ;
      LAYER via2 ;
        RECT 3377.690 2234.495 3377.990 2236.280 ;
        RECT 3383.130 2234.495 3383.430 2236.280 ;
      LAYER met3 ;
        RECT 3377.620 2234.465 3387.875 2236.315 ;
    END
    PORT
      LAYER li1 ;
        RECT 3377.780 3638.085 3377.950 3638.255 ;
        RECT 3383.220 3638.085 3383.390 3638.255 ;
      LAYER li1 ;
        RECT 3377.780 3637.855 3377.950 3637.940 ;
        RECT 3377.780 3634.450 3378.385 3637.855 ;
      LAYER li1 ;
        RECT 3383.220 3637.625 3383.390 3637.795 ;
        RECT 3383.220 3637.165 3383.390 3637.335 ;
        RECT 3383.220 3636.705 3383.390 3636.875 ;
        RECT 3383.220 3636.245 3383.390 3636.415 ;
        RECT 3383.220 3635.785 3383.390 3635.955 ;
        RECT 3383.220 3635.325 3383.390 3635.495 ;
        RECT 3383.220 3634.865 3383.390 3635.035 ;
      LAYER li1 ;
        RECT 3377.780 3634.100 3379.635 3634.450 ;
      LAYER li1 ;
        RECT 3383.220 3634.405 3383.390 3634.575 ;
      LAYER li1 ;
        RECT 3377.780 3632.510 3378.385 3634.100 ;
      LAYER li1 ;
        RECT 3383.220 3633.945 3383.390 3634.115 ;
        RECT 3383.220 3633.485 3383.390 3633.655 ;
        RECT 3383.220 3633.025 3383.390 3633.195 ;
        RECT 3383.220 3632.565 3383.390 3632.735 ;
      LAYER li1 ;
        RECT 3377.780 3632.420 3377.950 3632.510 ;
      LAYER li1 ;
        RECT 3377.780 3632.105 3377.950 3632.275 ;
        RECT 3383.220 3632.105 3383.390 3632.275 ;
      LAYER li1 ;
        RECT 3377.780 3631.875 3377.950 3631.960 ;
        RECT 3377.780 3628.470 3378.385 3631.875 ;
      LAYER li1 ;
        RECT 3383.220 3631.645 3383.390 3631.815 ;
        RECT 3383.220 3631.185 3383.390 3631.355 ;
        RECT 3383.220 3630.725 3383.390 3630.895 ;
        RECT 3383.220 3630.265 3383.390 3630.435 ;
        RECT 3383.220 3629.805 3383.390 3629.975 ;
        RECT 3383.220 3629.345 3383.390 3629.515 ;
        RECT 3383.220 3628.885 3383.390 3629.055 ;
      LAYER li1 ;
        RECT 3377.780 3628.120 3379.635 3628.470 ;
      LAYER li1 ;
        RECT 3383.220 3628.425 3383.390 3628.595 ;
      LAYER li1 ;
        RECT 3377.780 3626.530 3378.385 3628.120 ;
      LAYER li1 ;
        RECT 3383.220 3627.965 3383.390 3628.135 ;
        RECT 3383.220 3627.505 3383.390 3627.675 ;
        RECT 3383.220 3627.045 3383.390 3627.215 ;
        RECT 3383.220 3626.585 3383.390 3626.755 ;
      LAYER li1 ;
        RECT 3377.780 3626.440 3377.950 3626.530 ;
      LAYER li1 ;
        RECT 3377.780 3626.125 3377.950 3626.295 ;
        RECT 3383.220 3626.125 3383.390 3626.295 ;
      LAYER li1 ;
        RECT 3377.780 3625.895 3377.950 3625.980 ;
        RECT 3377.780 3622.490 3378.385 3625.895 ;
      LAYER li1 ;
        RECT 3383.220 3625.665 3383.390 3625.835 ;
        RECT 3383.220 3625.205 3383.390 3625.375 ;
        RECT 3383.220 3624.745 3383.390 3624.915 ;
        RECT 3383.220 3624.285 3383.390 3624.455 ;
        RECT 3383.220 3623.825 3383.390 3623.995 ;
        RECT 3383.220 3623.365 3383.390 3623.535 ;
        RECT 3383.220 3622.905 3383.390 3623.075 ;
      LAYER li1 ;
        RECT 3377.780 3622.140 3379.635 3622.490 ;
      LAYER li1 ;
        RECT 3383.220 3622.445 3383.390 3622.615 ;
      LAYER li1 ;
        RECT 3377.780 3620.550 3378.385 3622.140 ;
      LAYER li1 ;
        RECT 3383.220 3621.985 3383.390 3622.155 ;
        RECT 3383.220 3621.525 3383.390 3621.695 ;
        RECT 3383.220 3621.065 3383.390 3621.235 ;
        RECT 3383.220 3620.605 3383.390 3620.775 ;
      LAYER li1 ;
        RECT 3377.780 3620.460 3377.950 3620.550 ;
      LAYER li1 ;
        RECT 3377.780 3620.145 3377.950 3620.315 ;
        RECT 3383.220 3620.145 3383.390 3620.315 ;
      LAYER li1 ;
        RECT 3377.780 3619.915 3377.950 3620.000 ;
        RECT 3377.780 3616.510 3378.385 3619.915 ;
      LAYER li1 ;
        RECT 3383.220 3619.685 3383.390 3619.855 ;
        RECT 3383.220 3619.225 3383.390 3619.395 ;
        RECT 3383.220 3618.765 3383.390 3618.935 ;
        RECT 3383.220 3618.305 3383.390 3618.475 ;
        RECT 3383.220 3617.845 3383.390 3618.015 ;
        RECT 3383.220 3617.385 3383.390 3617.555 ;
        RECT 3383.220 3616.925 3383.390 3617.095 ;
      LAYER li1 ;
        RECT 3377.780 3616.160 3379.635 3616.510 ;
      LAYER li1 ;
        RECT 3383.220 3616.465 3383.390 3616.635 ;
      LAYER li1 ;
        RECT 3377.780 3614.570 3378.385 3616.160 ;
      LAYER li1 ;
        RECT 3383.220 3616.005 3383.390 3616.175 ;
        RECT 3383.220 3615.545 3383.390 3615.715 ;
        RECT 3383.220 3615.085 3383.390 3615.255 ;
        RECT 3383.220 3614.625 3383.390 3614.795 ;
      LAYER li1 ;
        RECT 3377.780 3614.480 3377.950 3614.570 ;
      LAYER li1 ;
        RECT 3377.780 3614.165 3377.950 3614.335 ;
        RECT 3383.220 3614.165 3383.390 3614.335 ;
      LAYER li1 ;
        RECT 3377.780 3613.935 3377.950 3614.020 ;
        RECT 3377.780 3610.530 3378.385 3613.935 ;
      LAYER li1 ;
        RECT 3383.220 3613.705 3383.390 3613.875 ;
        RECT 3383.220 3613.245 3383.390 3613.415 ;
        RECT 3383.220 3612.785 3383.390 3612.955 ;
        RECT 3383.220 3612.325 3383.390 3612.495 ;
        RECT 3383.220 3611.865 3383.390 3612.035 ;
        RECT 3383.220 3611.405 3383.390 3611.575 ;
        RECT 3383.220 3610.945 3383.390 3611.115 ;
      LAYER li1 ;
        RECT 3377.780 3610.180 3379.635 3610.530 ;
      LAYER li1 ;
        RECT 3383.220 3610.485 3383.390 3610.655 ;
      LAYER li1 ;
        RECT 3377.780 3608.590 3378.385 3610.180 ;
      LAYER li1 ;
        RECT 3383.220 3610.025 3383.390 3610.195 ;
        RECT 3383.220 3609.565 3383.390 3609.735 ;
        RECT 3383.220 3609.105 3383.390 3609.275 ;
        RECT 3383.220 3608.645 3383.390 3608.815 ;
      LAYER li1 ;
        RECT 3377.780 3608.500 3377.950 3608.590 ;
      LAYER li1 ;
        RECT 3377.780 3608.185 3377.950 3608.355 ;
        RECT 3383.220 3608.185 3383.390 3608.355 ;
      LAYER li1 ;
        RECT 3377.780 3607.955 3377.950 3608.040 ;
        RECT 3377.780 3604.550 3378.385 3607.955 ;
      LAYER li1 ;
        RECT 3383.220 3607.725 3383.390 3607.895 ;
        RECT 3383.220 3607.265 3383.390 3607.435 ;
        RECT 3383.220 3606.805 3383.390 3606.975 ;
        RECT 3383.220 3606.345 3383.390 3606.515 ;
        RECT 3383.220 3605.885 3383.390 3606.055 ;
        RECT 3383.220 3605.425 3383.390 3605.595 ;
        RECT 3383.220 3604.965 3383.390 3605.135 ;
      LAYER li1 ;
        RECT 3377.780 3604.200 3379.635 3604.550 ;
      LAYER li1 ;
        RECT 3383.220 3604.505 3383.390 3604.675 ;
      LAYER li1 ;
        RECT 3377.780 3602.610 3378.385 3604.200 ;
      LAYER li1 ;
        RECT 3383.220 3604.045 3383.390 3604.215 ;
        RECT 3383.220 3603.585 3383.390 3603.755 ;
        RECT 3383.220 3603.125 3383.390 3603.295 ;
        RECT 3383.220 3602.665 3383.390 3602.835 ;
      LAYER li1 ;
        RECT 3377.780 3602.520 3377.950 3602.610 ;
      LAYER li1 ;
        RECT 3377.780 3602.205 3377.950 3602.375 ;
        RECT 3383.220 3602.205 3383.390 3602.375 ;
      LAYER mcon ;
        RECT 3377.780 3637.165 3377.950 3637.335 ;
        RECT 3377.780 3636.705 3377.950 3636.875 ;
        RECT 3377.780 3636.245 3377.950 3636.415 ;
        RECT 3377.780 3635.785 3377.950 3635.955 ;
        RECT 3377.780 3635.325 3377.950 3635.495 ;
        RECT 3377.780 3634.865 3377.950 3635.035 ;
        RECT 3377.780 3634.405 3377.950 3634.575 ;
        RECT 3377.780 3633.945 3377.950 3634.115 ;
        RECT 3377.780 3633.485 3377.950 3633.655 ;
        RECT 3377.780 3633.025 3377.950 3633.195 ;
        RECT 3377.780 3632.565 3377.950 3632.735 ;
        RECT 3377.780 3631.185 3377.950 3631.355 ;
        RECT 3377.780 3630.725 3377.950 3630.895 ;
        RECT 3377.780 3630.265 3377.950 3630.435 ;
        RECT 3377.780 3629.805 3377.950 3629.975 ;
        RECT 3377.780 3629.345 3377.950 3629.515 ;
        RECT 3377.780 3628.885 3377.950 3629.055 ;
        RECT 3377.780 3628.425 3377.950 3628.595 ;
        RECT 3377.780 3627.965 3377.950 3628.135 ;
        RECT 3377.780 3627.505 3377.950 3627.675 ;
        RECT 3377.780 3627.045 3377.950 3627.215 ;
        RECT 3377.780 3626.585 3377.950 3626.755 ;
        RECT 3377.780 3625.205 3377.950 3625.375 ;
        RECT 3377.780 3624.745 3377.950 3624.915 ;
        RECT 3377.780 3624.285 3377.950 3624.455 ;
        RECT 3377.780 3623.825 3377.950 3623.995 ;
        RECT 3377.780 3623.365 3377.950 3623.535 ;
        RECT 3377.780 3622.905 3377.950 3623.075 ;
        RECT 3377.780 3622.445 3377.950 3622.615 ;
        RECT 3377.780 3621.985 3377.950 3622.155 ;
        RECT 3377.780 3621.525 3377.950 3621.695 ;
        RECT 3377.780 3621.065 3377.950 3621.235 ;
        RECT 3377.780 3620.605 3377.950 3620.775 ;
        RECT 3377.780 3619.225 3377.950 3619.395 ;
        RECT 3377.780 3618.765 3377.950 3618.935 ;
        RECT 3377.780 3618.305 3377.950 3618.475 ;
        RECT 3377.780 3617.845 3377.950 3618.015 ;
        RECT 3377.780 3617.385 3377.950 3617.555 ;
        RECT 3377.780 3616.925 3377.950 3617.095 ;
        RECT 3377.780 3616.465 3377.950 3616.635 ;
        RECT 3377.780 3616.005 3377.950 3616.175 ;
        RECT 3377.780 3615.545 3377.950 3615.715 ;
        RECT 3377.780 3615.085 3377.950 3615.255 ;
        RECT 3377.780 3614.625 3377.950 3614.795 ;
        RECT 3377.780 3613.245 3377.950 3613.415 ;
        RECT 3377.780 3612.785 3377.950 3612.955 ;
        RECT 3377.780 3612.325 3377.950 3612.495 ;
        RECT 3377.780 3611.865 3377.950 3612.035 ;
        RECT 3377.780 3611.405 3377.950 3611.575 ;
        RECT 3377.780 3610.945 3377.950 3611.115 ;
        RECT 3377.780 3610.485 3377.950 3610.655 ;
        RECT 3377.780 3610.025 3377.950 3610.195 ;
        RECT 3377.780 3609.565 3377.950 3609.735 ;
        RECT 3377.780 3609.105 3377.950 3609.275 ;
        RECT 3377.780 3608.645 3377.950 3608.815 ;
        RECT 3377.780 3607.265 3377.950 3607.435 ;
        RECT 3377.780 3606.805 3377.950 3606.975 ;
        RECT 3377.780 3606.345 3377.950 3606.515 ;
        RECT 3377.780 3605.885 3377.950 3606.055 ;
        RECT 3377.780 3605.425 3377.950 3605.595 ;
        RECT 3377.780 3604.965 3377.950 3605.135 ;
        RECT 3377.780 3604.505 3377.950 3604.675 ;
        RECT 3377.780 3604.045 3377.950 3604.215 ;
        RECT 3377.780 3603.585 3377.950 3603.755 ;
        RECT 3377.780 3603.125 3377.950 3603.295 ;
        RECT 3377.780 3602.665 3377.950 3602.835 ;
      LAYER met1 ;
        RECT 3377.625 3602.060 3378.105 3638.400 ;
        RECT 3383.065 3602.060 3383.545 3638.400 ;
      LAYER via ;
        RECT 3377.730 3616.500 3378.030 3618.285 ;
        RECT 3383.170 3616.500 3383.470 3618.285 ;
      LAYER met2 ;
        RECT 3377.660 3616.460 3378.090 3618.325 ;
        RECT 3383.100 3616.460 3383.530 3618.325 ;
      LAYER via2 ;
        RECT 3377.730 3616.500 3378.030 3618.285 ;
        RECT 3383.170 3616.500 3383.470 3618.285 ;
      LAYER met3 ;
        RECT 3377.660 3616.470 3387.915 3618.320 ;
    END
    PORT
      LAYER li1 ;
        RECT 669.145 219.760 669.315 219.930 ;
      LAYER li1 ;
        RECT 669.460 219.760 674.980 219.930 ;
      LAYER li1 ;
        RECT 675.125 219.760 675.295 219.930 ;
      LAYER li1 ;
        RECT 675.440 219.760 680.960 219.930 ;
      LAYER li1 ;
        RECT 681.105 219.760 681.275 219.930 ;
      LAYER li1 ;
        RECT 681.420 219.760 686.940 219.930 ;
      LAYER li1 ;
        RECT 687.085 219.760 687.255 219.930 ;
      LAYER li1 ;
        RECT 687.400 219.760 692.920 219.930 ;
      LAYER li1 ;
        RECT 693.065 219.760 693.235 219.930 ;
      LAYER li1 ;
        RECT 693.380 219.760 698.900 219.930 ;
      LAYER li1 ;
        RECT 699.045 219.760 699.215 219.930 ;
      LAYER li1 ;
        RECT 699.360 219.760 704.880 219.930 ;
      LAYER li1 ;
        RECT 705.025 219.760 705.195 219.930 ;
      LAYER li1 ;
        RECT 705.340 219.760 710.860 219.930 ;
      LAYER li1 ;
        RECT 711.005 219.760 711.175 219.930 ;
      LAYER li1 ;
        RECT 711.320 219.760 716.840 219.930 ;
      LAYER li1 ;
        RECT 716.985 219.760 717.155 219.930 ;
      LAYER li1 ;
        RECT 717.300 219.760 722.820 219.930 ;
      LAYER li1 ;
        RECT 722.965 219.760 723.135 219.930 ;
      LAYER li1 ;
        RECT 723.280 219.760 728.800 219.930 ;
      LAYER li1 ;
        RECT 728.945 219.760 729.115 219.930 ;
      LAYER li1 ;
        RECT 729.260 219.760 734.780 219.930 ;
      LAYER li1 ;
        RECT 734.925 219.760 735.095 219.930 ;
      LAYER li1 ;
        RECT 735.240 219.760 740.760 219.930 ;
      LAYER li1 ;
        RECT 740.905 219.760 741.075 219.930 ;
      LAYER li1 ;
        RECT 741.220 219.760 746.740 219.930 ;
      LAYER li1 ;
        RECT 746.885 219.760 747.055 219.930 ;
      LAYER li1 ;
        RECT 747.200 219.760 752.720 219.930 ;
      LAYER li1 ;
        RECT 752.865 219.760 753.035 219.930 ;
      LAYER li1 ;
        RECT 753.180 219.760 758.700 219.930 ;
      LAYER li1 ;
        RECT 758.845 219.760 759.015 219.930 ;
      LAYER li1 ;
        RECT 759.160 219.760 764.680 219.930 ;
      LAYER li1 ;
        RECT 764.825 219.760 764.995 219.930 ;
      LAYER li1 ;
        RECT 765.140 219.760 770.660 219.930 ;
      LAYER li1 ;
        RECT 770.805 219.760 770.975 219.930 ;
      LAYER li1 ;
        RECT 771.120 219.760 776.640 219.930 ;
      LAYER li1 ;
        RECT 776.785 219.760 776.955 219.930 ;
      LAYER li1 ;
        RECT 777.100 219.760 782.620 219.930 ;
      LAYER li1 ;
        RECT 782.765 219.760 782.935 219.930 ;
      LAYER li1 ;
        RECT 783.080 219.760 788.600 219.930 ;
      LAYER li1 ;
        RECT 788.745 219.760 788.915 219.930 ;
      LAYER li1 ;
        RECT 789.060 219.760 794.580 219.930 ;
      LAYER li1 ;
        RECT 794.725 219.760 794.895 219.930 ;
      LAYER li1 ;
        RECT 669.545 219.325 674.890 219.760 ;
        RECT 675.525 219.325 680.870 219.760 ;
        RECT 681.505 219.325 686.850 219.760 ;
        RECT 687.485 219.325 692.830 219.760 ;
        RECT 693.465 219.325 698.810 219.760 ;
        RECT 699.445 219.325 704.790 219.760 ;
        RECT 705.425 219.325 710.770 219.760 ;
        RECT 711.405 219.325 716.750 219.760 ;
        RECT 717.385 219.325 722.730 219.760 ;
        RECT 723.365 219.325 728.710 219.760 ;
        RECT 729.345 219.325 734.690 219.760 ;
        RECT 735.325 219.325 740.670 219.760 ;
        RECT 741.305 219.325 746.650 219.760 ;
        RECT 747.285 219.325 752.630 219.760 ;
        RECT 753.265 219.325 758.610 219.760 ;
        RECT 759.245 219.325 764.590 219.760 ;
        RECT 765.225 219.325 770.570 219.760 ;
        RECT 771.205 219.325 776.550 219.760 ;
        RECT 777.185 219.325 782.530 219.760 ;
        RECT 783.165 219.325 788.510 219.760 ;
        RECT 789.145 219.325 794.490 219.760 ;
        RECT 672.950 218.075 673.300 219.325 ;
        RECT 678.930 218.075 679.280 219.325 ;
        RECT 684.910 218.075 685.260 219.325 ;
        RECT 690.890 218.075 691.240 219.325 ;
        RECT 696.870 218.075 697.220 219.325 ;
        RECT 702.850 218.075 703.200 219.325 ;
        RECT 708.830 218.075 709.180 219.325 ;
        RECT 714.810 218.075 715.160 219.325 ;
        RECT 720.790 218.075 721.140 219.325 ;
        RECT 726.770 218.075 727.120 219.325 ;
        RECT 732.750 218.075 733.100 219.325 ;
        RECT 738.730 218.075 739.080 219.325 ;
        RECT 744.710 218.075 745.060 219.325 ;
        RECT 750.690 218.075 751.040 219.325 ;
        RECT 756.670 218.075 757.020 219.325 ;
        RECT 762.650 218.075 763.000 219.325 ;
        RECT 768.630 218.075 768.980 219.325 ;
        RECT 774.610 218.075 774.960 219.325 ;
        RECT 780.590 218.075 780.940 219.325 ;
        RECT 786.570 218.075 786.920 219.325 ;
        RECT 792.550 218.075 792.900 219.325 ;
      LAYER li1 ;
        RECT 669.145 214.320 669.315 214.490 ;
        RECT 669.605 214.320 669.775 214.490 ;
        RECT 670.065 214.320 670.235 214.490 ;
        RECT 670.525 214.320 670.695 214.490 ;
        RECT 670.985 214.320 671.155 214.490 ;
        RECT 671.445 214.320 671.615 214.490 ;
        RECT 671.905 214.320 672.075 214.490 ;
        RECT 672.365 214.320 672.535 214.490 ;
        RECT 672.825 214.320 672.995 214.490 ;
        RECT 673.285 214.320 673.455 214.490 ;
        RECT 673.745 214.320 673.915 214.490 ;
        RECT 674.205 214.320 674.375 214.490 ;
        RECT 674.665 214.320 674.835 214.490 ;
        RECT 675.125 214.320 675.295 214.490 ;
        RECT 675.585 214.320 675.755 214.490 ;
        RECT 676.045 214.320 676.215 214.490 ;
        RECT 676.505 214.320 676.675 214.490 ;
        RECT 676.965 214.320 677.135 214.490 ;
        RECT 677.425 214.320 677.595 214.490 ;
        RECT 677.885 214.320 678.055 214.490 ;
        RECT 678.345 214.320 678.515 214.490 ;
        RECT 678.805 214.320 678.975 214.490 ;
        RECT 679.265 214.320 679.435 214.490 ;
        RECT 679.725 214.320 679.895 214.490 ;
        RECT 680.185 214.320 680.355 214.490 ;
        RECT 680.645 214.320 680.815 214.490 ;
        RECT 681.105 214.320 681.275 214.490 ;
        RECT 681.565 214.320 681.735 214.490 ;
        RECT 682.025 214.320 682.195 214.490 ;
        RECT 682.485 214.320 682.655 214.490 ;
        RECT 682.945 214.320 683.115 214.490 ;
        RECT 683.405 214.320 683.575 214.490 ;
        RECT 683.865 214.320 684.035 214.490 ;
        RECT 684.325 214.320 684.495 214.490 ;
        RECT 684.785 214.320 684.955 214.490 ;
        RECT 685.245 214.320 685.415 214.490 ;
        RECT 685.705 214.320 685.875 214.490 ;
        RECT 686.165 214.320 686.335 214.490 ;
        RECT 686.625 214.320 686.795 214.490 ;
        RECT 687.085 214.320 687.255 214.490 ;
        RECT 687.545 214.320 687.715 214.490 ;
        RECT 688.005 214.320 688.175 214.490 ;
        RECT 688.465 214.320 688.635 214.490 ;
        RECT 688.925 214.320 689.095 214.490 ;
        RECT 689.385 214.320 689.555 214.490 ;
        RECT 689.845 214.320 690.015 214.490 ;
        RECT 690.305 214.320 690.475 214.490 ;
        RECT 690.765 214.320 690.935 214.490 ;
        RECT 691.225 214.320 691.395 214.490 ;
        RECT 691.685 214.320 691.855 214.490 ;
        RECT 692.145 214.320 692.315 214.490 ;
        RECT 692.605 214.320 692.775 214.490 ;
        RECT 693.065 214.320 693.235 214.490 ;
        RECT 693.525 214.320 693.695 214.490 ;
        RECT 693.985 214.320 694.155 214.490 ;
        RECT 694.445 214.320 694.615 214.490 ;
        RECT 694.905 214.320 695.075 214.490 ;
        RECT 695.365 214.320 695.535 214.490 ;
        RECT 695.825 214.320 695.995 214.490 ;
        RECT 696.285 214.320 696.455 214.490 ;
        RECT 696.745 214.320 696.915 214.490 ;
        RECT 697.205 214.320 697.375 214.490 ;
        RECT 697.665 214.320 697.835 214.490 ;
        RECT 698.125 214.320 698.295 214.490 ;
        RECT 698.585 214.320 698.755 214.490 ;
        RECT 699.045 214.320 699.215 214.490 ;
        RECT 699.505 214.320 699.675 214.490 ;
        RECT 699.965 214.320 700.135 214.490 ;
        RECT 700.425 214.320 700.595 214.490 ;
        RECT 700.885 214.320 701.055 214.490 ;
        RECT 701.345 214.320 701.515 214.490 ;
        RECT 701.805 214.320 701.975 214.490 ;
        RECT 702.265 214.320 702.435 214.490 ;
        RECT 702.725 214.320 702.895 214.490 ;
        RECT 703.185 214.320 703.355 214.490 ;
        RECT 703.645 214.320 703.815 214.490 ;
        RECT 704.105 214.320 704.275 214.490 ;
        RECT 704.565 214.320 704.735 214.490 ;
        RECT 705.025 214.320 705.195 214.490 ;
        RECT 705.485 214.320 705.655 214.490 ;
        RECT 705.945 214.320 706.115 214.490 ;
        RECT 706.405 214.320 706.575 214.490 ;
        RECT 706.865 214.320 707.035 214.490 ;
        RECT 707.325 214.320 707.495 214.490 ;
        RECT 707.785 214.320 707.955 214.490 ;
        RECT 708.245 214.320 708.415 214.490 ;
        RECT 708.705 214.320 708.875 214.490 ;
        RECT 709.165 214.320 709.335 214.490 ;
        RECT 709.625 214.320 709.795 214.490 ;
        RECT 710.085 214.320 710.255 214.490 ;
        RECT 710.545 214.320 710.715 214.490 ;
        RECT 711.005 214.320 711.175 214.490 ;
        RECT 711.465 214.320 711.635 214.490 ;
        RECT 711.925 214.320 712.095 214.490 ;
        RECT 712.385 214.320 712.555 214.490 ;
        RECT 712.845 214.320 713.015 214.490 ;
        RECT 713.305 214.320 713.475 214.490 ;
        RECT 713.765 214.320 713.935 214.490 ;
        RECT 714.225 214.320 714.395 214.490 ;
        RECT 714.685 214.320 714.855 214.490 ;
        RECT 715.145 214.320 715.315 214.490 ;
        RECT 715.605 214.320 715.775 214.490 ;
        RECT 716.065 214.320 716.235 214.490 ;
        RECT 716.525 214.320 716.695 214.490 ;
        RECT 716.985 214.320 717.155 214.490 ;
        RECT 717.445 214.320 717.615 214.490 ;
        RECT 717.905 214.320 718.075 214.490 ;
        RECT 718.365 214.320 718.535 214.490 ;
        RECT 718.825 214.320 718.995 214.490 ;
        RECT 719.285 214.320 719.455 214.490 ;
        RECT 719.745 214.320 719.915 214.490 ;
        RECT 720.205 214.320 720.375 214.490 ;
        RECT 720.665 214.320 720.835 214.490 ;
        RECT 721.125 214.320 721.295 214.490 ;
        RECT 721.585 214.320 721.755 214.490 ;
        RECT 722.045 214.320 722.215 214.490 ;
        RECT 722.505 214.320 722.675 214.490 ;
        RECT 722.965 214.320 723.135 214.490 ;
        RECT 723.425 214.320 723.595 214.490 ;
        RECT 723.885 214.320 724.055 214.490 ;
        RECT 724.345 214.320 724.515 214.490 ;
        RECT 724.805 214.320 724.975 214.490 ;
        RECT 725.265 214.320 725.435 214.490 ;
        RECT 725.725 214.320 725.895 214.490 ;
        RECT 726.185 214.320 726.355 214.490 ;
        RECT 726.645 214.320 726.815 214.490 ;
        RECT 727.105 214.320 727.275 214.490 ;
        RECT 727.565 214.320 727.735 214.490 ;
        RECT 728.025 214.320 728.195 214.490 ;
        RECT 728.485 214.320 728.655 214.490 ;
        RECT 728.945 214.320 729.115 214.490 ;
        RECT 729.405 214.320 729.575 214.490 ;
        RECT 729.865 214.320 730.035 214.490 ;
        RECT 730.325 214.320 730.495 214.490 ;
        RECT 730.785 214.320 730.955 214.490 ;
        RECT 731.245 214.320 731.415 214.490 ;
        RECT 731.705 214.320 731.875 214.490 ;
        RECT 732.165 214.320 732.335 214.490 ;
        RECT 732.625 214.320 732.795 214.490 ;
        RECT 733.085 214.320 733.255 214.490 ;
        RECT 733.545 214.320 733.715 214.490 ;
        RECT 734.005 214.320 734.175 214.490 ;
        RECT 734.465 214.320 734.635 214.490 ;
        RECT 734.925 214.320 735.095 214.490 ;
        RECT 735.385 214.320 735.555 214.490 ;
        RECT 735.845 214.320 736.015 214.490 ;
        RECT 736.305 214.320 736.475 214.490 ;
        RECT 736.765 214.320 736.935 214.490 ;
        RECT 737.225 214.320 737.395 214.490 ;
        RECT 737.685 214.320 737.855 214.490 ;
        RECT 738.145 214.320 738.315 214.490 ;
        RECT 738.605 214.320 738.775 214.490 ;
        RECT 739.065 214.320 739.235 214.490 ;
        RECT 739.525 214.320 739.695 214.490 ;
        RECT 739.985 214.320 740.155 214.490 ;
        RECT 740.445 214.320 740.615 214.490 ;
        RECT 740.905 214.320 741.075 214.490 ;
        RECT 741.365 214.320 741.535 214.490 ;
        RECT 741.825 214.320 741.995 214.490 ;
        RECT 742.285 214.320 742.455 214.490 ;
        RECT 742.745 214.320 742.915 214.490 ;
        RECT 743.205 214.320 743.375 214.490 ;
        RECT 743.665 214.320 743.835 214.490 ;
        RECT 744.125 214.320 744.295 214.490 ;
        RECT 744.585 214.320 744.755 214.490 ;
        RECT 745.045 214.320 745.215 214.490 ;
        RECT 745.505 214.320 745.675 214.490 ;
        RECT 745.965 214.320 746.135 214.490 ;
        RECT 746.425 214.320 746.595 214.490 ;
        RECT 746.885 214.320 747.055 214.490 ;
        RECT 747.345 214.320 747.515 214.490 ;
        RECT 747.805 214.320 747.975 214.490 ;
        RECT 748.265 214.320 748.435 214.490 ;
        RECT 748.725 214.320 748.895 214.490 ;
        RECT 749.185 214.320 749.355 214.490 ;
        RECT 749.645 214.320 749.815 214.490 ;
        RECT 750.105 214.320 750.275 214.490 ;
        RECT 750.565 214.320 750.735 214.490 ;
        RECT 751.025 214.320 751.195 214.490 ;
        RECT 751.485 214.320 751.655 214.490 ;
        RECT 751.945 214.320 752.115 214.490 ;
        RECT 752.405 214.320 752.575 214.490 ;
        RECT 752.865 214.320 753.035 214.490 ;
        RECT 753.325 214.320 753.495 214.490 ;
        RECT 753.785 214.320 753.955 214.490 ;
        RECT 754.245 214.320 754.415 214.490 ;
        RECT 754.705 214.320 754.875 214.490 ;
        RECT 755.165 214.320 755.335 214.490 ;
        RECT 755.625 214.320 755.795 214.490 ;
        RECT 756.085 214.320 756.255 214.490 ;
        RECT 756.545 214.320 756.715 214.490 ;
        RECT 757.005 214.320 757.175 214.490 ;
        RECT 757.465 214.320 757.635 214.490 ;
        RECT 757.925 214.320 758.095 214.490 ;
        RECT 758.385 214.320 758.555 214.490 ;
        RECT 758.845 214.320 759.015 214.490 ;
        RECT 759.305 214.320 759.475 214.490 ;
        RECT 759.765 214.320 759.935 214.490 ;
        RECT 760.225 214.320 760.395 214.490 ;
        RECT 760.685 214.320 760.855 214.490 ;
        RECT 761.145 214.320 761.315 214.490 ;
        RECT 761.605 214.320 761.775 214.490 ;
        RECT 762.065 214.320 762.235 214.490 ;
        RECT 762.525 214.320 762.695 214.490 ;
        RECT 762.985 214.320 763.155 214.490 ;
        RECT 763.445 214.320 763.615 214.490 ;
        RECT 763.905 214.320 764.075 214.490 ;
        RECT 764.365 214.320 764.535 214.490 ;
        RECT 764.825 214.320 764.995 214.490 ;
        RECT 765.285 214.320 765.455 214.490 ;
        RECT 765.745 214.320 765.915 214.490 ;
        RECT 766.205 214.320 766.375 214.490 ;
        RECT 766.665 214.320 766.835 214.490 ;
        RECT 767.125 214.320 767.295 214.490 ;
        RECT 767.585 214.320 767.755 214.490 ;
        RECT 768.045 214.320 768.215 214.490 ;
        RECT 768.505 214.320 768.675 214.490 ;
        RECT 768.965 214.320 769.135 214.490 ;
        RECT 769.425 214.320 769.595 214.490 ;
        RECT 769.885 214.320 770.055 214.490 ;
        RECT 770.345 214.320 770.515 214.490 ;
        RECT 770.805 214.320 770.975 214.490 ;
        RECT 771.265 214.320 771.435 214.490 ;
        RECT 771.725 214.320 771.895 214.490 ;
        RECT 772.185 214.320 772.355 214.490 ;
        RECT 772.645 214.320 772.815 214.490 ;
        RECT 773.105 214.320 773.275 214.490 ;
        RECT 773.565 214.320 773.735 214.490 ;
        RECT 774.025 214.320 774.195 214.490 ;
        RECT 774.485 214.320 774.655 214.490 ;
        RECT 774.945 214.320 775.115 214.490 ;
        RECT 775.405 214.320 775.575 214.490 ;
        RECT 775.865 214.320 776.035 214.490 ;
        RECT 776.325 214.320 776.495 214.490 ;
        RECT 776.785 214.320 776.955 214.490 ;
        RECT 777.245 214.320 777.415 214.490 ;
        RECT 777.705 214.320 777.875 214.490 ;
        RECT 778.165 214.320 778.335 214.490 ;
        RECT 778.625 214.320 778.795 214.490 ;
        RECT 779.085 214.320 779.255 214.490 ;
        RECT 779.545 214.320 779.715 214.490 ;
        RECT 780.005 214.320 780.175 214.490 ;
        RECT 780.465 214.320 780.635 214.490 ;
        RECT 780.925 214.320 781.095 214.490 ;
        RECT 781.385 214.320 781.555 214.490 ;
        RECT 781.845 214.320 782.015 214.490 ;
        RECT 782.305 214.320 782.475 214.490 ;
        RECT 782.765 214.320 782.935 214.490 ;
        RECT 783.225 214.320 783.395 214.490 ;
        RECT 783.685 214.320 783.855 214.490 ;
        RECT 784.145 214.320 784.315 214.490 ;
        RECT 784.605 214.320 784.775 214.490 ;
        RECT 785.065 214.320 785.235 214.490 ;
        RECT 785.525 214.320 785.695 214.490 ;
        RECT 785.985 214.320 786.155 214.490 ;
        RECT 786.445 214.320 786.615 214.490 ;
        RECT 786.905 214.320 787.075 214.490 ;
        RECT 787.365 214.320 787.535 214.490 ;
        RECT 787.825 214.320 787.995 214.490 ;
        RECT 788.285 214.320 788.455 214.490 ;
        RECT 788.745 214.320 788.915 214.490 ;
        RECT 789.205 214.320 789.375 214.490 ;
        RECT 789.665 214.320 789.835 214.490 ;
        RECT 790.125 214.320 790.295 214.490 ;
        RECT 790.585 214.320 790.755 214.490 ;
        RECT 791.045 214.320 791.215 214.490 ;
        RECT 791.505 214.320 791.675 214.490 ;
        RECT 791.965 214.320 792.135 214.490 ;
        RECT 792.425 214.320 792.595 214.490 ;
        RECT 792.885 214.320 793.055 214.490 ;
        RECT 793.345 214.320 793.515 214.490 ;
        RECT 793.805 214.320 793.975 214.490 ;
        RECT 794.265 214.320 794.435 214.490 ;
        RECT 794.725 214.320 794.895 214.490 ;
      LAYER mcon ;
        RECT 670.065 219.760 670.235 219.930 ;
        RECT 670.525 219.760 670.695 219.930 ;
        RECT 670.985 219.760 671.155 219.930 ;
        RECT 671.445 219.760 671.615 219.930 ;
        RECT 671.905 219.760 672.075 219.930 ;
        RECT 672.365 219.760 672.535 219.930 ;
        RECT 672.825 219.760 672.995 219.930 ;
        RECT 673.285 219.760 673.455 219.930 ;
        RECT 673.745 219.760 673.915 219.930 ;
        RECT 674.205 219.760 674.375 219.930 ;
        RECT 674.665 219.760 674.835 219.930 ;
        RECT 676.045 219.760 676.215 219.930 ;
        RECT 676.505 219.760 676.675 219.930 ;
        RECT 676.965 219.760 677.135 219.930 ;
        RECT 677.425 219.760 677.595 219.930 ;
        RECT 677.885 219.760 678.055 219.930 ;
        RECT 678.345 219.760 678.515 219.930 ;
        RECT 678.805 219.760 678.975 219.930 ;
        RECT 679.265 219.760 679.435 219.930 ;
        RECT 679.725 219.760 679.895 219.930 ;
        RECT 680.185 219.760 680.355 219.930 ;
        RECT 680.645 219.760 680.815 219.930 ;
        RECT 682.025 219.760 682.195 219.930 ;
        RECT 682.485 219.760 682.655 219.930 ;
        RECT 682.945 219.760 683.115 219.930 ;
        RECT 683.405 219.760 683.575 219.930 ;
        RECT 683.865 219.760 684.035 219.930 ;
        RECT 684.325 219.760 684.495 219.930 ;
        RECT 684.785 219.760 684.955 219.930 ;
        RECT 685.245 219.760 685.415 219.930 ;
        RECT 685.705 219.760 685.875 219.930 ;
        RECT 686.165 219.760 686.335 219.930 ;
        RECT 686.625 219.760 686.795 219.930 ;
        RECT 688.005 219.760 688.175 219.930 ;
        RECT 688.465 219.760 688.635 219.930 ;
        RECT 688.925 219.760 689.095 219.930 ;
        RECT 689.385 219.760 689.555 219.930 ;
        RECT 689.845 219.760 690.015 219.930 ;
        RECT 690.305 219.760 690.475 219.930 ;
        RECT 690.765 219.760 690.935 219.930 ;
        RECT 691.225 219.760 691.395 219.930 ;
        RECT 691.685 219.760 691.855 219.930 ;
        RECT 692.145 219.760 692.315 219.930 ;
        RECT 692.605 219.760 692.775 219.930 ;
        RECT 693.985 219.760 694.155 219.930 ;
        RECT 694.445 219.760 694.615 219.930 ;
        RECT 694.905 219.760 695.075 219.930 ;
        RECT 695.365 219.760 695.535 219.930 ;
        RECT 695.825 219.760 695.995 219.930 ;
        RECT 696.285 219.760 696.455 219.930 ;
        RECT 696.745 219.760 696.915 219.930 ;
        RECT 697.205 219.760 697.375 219.930 ;
        RECT 697.665 219.760 697.835 219.930 ;
        RECT 698.125 219.760 698.295 219.930 ;
        RECT 698.585 219.760 698.755 219.930 ;
        RECT 699.965 219.760 700.135 219.930 ;
        RECT 700.425 219.760 700.595 219.930 ;
        RECT 700.885 219.760 701.055 219.930 ;
        RECT 701.345 219.760 701.515 219.930 ;
        RECT 701.805 219.760 701.975 219.930 ;
        RECT 702.265 219.760 702.435 219.930 ;
        RECT 702.725 219.760 702.895 219.930 ;
        RECT 703.185 219.760 703.355 219.930 ;
        RECT 703.645 219.760 703.815 219.930 ;
        RECT 704.105 219.760 704.275 219.930 ;
        RECT 704.565 219.760 704.735 219.930 ;
        RECT 705.945 219.760 706.115 219.930 ;
        RECT 706.405 219.760 706.575 219.930 ;
        RECT 706.865 219.760 707.035 219.930 ;
        RECT 707.325 219.760 707.495 219.930 ;
        RECT 707.785 219.760 707.955 219.930 ;
        RECT 708.245 219.760 708.415 219.930 ;
        RECT 708.705 219.760 708.875 219.930 ;
        RECT 709.165 219.760 709.335 219.930 ;
        RECT 709.625 219.760 709.795 219.930 ;
        RECT 710.085 219.760 710.255 219.930 ;
        RECT 710.545 219.760 710.715 219.930 ;
        RECT 711.925 219.760 712.095 219.930 ;
        RECT 712.385 219.760 712.555 219.930 ;
        RECT 712.845 219.760 713.015 219.930 ;
        RECT 713.305 219.760 713.475 219.930 ;
        RECT 713.765 219.760 713.935 219.930 ;
        RECT 714.225 219.760 714.395 219.930 ;
        RECT 714.685 219.760 714.855 219.930 ;
        RECT 715.145 219.760 715.315 219.930 ;
        RECT 715.605 219.760 715.775 219.930 ;
        RECT 716.065 219.760 716.235 219.930 ;
        RECT 716.525 219.760 716.695 219.930 ;
        RECT 717.905 219.760 718.075 219.930 ;
        RECT 718.365 219.760 718.535 219.930 ;
        RECT 718.825 219.760 718.995 219.930 ;
        RECT 719.285 219.760 719.455 219.930 ;
        RECT 719.745 219.760 719.915 219.930 ;
        RECT 720.205 219.760 720.375 219.930 ;
        RECT 720.665 219.760 720.835 219.930 ;
        RECT 721.125 219.760 721.295 219.930 ;
        RECT 721.585 219.760 721.755 219.930 ;
        RECT 722.045 219.760 722.215 219.930 ;
        RECT 722.505 219.760 722.675 219.930 ;
        RECT 723.885 219.760 724.055 219.930 ;
        RECT 724.345 219.760 724.515 219.930 ;
        RECT 724.805 219.760 724.975 219.930 ;
        RECT 725.265 219.760 725.435 219.930 ;
        RECT 725.725 219.760 725.895 219.930 ;
        RECT 726.185 219.760 726.355 219.930 ;
        RECT 726.645 219.760 726.815 219.930 ;
        RECT 727.105 219.760 727.275 219.930 ;
        RECT 727.565 219.760 727.735 219.930 ;
        RECT 728.025 219.760 728.195 219.930 ;
        RECT 728.485 219.760 728.655 219.930 ;
        RECT 729.865 219.760 730.035 219.930 ;
        RECT 730.325 219.760 730.495 219.930 ;
        RECT 730.785 219.760 730.955 219.930 ;
        RECT 731.245 219.760 731.415 219.930 ;
        RECT 731.705 219.760 731.875 219.930 ;
        RECT 732.165 219.760 732.335 219.930 ;
        RECT 732.625 219.760 732.795 219.930 ;
        RECT 733.085 219.760 733.255 219.930 ;
        RECT 733.545 219.760 733.715 219.930 ;
        RECT 734.005 219.760 734.175 219.930 ;
        RECT 734.465 219.760 734.635 219.930 ;
        RECT 735.845 219.760 736.015 219.930 ;
        RECT 736.305 219.760 736.475 219.930 ;
        RECT 736.765 219.760 736.935 219.930 ;
        RECT 737.225 219.760 737.395 219.930 ;
        RECT 737.685 219.760 737.855 219.930 ;
        RECT 738.145 219.760 738.315 219.930 ;
        RECT 738.605 219.760 738.775 219.930 ;
        RECT 739.065 219.760 739.235 219.930 ;
        RECT 739.525 219.760 739.695 219.930 ;
        RECT 739.985 219.760 740.155 219.930 ;
        RECT 740.445 219.760 740.615 219.930 ;
        RECT 741.825 219.760 741.995 219.930 ;
        RECT 742.285 219.760 742.455 219.930 ;
        RECT 742.745 219.760 742.915 219.930 ;
        RECT 743.205 219.760 743.375 219.930 ;
        RECT 743.665 219.760 743.835 219.930 ;
        RECT 744.125 219.760 744.295 219.930 ;
        RECT 744.585 219.760 744.755 219.930 ;
        RECT 745.045 219.760 745.215 219.930 ;
        RECT 745.505 219.760 745.675 219.930 ;
        RECT 745.965 219.760 746.135 219.930 ;
        RECT 746.425 219.760 746.595 219.930 ;
        RECT 747.805 219.760 747.975 219.930 ;
        RECT 748.265 219.760 748.435 219.930 ;
        RECT 748.725 219.760 748.895 219.930 ;
        RECT 749.185 219.760 749.355 219.930 ;
        RECT 749.645 219.760 749.815 219.930 ;
        RECT 750.105 219.760 750.275 219.930 ;
        RECT 750.565 219.760 750.735 219.930 ;
        RECT 751.025 219.760 751.195 219.930 ;
        RECT 751.485 219.760 751.655 219.930 ;
        RECT 751.945 219.760 752.115 219.930 ;
        RECT 752.405 219.760 752.575 219.930 ;
        RECT 753.785 219.760 753.955 219.930 ;
        RECT 754.245 219.760 754.415 219.930 ;
        RECT 754.705 219.760 754.875 219.930 ;
        RECT 755.165 219.760 755.335 219.930 ;
        RECT 755.625 219.760 755.795 219.930 ;
        RECT 756.085 219.760 756.255 219.930 ;
        RECT 756.545 219.760 756.715 219.930 ;
        RECT 757.005 219.760 757.175 219.930 ;
        RECT 757.465 219.760 757.635 219.930 ;
        RECT 757.925 219.760 758.095 219.930 ;
        RECT 758.385 219.760 758.555 219.930 ;
        RECT 759.765 219.760 759.935 219.930 ;
        RECT 760.225 219.760 760.395 219.930 ;
        RECT 760.685 219.760 760.855 219.930 ;
        RECT 761.145 219.760 761.315 219.930 ;
        RECT 761.605 219.760 761.775 219.930 ;
        RECT 762.065 219.760 762.235 219.930 ;
        RECT 762.525 219.760 762.695 219.930 ;
        RECT 762.985 219.760 763.155 219.930 ;
        RECT 763.445 219.760 763.615 219.930 ;
        RECT 763.905 219.760 764.075 219.930 ;
        RECT 764.365 219.760 764.535 219.930 ;
        RECT 765.745 219.760 765.915 219.930 ;
        RECT 766.205 219.760 766.375 219.930 ;
        RECT 766.665 219.760 766.835 219.930 ;
        RECT 767.125 219.760 767.295 219.930 ;
        RECT 767.585 219.760 767.755 219.930 ;
        RECT 768.045 219.760 768.215 219.930 ;
        RECT 768.505 219.760 768.675 219.930 ;
        RECT 768.965 219.760 769.135 219.930 ;
        RECT 769.425 219.760 769.595 219.930 ;
        RECT 769.885 219.760 770.055 219.930 ;
        RECT 770.345 219.760 770.515 219.930 ;
        RECT 771.725 219.760 771.895 219.930 ;
        RECT 772.185 219.760 772.355 219.930 ;
        RECT 772.645 219.760 772.815 219.930 ;
        RECT 773.105 219.760 773.275 219.930 ;
        RECT 773.565 219.760 773.735 219.930 ;
        RECT 774.025 219.760 774.195 219.930 ;
        RECT 774.485 219.760 774.655 219.930 ;
        RECT 774.945 219.760 775.115 219.930 ;
        RECT 775.405 219.760 775.575 219.930 ;
        RECT 775.865 219.760 776.035 219.930 ;
        RECT 776.325 219.760 776.495 219.930 ;
        RECT 777.705 219.760 777.875 219.930 ;
        RECT 778.165 219.760 778.335 219.930 ;
        RECT 778.625 219.760 778.795 219.930 ;
        RECT 779.085 219.760 779.255 219.930 ;
        RECT 779.545 219.760 779.715 219.930 ;
        RECT 780.005 219.760 780.175 219.930 ;
        RECT 780.465 219.760 780.635 219.930 ;
        RECT 780.925 219.760 781.095 219.930 ;
        RECT 781.385 219.760 781.555 219.930 ;
        RECT 781.845 219.760 782.015 219.930 ;
        RECT 782.305 219.760 782.475 219.930 ;
        RECT 783.685 219.760 783.855 219.930 ;
        RECT 784.145 219.760 784.315 219.930 ;
        RECT 784.605 219.760 784.775 219.930 ;
        RECT 785.065 219.760 785.235 219.930 ;
        RECT 785.525 219.760 785.695 219.930 ;
        RECT 785.985 219.760 786.155 219.930 ;
        RECT 786.445 219.760 786.615 219.930 ;
        RECT 786.905 219.760 787.075 219.930 ;
        RECT 787.365 219.760 787.535 219.930 ;
        RECT 787.825 219.760 787.995 219.930 ;
        RECT 788.285 219.760 788.455 219.930 ;
        RECT 789.665 219.760 789.835 219.930 ;
        RECT 790.125 219.760 790.295 219.930 ;
        RECT 790.585 219.760 790.755 219.930 ;
        RECT 791.045 219.760 791.215 219.930 ;
        RECT 791.505 219.760 791.675 219.930 ;
        RECT 791.965 219.760 792.135 219.930 ;
        RECT 792.425 219.760 792.595 219.930 ;
        RECT 792.885 219.760 793.055 219.930 ;
        RECT 793.345 219.760 793.515 219.930 ;
        RECT 793.805 219.760 793.975 219.930 ;
        RECT 794.265 219.760 794.435 219.930 ;
      LAYER met1 ;
        RECT 669.000 219.605 795.040 220.085 ;
        RECT 669.000 214.165 795.040 214.645 ;
      LAYER via ;
        RECT 730.995 219.720 732.780 220.020 ;
        RECT 730.995 214.280 732.780 214.580 ;
      LAYER met2 ;
        RECT 730.955 219.660 732.820 220.090 ;
        RECT 730.955 214.220 732.820 214.650 ;
      LAYER via2 ;
        RECT 730.995 219.720 732.780 220.020 ;
        RECT 730.995 214.280 732.780 214.580 ;
      LAYER met3 ;
        RECT 730.965 209.835 732.815 220.090 ;
    END
    PORT
      LAYER li1 ;
        RECT 2146.145 219.760 2146.315 219.930 ;
      LAYER li1 ;
        RECT 2146.460 219.760 2151.980 219.930 ;
      LAYER li1 ;
        RECT 2152.125 219.760 2152.295 219.930 ;
      LAYER li1 ;
        RECT 2152.440 219.760 2157.960 219.930 ;
      LAYER li1 ;
        RECT 2158.105 219.760 2158.275 219.930 ;
      LAYER li1 ;
        RECT 2158.420 219.760 2163.940 219.930 ;
      LAYER li1 ;
        RECT 2164.085 219.760 2164.255 219.930 ;
      LAYER li1 ;
        RECT 2164.400 219.760 2169.920 219.930 ;
      LAYER li1 ;
        RECT 2170.065 219.760 2170.235 219.930 ;
      LAYER li1 ;
        RECT 2170.380 219.760 2175.900 219.930 ;
      LAYER li1 ;
        RECT 2176.045 219.760 2176.215 219.930 ;
      LAYER li1 ;
        RECT 2176.360 219.760 2181.880 219.930 ;
      LAYER li1 ;
        RECT 2182.025 219.760 2182.195 219.930 ;
      LAYER li1 ;
        RECT 2182.340 219.760 2187.860 219.930 ;
      LAYER li1 ;
        RECT 2188.005 219.760 2188.175 219.930 ;
      LAYER li1 ;
        RECT 2188.320 219.760 2193.840 219.930 ;
      LAYER li1 ;
        RECT 2193.985 219.760 2194.155 219.930 ;
      LAYER li1 ;
        RECT 2194.300 219.760 2199.820 219.930 ;
      LAYER li1 ;
        RECT 2199.965 219.760 2200.135 219.930 ;
      LAYER li1 ;
        RECT 2200.280 219.760 2205.800 219.930 ;
      LAYER li1 ;
        RECT 2205.945 219.760 2206.115 219.930 ;
      LAYER li1 ;
        RECT 2206.260 219.760 2211.780 219.930 ;
      LAYER li1 ;
        RECT 2211.925 219.760 2212.095 219.930 ;
      LAYER li1 ;
        RECT 2212.240 219.760 2217.760 219.930 ;
      LAYER li1 ;
        RECT 2217.905 219.760 2218.075 219.930 ;
      LAYER li1 ;
        RECT 2218.220 219.760 2223.740 219.930 ;
      LAYER li1 ;
        RECT 2223.885 219.760 2224.055 219.930 ;
      LAYER li1 ;
        RECT 2224.200 219.760 2229.720 219.930 ;
      LAYER li1 ;
        RECT 2229.865 219.760 2230.035 219.930 ;
      LAYER li1 ;
        RECT 2230.180 219.760 2235.700 219.930 ;
      LAYER li1 ;
        RECT 2235.845 219.760 2236.015 219.930 ;
      LAYER li1 ;
        RECT 2236.160 219.760 2241.680 219.930 ;
      LAYER li1 ;
        RECT 2241.825 219.760 2241.995 219.930 ;
      LAYER li1 ;
        RECT 2242.140 219.760 2247.660 219.930 ;
      LAYER li1 ;
        RECT 2247.805 219.760 2247.975 219.930 ;
      LAYER li1 ;
        RECT 2248.120 219.760 2253.640 219.930 ;
      LAYER li1 ;
        RECT 2253.785 219.760 2253.955 219.930 ;
      LAYER li1 ;
        RECT 2254.100 219.760 2259.620 219.930 ;
      LAYER li1 ;
        RECT 2259.765 219.760 2259.935 219.930 ;
      LAYER li1 ;
        RECT 2260.080 219.760 2265.600 219.930 ;
      LAYER li1 ;
        RECT 2265.745 219.760 2265.915 219.930 ;
      LAYER li1 ;
        RECT 2266.060 219.760 2271.580 219.930 ;
      LAYER li1 ;
        RECT 2271.725 219.760 2271.895 219.930 ;
      LAYER li1 ;
        RECT 2146.545 219.325 2151.890 219.760 ;
        RECT 2152.525 219.325 2157.870 219.760 ;
        RECT 2158.505 219.325 2163.850 219.760 ;
        RECT 2164.485 219.325 2169.830 219.760 ;
        RECT 2170.465 219.325 2175.810 219.760 ;
        RECT 2176.445 219.325 2181.790 219.760 ;
        RECT 2182.425 219.325 2187.770 219.760 ;
        RECT 2188.405 219.325 2193.750 219.760 ;
        RECT 2194.385 219.325 2199.730 219.760 ;
        RECT 2200.365 219.325 2205.710 219.760 ;
        RECT 2206.345 219.325 2211.690 219.760 ;
        RECT 2212.325 219.325 2217.670 219.760 ;
        RECT 2218.305 219.325 2223.650 219.760 ;
        RECT 2224.285 219.325 2229.630 219.760 ;
        RECT 2230.265 219.325 2235.610 219.760 ;
        RECT 2236.245 219.325 2241.590 219.760 ;
        RECT 2242.225 219.325 2247.570 219.760 ;
        RECT 2248.205 219.325 2253.550 219.760 ;
        RECT 2254.185 219.325 2259.530 219.760 ;
        RECT 2260.165 219.325 2265.510 219.760 ;
        RECT 2266.145 219.325 2271.490 219.760 ;
        RECT 2149.950 218.075 2150.300 219.325 ;
        RECT 2155.930 218.075 2156.280 219.325 ;
        RECT 2161.910 218.075 2162.260 219.325 ;
        RECT 2167.890 218.075 2168.240 219.325 ;
        RECT 2173.870 218.075 2174.220 219.325 ;
        RECT 2179.850 218.075 2180.200 219.325 ;
        RECT 2185.830 218.075 2186.180 219.325 ;
        RECT 2191.810 218.075 2192.160 219.325 ;
        RECT 2197.790 218.075 2198.140 219.325 ;
        RECT 2203.770 218.075 2204.120 219.325 ;
        RECT 2209.750 218.075 2210.100 219.325 ;
        RECT 2215.730 218.075 2216.080 219.325 ;
        RECT 2221.710 218.075 2222.060 219.325 ;
        RECT 2227.690 218.075 2228.040 219.325 ;
        RECT 2233.670 218.075 2234.020 219.325 ;
        RECT 2239.650 218.075 2240.000 219.325 ;
        RECT 2245.630 218.075 2245.980 219.325 ;
        RECT 2251.610 218.075 2251.960 219.325 ;
        RECT 2257.590 218.075 2257.940 219.325 ;
        RECT 2263.570 218.075 2263.920 219.325 ;
        RECT 2269.550 218.075 2269.900 219.325 ;
      LAYER li1 ;
        RECT 2146.145 214.320 2146.315 214.490 ;
        RECT 2146.605 214.320 2146.775 214.490 ;
        RECT 2147.065 214.320 2147.235 214.490 ;
        RECT 2147.525 214.320 2147.695 214.490 ;
        RECT 2147.985 214.320 2148.155 214.490 ;
        RECT 2148.445 214.320 2148.615 214.490 ;
        RECT 2148.905 214.320 2149.075 214.490 ;
        RECT 2149.365 214.320 2149.535 214.490 ;
        RECT 2149.825 214.320 2149.995 214.490 ;
        RECT 2150.285 214.320 2150.455 214.490 ;
        RECT 2150.745 214.320 2150.915 214.490 ;
        RECT 2151.205 214.320 2151.375 214.490 ;
        RECT 2151.665 214.320 2151.835 214.490 ;
        RECT 2152.125 214.320 2152.295 214.490 ;
        RECT 2152.585 214.320 2152.755 214.490 ;
        RECT 2153.045 214.320 2153.215 214.490 ;
        RECT 2153.505 214.320 2153.675 214.490 ;
        RECT 2153.965 214.320 2154.135 214.490 ;
        RECT 2154.425 214.320 2154.595 214.490 ;
        RECT 2154.885 214.320 2155.055 214.490 ;
        RECT 2155.345 214.320 2155.515 214.490 ;
        RECT 2155.805 214.320 2155.975 214.490 ;
        RECT 2156.265 214.320 2156.435 214.490 ;
        RECT 2156.725 214.320 2156.895 214.490 ;
        RECT 2157.185 214.320 2157.355 214.490 ;
        RECT 2157.645 214.320 2157.815 214.490 ;
        RECT 2158.105 214.320 2158.275 214.490 ;
        RECT 2158.565 214.320 2158.735 214.490 ;
        RECT 2159.025 214.320 2159.195 214.490 ;
        RECT 2159.485 214.320 2159.655 214.490 ;
        RECT 2159.945 214.320 2160.115 214.490 ;
        RECT 2160.405 214.320 2160.575 214.490 ;
        RECT 2160.865 214.320 2161.035 214.490 ;
        RECT 2161.325 214.320 2161.495 214.490 ;
        RECT 2161.785 214.320 2161.955 214.490 ;
        RECT 2162.245 214.320 2162.415 214.490 ;
        RECT 2162.705 214.320 2162.875 214.490 ;
        RECT 2163.165 214.320 2163.335 214.490 ;
        RECT 2163.625 214.320 2163.795 214.490 ;
        RECT 2164.085 214.320 2164.255 214.490 ;
        RECT 2164.545 214.320 2164.715 214.490 ;
        RECT 2165.005 214.320 2165.175 214.490 ;
        RECT 2165.465 214.320 2165.635 214.490 ;
        RECT 2165.925 214.320 2166.095 214.490 ;
        RECT 2166.385 214.320 2166.555 214.490 ;
        RECT 2166.845 214.320 2167.015 214.490 ;
        RECT 2167.305 214.320 2167.475 214.490 ;
        RECT 2167.765 214.320 2167.935 214.490 ;
        RECT 2168.225 214.320 2168.395 214.490 ;
        RECT 2168.685 214.320 2168.855 214.490 ;
        RECT 2169.145 214.320 2169.315 214.490 ;
        RECT 2169.605 214.320 2169.775 214.490 ;
        RECT 2170.065 214.320 2170.235 214.490 ;
        RECT 2170.525 214.320 2170.695 214.490 ;
        RECT 2170.985 214.320 2171.155 214.490 ;
        RECT 2171.445 214.320 2171.615 214.490 ;
        RECT 2171.905 214.320 2172.075 214.490 ;
        RECT 2172.365 214.320 2172.535 214.490 ;
        RECT 2172.825 214.320 2172.995 214.490 ;
        RECT 2173.285 214.320 2173.455 214.490 ;
        RECT 2173.745 214.320 2173.915 214.490 ;
        RECT 2174.205 214.320 2174.375 214.490 ;
        RECT 2174.665 214.320 2174.835 214.490 ;
        RECT 2175.125 214.320 2175.295 214.490 ;
        RECT 2175.585 214.320 2175.755 214.490 ;
        RECT 2176.045 214.320 2176.215 214.490 ;
        RECT 2176.505 214.320 2176.675 214.490 ;
        RECT 2176.965 214.320 2177.135 214.490 ;
        RECT 2177.425 214.320 2177.595 214.490 ;
        RECT 2177.885 214.320 2178.055 214.490 ;
        RECT 2178.345 214.320 2178.515 214.490 ;
        RECT 2178.805 214.320 2178.975 214.490 ;
        RECT 2179.265 214.320 2179.435 214.490 ;
        RECT 2179.725 214.320 2179.895 214.490 ;
        RECT 2180.185 214.320 2180.355 214.490 ;
        RECT 2180.645 214.320 2180.815 214.490 ;
        RECT 2181.105 214.320 2181.275 214.490 ;
        RECT 2181.565 214.320 2181.735 214.490 ;
        RECT 2182.025 214.320 2182.195 214.490 ;
        RECT 2182.485 214.320 2182.655 214.490 ;
        RECT 2182.945 214.320 2183.115 214.490 ;
        RECT 2183.405 214.320 2183.575 214.490 ;
        RECT 2183.865 214.320 2184.035 214.490 ;
        RECT 2184.325 214.320 2184.495 214.490 ;
        RECT 2184.785 214.320 2184.955 214.490 ;
        RECT 2185.245 214.320 2185.415 214.490 ;
        RECT 2185.705 214.320 2185.875 214.490 ;
        RECT 2186.165 214.320 2186.335 214.490 ;
        RECT 2186.625 214.320 2186.795 214.490 ;
        RECT 2187.085 214.320 2187.255 214.490 ;
        RECT 2187.545 214.320 2187.715 214.490 ;
        RECT 2188.005 214.320 2188.175 214.490 ;
        RECT 2188.465 214.320 2188.635 214.490 ;
        RECT 2188.925 214.320 2189.095 214.490 ;
        RECT 2189.385 214.320 2189.555 214.490 ;
        RECT 2189.845 214.320 2190.015 214.490 ;
        RECT 2190.305 214.320 2190.475 214.490 ;
        RECT 2190.765 214.320 2190.935 214.490 ;
        RECT 2191.225 214.320 2191.395 214.490 ;
        RECT 2191.685 214.320 2191.855 214.490 ;
        RECT 2192.145 214.320 2192.315 214.490 ;
        RECT 2192.605 214.320 2192.775 214.490 ;
        RECT 2193.065 214.320 2193.235 214.490 ;
        RECT 2193.525 214.320 2193.695 214.490 ;
        RECT 2193.985 214.320 2194.155 214.490 ;
        RECT 2194.445 214.320 2194.615 214.490 ;
        RECT 2194.905 214.320 2195.075 214.490 ;
        RECT 2195.365 214.320 2195.535 214.490 ;
        RECT 2195.825 214.320 2195.995 214.490 ;
        RECT 2196.285 214.320 2196.455 214.490 ;
        RECT 2196.745 214.320 2196.915 214.490 ;
        RECT 2197.205 214.320 2197.375 214.490 ;
        RECT 2197.665 214.320 2197.835 214.490 ;
        RECT 2198.125 214.320 2198.295 214.490 ;
        RECT 2198.585 214.320 2198.755 214.490 ;
        RECT 2199.045 214.320 2199.215 214.490 ;
        RECT 2199.505 214.320 2199.675 214.490 ;
        RECT 2199.965 214.320 2200.135 214.490 ;
        RECT 2200.425 214.320 2200.595 214.490 ;
        RECT 2200.885 214.320 2201.055 214.490 ;
        RECT 2201.345 214.320 2201.515 214.490 ;
        RECT 2201.805 214.320 2201.975 214.490 ;
        RECT 2202.265 214.320 2202.435 214.490 ;
        RECT 2202.725 214.320 2202.895 214.490 ;
        RECT 2203.185 214.320 2203.355 214.490 ;
        RECT 2203.645 214.320 2203.815 214.490 ;
        RECT 2204.105 214.320 2204.275 214.490 ;
        RECT 2204.565 214.320 2204.735 214.490 ;
        RECT 2205.025 214.320 2205.195 214.490 ;
        RECT 2205.485 214.320 2205.655 214.490 ;
        RECT 2205.945 214.320 2206.115 214.490 ;
        RECT 2206.405 214.320 2206.575 214.490 ;
        RECT 2206.865 214.320 2207.035 214.490 ;
        RECT 2207.325 214.320 2207.495 214.490 ;
        RECT 2207.785 214.320 2207.955 214.490 ;
        RECT 2208.245 214.320 2208.415 214.490 ;
        RECT 2208.705 214.320 2208.875 214.490 ;
        RECT 2209.165 214.320 2209.335 214.490 ;
        RECT 2209.625 214.320 2209.795 214.490 ;
        RECT 2210.085 214.320 2210.255 214.490 ;
        RECT 2210.545 214.320 2210.715 214.490 ;
        RECT 2211.005 214.320 2211.175 214.490 ;
        RECT 2211.465 214.320 2211.635 214.490 ;
        RECT 2211.925 214.320 2212.095 214.490 ;
        RECT 2212.385 214.320 2212.555 214.490 ;
        RECT 2212.845 214.320 2213.015 214.490 ;
        RECT 2213.305 214.320 2213.475 214.490 ;
        RECT 2213.765 214.320 2213.935 214.490 ;
        RECT 2214.225 214.320 2214.395 214.490 ;
        RECT 2214.685 214.320 2214.855 214.490 ;
        RECT 2215.145 214.320 2215.315 214.490 ;
        RECT 2215.605 214.320 2215.775 214.490 ;
        RECT 2216.065 214.320 2216.235 214.490 ;
        RECT 2216.525 214.320 2216.695 214.490 ;
        RECT 2216.985 214.320 2217.155 214.490 ;
        RECT 2217.445 214.320 2217.615 214.490 ;
        RECT 2217.905 214.320 2218.075 214.490 ;
        RECT 2218.365 214.320 2218.535 214.490 ;
        RECT 2218.825 214.320 2218.995 214.490 ;
        RECT 2219.285 214.320 2219.455 214.490 ;
        RECT 2219.745 214.320 2219.915 214.490 ;
        RECT 2220.205 214.320 2220.375 214.490 ;
        RECT 2220.665 214.320 2220.835 214.490 ;
        RECT 2221.125 214.320 2221.295 214.490 ;
        RECT 2221.585 214.320 2221.755 214.490 ;
        RECT 2222.045 214.320 2222.215 214.490 ;
        RECT 2222.505 214.320 2222.675 214.490 ;
        RECT 2222.965 214.320 2223.135 214.490 ;
        RECT 2223.425 214.320 2223.595 214.490 ;
        RECT 2223.885 214.320 2224.055 214.490 ;
        RECT 2224.345 214.320 2224.515 214.490 ;
        RECT 2224.805 214.320 2224.975 214.490 ;
        RECT 2225.265 214.320 2225.435 214.490 ;
        RECT 2225.725 214.320 2225.895 214.490 ;
        RECT 2226.185 214.320 2226.355 214.490 ;
        RECT 2226.645 214.320 2226.815 214.490 ;
        RECT 2227.105 214.320 2227.275 214.490 ;
        RECT 2227.565 214.320 2227.735 214.490 ;
        RECT 2228.025 214.320 2228.195 214.490 ;
        RECT 2228.485 214.320 2228.655 214.490 ;
        RECT 2228.945 214.320 2229.115 214.490 ;
        RECT 2229.405 214.320 2229.575 214.490 ;
        RECT 2229.865 214.320 2230.035 214.490 ;
        RECT 2230.325 214.320 2230.495 214.490 ;
        RECT 2230.785 214.320 2230.955 214.490 ;
        RECT 2231.245 214.320 2231.415 214.490 ;
        RECT 2231.705 214.320 2231.875 214.490 ;
        RECT 2232.165 214.320 2232.335 214.490 ;
        RECT 2232.625 214.320 2232.795 214.490 ;
        RECT 2233.085 214.320 2233.255 214.490 ;
        RECT 2233.545 214.320 2233.715 214.490 ;
        RECT 2234.005 214.320 2234.175 214.490 ;
        RECT 2234.465 214.320 2234.635 214.490 ;
        RECT 2234.925 214.320 2235.095 214.490 ;
        RECT 2235.385 214.320 2235.555 214.490 ;
        RECT 2235.845 214.320 2236.015 214.490 ;
        RECT 2236.305 214.320 2236.475 214.490 ;
        RECT 2236.765 214.320 2236.935 214.490 ;
        RECT 2237.225 214.320 2237.395 214.490 ;
        RECT 2237.685 214.320 2237.855 214.490 ;
        RECT 2238.145 214.320 2238.315 214.490 ;
        RECT 2238.605 214.320 2238.775 214.490 ;
        RECT 2239.065 214.320 2239.235 214.490 ;
        RECT 2239.525 214.320 2239.695 214.490 ;
        RECT 2239.985 214.320 2240.155 214.490 ;
        RECT 2240.445 214.320 2240.615 214.490 ;
        RECT 2240.905 214.320 2241.075 214.490 ;
        RECT 2241.365 214.320 2241.535 214.490 ;
        RECT 2241.825 214.320 2241.995 214.490 ;
        RECT 2242.285 214.320 2242.455 214.490 ;
        RECT 2242.745 214.320 2242.915 214.490 ;
        RECT 2243.205 214.320 2243.375 214.490 ;
        RECT 2243.665 214.320 2243.835 214.490 ;
        RECT 2244.125 214.320 2244.295 214.490 ;
        RECT 2244.585 214.320 2244.755 214.490 ;
        RECT 2245.045 214.320 2245.215 214.490 ;
        RECT 2245.505 214.320 2245.675 214.490 ;
        RECT 2245.965 214.320 2246.135 214.490 ;
        RECT 2246.425 214.320 2246.595 214.490 ;
        RECT 2246.885 214.320 2247.055 214.490 ;
        RECT 2247.345 214.320 2247.515 214.490 ;
        RECT 2247.805 214.320 2247.975 214.490 ;
        RECT 2248.265 214.320 2248.435 214.490 ;
        RECT 2248.725 214.320 2248.895 214.490 ;
        RECT 2249.185 214.320 2249.355 214.490 ;
        RECT 2249.645 214.320 2249.815 214.490 ;
        RECT 2250.105 214.320 2250.275 214.490 ;
        RECT 2250.565 214.320 2250.735 214.490 ;
        RECT 2251.025 214.320 2251.195 214.490 ;
        RECT 2251.485 214.320 2251.655 214.490 ;
        RECT 2251.945 214.320 2252.115 214.490 ;
        RECT 2252.405 214.320 2252.575 214.490 ;
        RECT 2252.865 214.320 2253.035 214.490 ;
        RECT 2253.325 214.320 2253.495 214.490 ;
        RECT 2253.785 214.320 2253.955 214.490 ;
        RECT 2254.245 214.320 2254.415 214.490 ;
        RECT 2254.705 214.320 2254.875 214.490 ;
        RECT 2255.165 214.320 2255.335 214.490 ;
        RECT 2255.625 214.320 2255.795 214.490 ;
        RECT 2256.085 214.320 2256.255 214.490 ;
        RECT 2256.545 214.320 2256.715 214.490 ;
        RECT 2257.005 214.320 2257.175 214.490 ;
        RECT 2257.465 214.320 2257.635 214.490 ;
        RECT 2257.925 214.320 2258.095 214.490 ;
        RECT 2258.385 214.320 2258.555 214.490 ;
        RECT 2258.845 214.320 2259.015 214.490 ;
        RECT 2259.305 214.320 2259.475 214.490 ;
        RECT 2259.765 214.320 2259.935 214.490 ;
        RECT 2260.225 214.320 2260.395 214.490 ;
        RECT 2260.685 214.320 2260.855 214.490 ;
        RECT 2261.145 214.320 2261.315 214.490 ;
        RECT 2261.605 214.320 2261.775 214.490 ;
        RECT 2262.065 214.320 2262.235 214.490 ;
        RECT 2262.525 214.320 2262.695 214.490 ;
        RECT 2262.985 214.320 2263.155 214.490 ;
        RECT 2263.445 214.320 2263.615 214.490 ;
        RECT 2263.905 214.320 2264.075 214.490 ;
        RECT 2264.365 214.320 2264.535 214.490 ;
        RECT 2264.825 214.320 2264.995 214.490 ;
        RECT 2265.285 214.320 2265.455 214.490 ;
        RECT 2265.745 214.320 2265.915 214.490 ;
        RECT 2266.205 214.320 2266.375 214.490 ;
        RECT 2266.665 214.320 2266.835 214.490 ;
        RECT 2267.125 214.320 2267.295 214.490 ;
        RECT 2267.585 214.320 2267.755 214.490 ;
        RECT 2268.045 214.320 2268.215 214.490 ;
        RECT 2268.505 214.320 2268.675 214.490 ;
        RECT 2268.965 214.320 2269.135 214.490 ;
        RECT 2269.425 214.320 2269.595 214.490 ;
        RECT 2269.885 214.320 2270.055 214.490 ;
        RECT 2270.345 214.320 2270.515 214.490 ;
        RECT 2270.805 214.320 2270.975 214.490 ;
        RECT 2271.265 214.320 2271.435 214.490 ;
        RECT 2271.725 214.320 2271.895 214.490 ;
      LAYER mcon ;
        RECT 2147.065 219.760 2147.235 219.930 ;
        RECT 2147.525 219.760 2147.695 219.930 ;
        RECT 2147.985 219.760 2148.155 219.930 ;
        RECT 2148.445 219.760 2148.615 219.930 ;
        RECT 2148.905 219.760 2149.075 219.930 ;
        RECT 2149.365 219.760 2149.535 219.930 ;
        RECT 2149.825 219.760 2149.995 219.930 ;
        RECT 2150.285 219.760 2150.455 219.930 ;
        RECT 2150.745 219.760 2150.915 219.930 ;
        RECT 2151.205 219.760 2151.375 219.930 ;
        RECT 2151.665 219.760 2151.835 219.930 ;
        RECT 2153.045 219.760 2153.215 219.930 ;
        RECT 2153.505 219.760 2153.675 219.930 ;
        RECT 2153.965 219.760 2154.135 219.930 ;
        RECT 2154.425 219.760 2154.595 219.930 ;
        RECT 2154.885 219.760 2155.055 219.930 ;
        RECT 2155.345 219.760 2155.515 219.930 ;
        RECT 2155.805 219.760 2155.975 219.930 ;
        RECT 2156.265 219.760 2156.435 219.930 ;
        RECT 2156.725 219.760 2156.895 219.930 ;
        RECT 2157.185 219.760 2157.355 219.930 ;
        RECT 2157.645 219.760 2157.815 219.930 ;
        RECT 2159.025 219.760 2159.195 219.930 ;
        RECT 2159.485 219.760 2159.655 219.930 ;
        RECT 2159.945 219.760 2160.115 219.930 ;
        RECT 2160.405 219.760 2160.575 219.930 ;
        RECT 2160.865 219.760 2161.035 219.930 ;
        RECT 2161.325 219.760 2161.495 219.930 ;
        RECT 2161.785 219.760 2161.955 219.930 ;
        RECT 2162.245 219.760 2162.415 219.930 ;
        RECT 2162.705 219.760 2162.875 219.930 ;
        RECT 2163.165 219.760 2163.335 219.930 ;
        RECT 2163.625 219.760 2163.795 219.930 ;
        RECT 2165.005 219.760 2165.175 219.930 ;
        RECT 2165.465 219.760 2165.635 219.930 ;
        RECT 2165.925 219.760 2166.095 219.930 ;
        RECT 2166.385 219.760 2166.555 219.930 ;
        RECT 2166.845 219.760 2167.015 219.930 ;
        RECT 2167.305 219.760 2167.475 219.930 ;
        RECT 2167.765 219.760 2167.935 219.930 ;
        RECT 2168.225 219.760 2168.395 219.930 ;
        RECT 2168.685 219.760 2168.855 219.930 ;
        RECT 2169.145 219.760 2169.315 219.930 ;
        RECT 2169.605 219.760 2169.775 219.930 ;
        RECT 2170.985 219.760 2171.155 219.930 ;
        RECT 2171.445 219.760 2171.615 219.930 ;
        RECT 2171.905 219.760 2172.075 219.930 ;
        RECT 2172.365 219.760 2172.535 219.930 ;
        RECT 2172.825 219.760 2172.995 219.930 ;
        RECT 2173.285 219.760 2173.455 219.930 ;
        RECT 2173.745 219.760 2173.915 219.930 ;
        RECT 2174.205 219.760 2174.375 219.930 ;
        RECT 2174.665 219.760 2174.835 219.930 ;
        RECT 2175.125 219.760 2175.295 219.930 ;
        RECT 2175.585 219.760 2175.755 219.930 ;
        RECT 2176.965 219.760 2177.135 219.930 ;
        RECT 2177.425 219.760 2177.595 219.930 ;
        RECT 2177.885 219.760 2178.055 219.930 ;
        RECT 2178.345 219.760 2178.515 219.930 ;
        RECT 2178.805 219.760 2178.975 219.930 ;
        RECT 2179.265 219.760 2179.435 219.930 ;
        RECT 2179.725 219.760 2179.895 219.930 ;
        RECT 2180.185 219.760 2180.355 219.930 ;
        RECT 2180.645 219.760 2180.815 219.930 ;
        RECT 2181.105 219.760 2181.275 219.930 ;
        RECT 2181.565 219.760 2181.735 219.930 ;
        RECT 2182.945 219.760 2183.115 219.930 ;
        RECT 2183.405 219.760 2183.575 219.930 ;
        RECT 2183.865 219.760 2184.035 219.930 ;
        RECT 2184.325 219.760 2184.495 219.930 ;
        RECT 2184.785 219.760 2184.955 219.930 ;
        RECT 2185.245 219.760 2185.415 219.930 ;
        RECT 2185.705 219.760 2185.875 219.930 ;
        RECT 2186.165 219.760 2186.335 219.930 ;
        RECT 2186.625 219.760 2186.795 219.930 ;
        RECT 2187.085 219.760 2187.255 219.930 ;
        RECT 2187.545 219.760 2187.715 219.930 ;
        RECT 2188.925 219.760 2189.095 219.930 ;
        RECT 2189.385 219.760 2189.555 219.930 ;
        RECT 2189.845 219.760 2190.015 219.930 ;
        RECT 2190.305 219.760 2190.475 219.930 ;
        RECT 2190.765 219.760 2190.935 219.930 ;
        RECT 2191.225 219.760 2191.395 219.930 ;
        RECT 2191.685 219.760 2191.855 219.930 ;
        RECT 2192.145 219.760 2192.315 219.930 ;
        RECT 2192.605 219.760 2192.775 219.930 ;
        RECT 2193.065 219.760 2193.235 219.930 ;
        RECT 2193.525 219.760 2193.695 219.930 ;
        RECT 2194.905 219.760 2195.075 219.930 ;
        RECT 2195.365 219.760 2195.535 219.930 ;
        RECT 2195.825 219.760 2195.995 219.930 ;
        RECT 2196.285 219.760 2196.455 219.930 ;
        RECT 2196.745 219.760 2196.915 219.930 ;
        RECT 2197.205 219.760 2197.375 219.930 ;
        RECT 2197.665 219.760 2197.835 219.930 ;
        RECT 2198.125 219.760 2198.295 219.930 ;
        RECT 2198.585 219.760 2198.755 219.930 ;
        RECT 2199.045 219.760 2199.215 219.930 ;
        RECT 2199.505 219.760 2199.675 219.930 ;
        RECT 2200.885 219.760 2201.055 219.930 ;
        RECT 2201.345 219.760 2201.515 219.930 ;
        RECT 2201.805 219.760 2201.975 219.930 ;
        RECT 2202.265 219.760 2202.435 219.930 ;
        RECT 2202.725 219.760 2202.895 219.930 ;
        RECT 2203.185 219.760 2203.355 219.930 ;
        RECT 2203.645 219.760 2203.815 219.930 ;
        RECT 2204.105 219.760 2204.275 219.930 ;
        RECT 2204.565 219.760 2204.735 219.930 ;
        RECT 2205.025 219.760 2205.195 219.930 ;
        RECT 2205.485 219.760 2205.655 219.930 ;
        RECT 2206.865 219.760 2207.035 219.930 ;
        RECT 2207.325 219.760 2207.495 219.930 ;
        RECT 2207.785 219.760 2207.955 219.930 ;
        RECT 2208.245 219.760 2208.415 219.930 ;
        RECT 2208.705 219.760 2208.875 219.930 ;
        RECT 2209.165 219.760 2209.335 219.930 ;
        RECT 2209.625 219.760 2209.795 219.930 ;
        RECT 2210.085 219.760 2210.255 219.930 ;
        RECT 2210.545 219.760 2210.715 219.930 ;
        RECT 2211.005 219.760 2211.175 219.930 ;
        RECT 2211.465 219.760 2211.635 219.930 ;
        RECT 2212.845 219.760 2213.015 219.930 ;
        RECT 2213.305 219.760 2213.475 219.930 ;
        RECT 2213.765 219.760 2213.935 219.930 ;
        RECT 2214.225 219.760 2214.395 219.930 ;
        RECT 2214.685 219.760 2214.855 219.930 ;
        RECT 2215.145 219.760 2215.315 219.930 ;
        RECT 2215.605 219.760 2215.775 219.930 ;
        RECT 2216.065 219.760 2216.235 219.930 ;
        RECT 2216.525 219.760 2216.695 219.930 ;
        RECT 2216.985 219.760 2217.155 219.930 ;
        RECT 2217.445 219.760 2217.615 219.930 ;
        RECT 2218.825 219.760 2218.995 219.930 ;
        RECT 2219.285 219.760 2219.455 219.930 ;
        RECT 2219.745 219.760 2219.915 219.930 ;
        RECT 2220.205 219.760 2220.375 219.930 ;
        RECT 2220.665 219.760 2220.835 219.930 ;
        RECT 2221.125 219.760 2221.295 219.930 ;
        RECT 2221.585 219.760 2221.755 219.930 ;
        RECT 2222.045 219.760 2222.215 219.930 ;
        RECT 2222.505 219.760 2222.675 219.930 ;
        RECT 2222.965 219.760 2223.135 219.930 ;
        RECT 2223.425 219.760 2223.595 219.930 ;
        RECT 2224.805 219.760 2224.975 219.930 ;
        RECT 2225.265 219.760 2225.435 219.930 ;
        RECT 2225.725 219.760 2225.895 219.930 ;
        RECT 2226.185 219.760 2226.355 219.930 ;
        RECT 2226.645 219.760 2226.815 219.930 ;
        RECT 2227.105 219.760 2227.275 219.930 ;
        RECT 2227.565 219.760 2227.735 219.930 ;
        RECT 2228.025 219.760 2228.195 219.930 ;
        RECT 2228.485 219.760 2228.655 219.930 ;
        RECT 2228.945 219.760 2229.115 219.930 ;
        RECT 2229.405 219.760 2229.575 219.930 ;
        RECT 2230.785 219.760 2230.955 219.930 ;
        RECT 2231.245 219.760 2231.415 219.930 ;
        RECT 2231.705 219.760 2231.875 219.930 ;
        RECT 2232.165 219.760 2232.335 219.930 ;
        RECT 2232.625 219.760 2232.795 219.930 ;
        RECT 2233.085 219.760 2233.255 219.930 ;
        RECT 2233.545 219.760 2233.715 219.930 ;
        RECT 2234.005 219.760 2234.175 219.930 ;
        RECT 2234.465 219.760 2234.635 219.930 ;
        RECT 2234.925 219.760 2235.095 219.930 ;
        RECT 2235.385 219.760 2235.555 219.930 ;
        RECT 2236.765 219.760 2236.935 219.930 ;
        RECT 2237.225 219.760 2237.395 219.930 ;
        RECT 2237.685 219.760 2237.855 219.930 ;
        RECT 2238.145 219.760 2238.315 219.930 ;
        RECT 2238.605 219.760 2238.775 219.930 ;
        RECT 2239.065 219.760 2239.235 219.930 ;
        RECT 2239.525 219.760 2239.695 219.930 ;
        RECT 2239.985 219.760 2240.155 219.930 ;
        RECT 2240.445 219.760 2240.615 219.930 ;
        RECT 2240.905 219.760 2241.075 219.930 ;
        RECT 2241.365 219.760 2241.535 219.930 ;
        RECT 2242.745 219.760 2242.915 219.930 ;
        RECT 2243.205 219.760 2243.375 219.930 ;
        RECT 2243.665 219.760 2243.835 219.930 ;
        RECT 2244.125 219.760 2244.295 219.930 ;
        RECT 2244.585 219.760 2244.755 219.930 ;
        RECT 2245.045 219.760 2245.215 219.930 ;
        RECT 2245.505 219.760 2245.675 219.930 ;
        RECT 2245.965 219.760 2246.135 219.930 ;
        RECT 2246.425 219.760 2246.595 219.930 ;
        RECT 2246.885 219.760 2247.055 219.930 ;
        RECT 2247.345 219.760 2247.515 219.930 ;
        RECT 2248.725 219.760 2248.895 219.930 ;
        RECT 2249.185 219.760 2249.355 219.930 ;
        RECT 2249.645 219.760 2249.815 219.930 ;
        RECT 2250.105 219.760 2250.275 219.930 ;
        RECT 2250.565 219.760 2250.735 219.930 ;
        RECT 2251.025 219.760 2251.195 219.930 ;
        RECT 2251.485 219.760 2251.655 219.930 ;
        RECT 2251.945 219.760 2252.115 219.930 ;
        RECT 2252.405 219.760 2252.575 219.930 ;
        RECT 2252.865 219.760 2253.035 219.930 ;
        RECT 2253.325 219.760 2253.495 219.930 ;
        RECT 2254.705 219.760 2254.875 219.930 ;
        RECT 2255.165 219.760 2255.335 219.930 ;
        RECT 2255.625 219.760 2255.795 219.930 ;
        RECT 2256.085 219.760 2256.255 219.930 ;
        RECT 2256.545 219.760 2256.715 219.930 ;
        RECT 2257.005 219.760 2257.175 219.930 ;
        RECT 2257.465 219.760 2257.635 219.930 ;
        RECT 2257.925 219.760 2258.095 219.930 ;
        RECT 2258.385 219.760 2258.555 219.930 ;
        RECT 2258.845 219.760 2259.015 219.930 ;
        RECT 2259.305 219.760 2259.475 219.930 ;
        RECT 2260.685 219.760 2260.855 219.930 ;
        RECT 2261.145 219.760 2261.315 219.930 ;
        RECT 2261.605 219.760 2261.775 219.930 ;
        RECT 2262.065 219.760 2262.235 219.930 ;
        RECT 2262.525 219.760 2262.695 219.930 ;
        RECT 2262.985 219.760 2263.155 219.930 ;
        RECT 2263.445 219.760 2263.615 219.930 ;
        RECT 2263.905 219.760 2264.075 219.930 ;
        RECT 2264.365 219.760 2264.535 219.930 ;
        RECT 2264.825 219.760 2264.995 219.930 ;
        RECT 2265.285 219.760 2265.455 219.930 ;
        RECT 2266.665 219.760 2266.835 219.930 ;
        RECT 2267.125 219.760 2267.295 219.930 ;
        RECT 2267.585 219.760 2267.755 219.930 ;
        RECT 2268.045 219.760 2268.215 219.930 ;
        RECT 2268.505 219.760 2268.675 219.930 ;
        RECT 2268.965 219.760 2269.135 219.930 ;
        RECT 2269.425 219.760 2269.595 219.930 ;
        RECT 2269.885 219.760 2270.055 219.930 ;
        RECT 2270.345 219.760 2270.515 219.930 ;
        RECT 2270.805 219.760 2270.975 219.930 ;
        RECT 2271.265 219.760 2271.435 219.930 ;
      LAYER met1 ;
        RECT 2146.000 219.605 2272.040 220.085 ;
        RECT 2146.000 214.165 2272.040 214.645 ;
      LAYER via ;
        RECT 2202.150 219.685 2203.935 219.985 ;
        RECT 2202.150 214.245 2203.935 214.545 ;
      LAYER met2 ;
        RECT 2202.110 219.625 2203.975 220.055 ;
        RECT 2202.110 214.185 2203.975 214.615 ;
      LAYER via2 ;
        RECT 2202.150 219.685 2203.935 219.985 ;
        RECT 2202.150 214.245 2203.935 214.545 ;
      LAYER met3 ;
        RECT 2202.120 209.800 2203.970 220.055 ;
    END
    PORT
      LAYER li1 ;
        RECT 204.715 1762.750 204.885 1762.920 ;
        RECT 210.155 1762.750 210.325 1762.920 ;
      LAYER li1 ;
        RECT 210.155 1762.520 210.325 1762.605 ;
      LAYER li1 ;
        RECT 204.715 1762.290 204.885 1762.460 ;
        RECT 204.715 1761.830 204.885 1762.000 ;
        RECT 204.715 1761.370 204.885 1761.540 ;
        RECT 204.715 1760.910 204.885 1761.080 ;
        RECT 204.715 1760.450 204.885 1760.620 ;
        RECT 204.715 1759.990 204.885 1760.160 ;
        RECT 204.715 1759.530 204.885 1759.700 ;
        RECT 204.715 1759.070 204.885 1759.240 ;
      LAYER li1 ;
        RECT 209.720 1759.115 210.325 1762.520 ;
      LAYER li1 ;
        RECT 204.715 1758.610 204.885 1758.780 ;
      LAYER li1 ;
        RECT 208.470 1758.765 210.325 1759.115 ;
      LAYER li1 ;
        RECT 204.715 1758.150 204.885 1758.320 ;
        RECT 204.715 1757.690 204.885 1757.860 ;
        RECT 204.715 1757.230 204.885 1757.400 ;
      LAYER li1 ;
        RECT 209.720 1757.175 210.325 1758.765 ;
        RECT 210.155 1757.085 210.325 1757.175 ;
      LAYER li1 ;
        RECT 204.715 1756.770 204.885 1756.940 ;
        RECT 210.155 1756.770 210.325 1756.940 ;
      LAYER li1 ;
        RECT 210.155 1756.540 210.325 1756.625 ;
      LAYER li1 ;
        RECT 204.715 1756.310 204.885 1756.480 ;
        RECT 204.715 1755.850 204.885 1756.020 ;
        RECT 204.715 1755.390 204.885 1755.560 ;
        RECT 204.715 1754.930 204.885 1755.100 ;
        RECT 204.715 1754.470 204.885 1754.640 ;
        RECT 204.715 1754.010 204.885 1754.180 ;
        RECT 204.715 1753.550 204.885 1753.720 ;
        RECT 204.715 1753.090 204.885 1753.260 ;
      LAYER li1 ;
        RECT 209.720 1753.135 210.325 1756.540 ;
      LAYER li1 ;
        RECT 204.715 1752.630 204.885 1752.800 ;
      LAYER li1 ;
        RECT 208.470 1752.785 210.325 1753.135 ;
      LAYER li1 ;
        RECT 204.715 1752.170 204.885 1752.340 ;
        RECT 204.715 1751.710 204.885 1751.880 ;
        RECT 204.715 1751.250 204.885 1751.420 ;
      LAYER li1 ;
        RECT 209.720 1751.195 210.325 1752.785 ;
        RECT 210.155 1751.105 210.325 1751.195 ;
      LAYER li1 ;
        RECT 204.715 1750.790 204.885 1750.960 ;
        RECT 210.155 1750.790 210.325 1750.960 ;
        RECT 204.715 1750.330 204.885 1750.500 ;
        RECT 210.155 1750.330 210.325 1750.500 ;
        RECT 204.715 1749.870 204.885 1750.040 ;
        RECT 210.155 1749.870 210.325 1750.040 ;
        RECT 204.715 1749.410 204.885 1749.580 ;
        RECT 210.155 1749.410 210.325 1749.580 ;
        RECT 204.715 1748.950 204.885 1749.120 ;
        RECT 210.155 1748.950 210.325 1749.120 ;
        RECT 204.715 1748.490 204.885 1748.660 ;
        RECT 210.155 1748.490 210.325 1748.660 ;
        RECT 204.715 1748.030 204.885 1748.200 ;
        RECT 210.155 1748.030 210.325 1748.200 ;
        RECT 204.715 1747.570 204.885 1747.740 ;
        RECT 210.155 1747.570 210.325 1747.740 ;
        RECT 204.715 1747.110 204.885 1747.280 ;
        RECT 210.155 1747.110 210.325 1747.280 ;
        RECT 204.715 1746.650 204.885 1746.820 ;
        RECT 210.155 1746.650 210.325 1746.820 ;
        RECT 204.715 1746.190 204.885 1746.360 ;
        RECT 210.155 1746.190 210.325 1746.360 ;
        RECT 204.715 1745.730 204.885 1745.900 ;
        RECT 210.155 1745.730 210.325 1745.900 ;
        RECT 204.715 1745.270 204.885 1745.440 ;
        RECT 210.155 1745.270 210.325 1745.440 ;
        RECT 204.715 1744.810 204.885 1744.980 ;
        RECT 210.155 1744.810 210.325 1744.980 ;
      LAYER li1 ;
        RECT 210.155 1744.580 210.325 1744.665 ;
      LAYER li1 ;
        RECT 204.715 1744.350 204.885 1744.520 ;
        RECT 204.715 1743.890 204.885 1744.060 ;
        RECT 204.715 1743.430 204.885 1743.600 ;
        RECT 204.715 1742.970 204.885 1743.140 ;
        RECT 204.715 1742.510 204.885 1742.680 ;
        RECT 204.715 1742.050 204.885 1742.220 ;
        RECT 204.715 1741.590 204.885 1741.760 ;
        RECT 204.715 1741.130 204.885 1741.300 ;
      LAYER li1 ;
        RECT 209.720 1741.175 210.325 1744.580 ;
      LAYER li1 ;
        RECT 204.715 1740.670 204.885 1740.840 ;
      LAYER li1 ;
        RECT 208.470 1740.825 210.325 1741.175 ;
      LAYER li1 ;
        RECT 204.715 1740.210 204.885 1740.380 ;
        RECT 204.715 1739.750 204.885 1739.920 ;
        RECT 204.715 1739.290 204.885 1739.460 ;
      LAYER li1 ;
        RECT 209.720 1739.235 210.325 1740.825 ;
        RECT 210.155 1739.145 210.325 1739.235 ;
      LAYER li1 ;
        RECT 204.715 1738.830 204.885 1739.000 ;
        RECT 210.155 1738.830 210.325 1739.000 ;
      LAYER li1 ;
        RECT 210.155 1738.600 210.325 1738.685 ;
      LAYER li1 ;
        RECT 204.715 1738.370 204.885 1738.540 ;
        RECT 204.715 1737.910 204.885 1738.080 ;
        RECT 204.715 1737.450 204.885 1737.620 ;
        RECT 204.715 1736.990 204.885 1737.160 ;
        RECT 204.715 1736.530 204.885 1736.700 ;
        RECT 204.715 1736.070 204.885 1736.240 ;
        RECT 204.715 1735.610 204.885 1735.780 ;
        RECT 204.715 1735.150 204.885 1735.320 ;
      LAYER li1 ;
        RECT 209.720 1735.195 210.325 1738.600 ;
      LAYER li1 ;
        RECT 204.715 1734.690 204.885 1734.860 ;
      LAYER li1 ;
        RECT 208.470 1734.845 210.325 1735.195 ;
      LAYER li1 ;
        RECT 204.715 1734.230 204.885 1734.400 ;
        RECT 204.715 1733.770 204.885 1733.940 ;
        RECT 204.715 1733.310 204.885 1733.480 ;
      LAYER li1 ;
        RECT 209.720 1733.255 210.325 1734.845 ;
        RECT 210.155 1733.165 210.325 1733.255 ;
      LAYER li1 ;
        RECT 204.715 1732.850 204.885 1733.020 ;
        RECT 210.155 1732.850 210.325 1733.020 ;
      LAYER li1 ;
        RECT 210.155 1732.620 210.325 1732.705 ;
      LAYER li1 ;
        RECT 204.715 1732.390 204.885 1732.560 ;
        RECT 204.715 1731.930 204.885 1732.100 ;
        RECT 204.715 1731.470 204.885 1731.640 ;
        RECT 204.715 1731.010 204.885 1731.180 ;
        RECT 204.715 1730.550 204.885 1730.720 ;
        RECT 204.715 1730.090 204.885 1730.260 ;
        RECT 204.715 1729.630 204.885 1729.800 ;
        RECT 204.715 1729.170 204.885 1729.340 ;
      LAYER li1 ;
        RECT 209.720 1729.215 210.325 1732.620 ;
      LAYER li1 ;
        RECT 204.715 1728.710 204.885 1728.880 ;
      LAYER li1 ;
        RECT 208.470 1728.865 210.325 1729.215 ;
      LAYER li1 ;
        RECT 204.715 1728.250 204.885 1728.420 ;
        RECT 204.715 1727.790 204.885 1727.960 ;
        RECT 204.715 1727.330 204.885 1727.500 ;
      LAYER li1 ;
        RECT 209.720 1727.275 210.325 1728.865 ;
        RECT 210.155 1727.185 210.325 1727.275 ;
      LAYER li1 ;
        RECT 204.715 1726.870 204.885 1727.040 ;
        RECT 210.155 1726.870 210.325 1727.040 ;
      LAYER li1 ;
        RECT 210.155 1726.640 210.325 1726.725 ;
      LAYER li1 ;
        RECT 204.715 1726.410 204.885 1726.580 ;
        RECT 204.715 1725.950 204.885 1726.120 ;
        RECT 204.715 1725.490 204.885 1725.660 ;
        RECT 204.715 1725.030 204.885 1725.200 ;
        RECT 204.715 1724.570 204.885 1724.740 ;
        RECT 204.715 1724.110 204.885 1724.280 ;
        RECT 204.715 1723.650 204.885 1723.820 ;
        RECT 204.715 1723.190 204.885 1723.360 ;
      LAYER li1 ;
        RECT 209.720 1723.235 210.325 1726.640 ;
      LAYER li1 ;
        RECT 204.715 1722.730 204.885 1722.900 ;
      LAYER li1 ;
        RECT 208.470 1722.885 210.325 1723.235 ;
      LAYER li1 ;
        RECT 204.715 1722.270 204.885 1722.440 ;
        RECT 204.715 1721.810 204.885 1721.980 ;
        RECT 204.715 1721.350 204.885 1721.520 ;
      LAYER li1 ;
        RECT 209.720 1721.295 210.325 1722.885 ;
        RECT 210.155 1721.205 210.325 1721.295 ;
      LAYER li1 ;
        RECT 204.715 1720.890 204.885 1721.060 ;
        RECT 210.155 1720.890 210.325 1721.060 ;
      LAYER li1 ;
        RECT 210.155 1720.660 210.325 1720.745 ;
      LAYER li1 ;
        RECT 204.715 1720.430 204.885 1720.600 ;
        RECT 204.715 1719.970 204.885 1720.140 ;
        RECT 204.715 1719.510 204.885 1719.680 ;
        RECT 204.715 1719.050 204.885 1719.220 ;
        RECT 204.715 1718.590 204.885 1718.760 ;
        RECT 204.715 1718.130 204.885 1718.300 ;
        RECT 204.715 1717.670 204.885 1717.840 ;
        RECT 204.715 1717.210 204.885 1717.380 ;
      LAYER li1 ;
        RECT 209.720 1717.255 210.325 1720.660 ;
      LAYER li1 ;
        RECT 204.715 1716.750 204.885 1716.920 ;
      LAYER li1 ;
        RECT 208.470 1716.905 210.325 1717.255 ;
      LAYER li1 ;
        RECT 204.715 1716.290 204.885 1716.460 ;
        RECT 204.715 1715.830 204.885 1716.000 ;
        RECT 204.715 1715.370 204.885 1715.540 ;
      LAYER li1 ;
        RECT 209.720 1715.315 210.325 1716.905 ;
        RECT 210.155 1715.225 210.325 1715.315 ;
      LAYER li1 ;
        RECT 204.715 1714.910 204.885 1715.080 ;
        RECT 210.155 1714.910 210.325 1715.080 ;
      LAYER li1 ;
        RECT 210.155 1714.680 210.325 1714.765 ;
      LAYER li1 ;
        RECT 204.715 1714.450 204.885 1714.620 ;
        RECT 204.715 1713.990 204.885 1714.160 ;
        RECT 204.715 1713.530 204.885 1713.700 ;
        RECT 204.715 1713.070 204.885 1713.240 ;
        RECT 204.715 1712.610 204.885 1712.780 ;
        RECT 204.715 1712.150 204.885 1712.320 ;
        RECT 204.715 1711.690 204.885 1711.860 ;
        RECT 204.715 1711.230 204.885 1711.400 ;
      LAYER li1 ;
        RECT 209.720 1711.275 210.325 1714.680 ;
      LAYER li1 ;
        RECT 204.715 1710.770 204.885 1710.940 ;
      LAYER li1 ;
        RECT 208.470 1710.925 210.325 1711.275 ;
      LAYER li1 ;
        RECT 204.715 1710.310 204.885 1710.480 ;
        RECT 204.715 1709.850 204.885 1710.020 ;
        RECT 204.715 1709.390 204.885 1709.560 ;
      LAYER li1 ;
        RECT 209.720 1709.335 210.325 1710.925 ;
        RECT 210.155 1709.245 210.325 1709.335 ;
      LAYER li1 ;
        RECT 204.715 1708.930 204.885 1709.100 ;
        RECT 210.155 1708.930 210.325 1709.100 ;
      LAYER li1 ;
        RECT 210.155 1708.700 210.325 1708.785 ;
      LAYER li1 ;
        RECT 204.715 1708.470 204.885 1708.640 ;
        RECT 204.715 1708.010 204.885 1708.180 ;
        RECT 204.715 1707.550 204.885 1707.720 ;
        RECT 204.715 1707.090 204.885 1707.260 ;
        RECT 204.715 1706.630 204.885 1706.800 ;
        RECT 204.715 1706.170 204.885 1706.340 ;
        RECT 204.715 1705.710 204.885 1705.880 ;
        RECT 204.715 1705.250 204.885 1705.420 ;
      LAYER li1 ;
        RECT 209.720 1705.295 210.325 1708.700 ;
      LAYER li1 ;
        RECT 204.715 1704.790 204.885 1704.960 ;
      LAYER li1 ;
        RECT 208.470 1704.945 210.325 1705.295 ;
      LAYER li1 ;
        RECT 204.715 1704.330 204.885 1704.500 ;
        RECT 204.715 1703.870 204.885 1704.040 ;
        RECT 204.715 1703.410 204.885 1703.580 ;
      LAYER li1 ;
        RECT 209.720 1703.355 210.325 1704.945 ;
        RECT 210.155 1703.265 210.325 1703.355 ;
      LAYER li1 ;
        RECT 204.715 1702.950 204.885 1703.120 ;
        RECT 210.155 1702.950 210.325 1703.120 ;
      LAYER li1 ;
        RECT 210.155 1702.720 210.325 1702.805 ;
      LAYER li1 ;
        RECT 204.715 1702.490 204.885 1702.660 ;
        RECT 204.715 1702.030 204.885 1702.200 ;
        RECT 204.715 1701.570 204.885 1701.740 ;
        RECT 204.715 1701.110 204.885 1701.280 ;
        RECT 204.715 1700.650 204.885 1700.820 ;
        RECT 204.715 1700.190 204.885 1700.360 ;
        RECT 204.715 1699.730 204.885 1699.900 ;
        RECT 204.715 1699.270 204.885 1699.440 ;
      LAYER li1 ;
        RECT 209.720 1699.315 210.325 1702.720 ;
      LAYER li1 ;
        RECT 204.715 1698.810 204.885 1698.980 ;
      LAYER li1 ;
        RECT 208.470 1698.965 210.325 1699.315 ;
      LAYER li1 ;
        RECT 204.715 1698.350 204.885 1698.520 ;
        RECT 204.715 1697.890 204.885 1698.060 ;
        RECT 204.715 1697.430 204.885 1697.600 ;
      LAYER li1 ;
        RECT 209.720 1697.375 210.325 1698.965 ;
        RECT 210.155 1697.285 210.325 1697.375 ;
      LAYER li1 ;
        RECT 204.715 1696.970 204.885 1697.140 ;
        RECT 210.155 1696.970 210.325 1697.140 ;
      LAYER li1 ;
        RECT 210.155 1696.740 210.325 1696.825 ;
      LAYER li1 ;
        RECT 204.715 1696.510 204.885 1696.680 ;
        RECT 204.715 1696.050 204.885 1696.220 ;
        RECT 204.715 1695.590 204.885 1695.760 ;
        RECT 204.715 1695.130 204.885 1695.300 ;
        RECT 204.715 1694.670 204.885 1694.840 ;
        RECT 204.715 1694.210 204.885 1694.380 ;
        RECT 204.715 1693.750 204.885 1693.920 ;
        RECT 204.715 1693.290 204.885 1693.460 ;
      LAYER li1 ;
        RECT 209.720 1693.335 210.325 1696.740 ;
      LAYER li1 ;
        RECT 204.715 1692.830 204.885 1693.000 ;
      LAYER li1 ;
        RECT 208.470 1692.985 210.325 1693.335 ;
      LAYER li1 ;
        RECT 204.715 1692.370 204.885 1692.540 ;
        RECT 204.715 1691.910 204.885 1692.080 ;
        RECT 204.715 1691.450 204.885 1691.620 ;
      LAYER li1 ;
        RECT 209.720 1691.395 210.325 1692.985 ;
        RECT 210.155 1691.305 210.325 1691.395 ;
      LAYER li1 ;
        RECT 204.715 1690.990 204.885 1691.160 ;
        RECT 210.155 1690.990 210.325 1691.160 ;
      LAYER li1 ;
        RECT 210.155 1690.760 210.325 1690.845 ;
      LAYER li1 ;
        RECT 204.715 1690.530 204.885 1690.700 ;
        RECT 204.715 1690.070 204.885 1690.240 ;
        RECT 204.715 1689.610 204.885 1689.780 ;
        RECT 204.715 1689.150 204.885 1689.320 ;
        RECT 204.715 1688.690 204.885 1688.860 ;
        RECT 204.715 1688.230 204.885 1688.400 ;
        RECT 204.715 1687.770 204.885 1687.940 ;
        RECT 204.715 1687.310 204.885 1687.480 ;
      LAYER li1 ;
        RECT 209.720 1687.355 210.325 1690.760 ;
      LAYER li1 ;
        RECT 204.715 1686.850 204.885 1687.020 ;
      LAYER li1 ;
        RECT 208.470 1687.005 210.325 1687.355 ;
      LAYER li1 ;
        RECT 204.715 1686.390 204.885 1686.560 ;
        RECT 204.715 1685.930 204.885 1686.100 ;
        RECT 204.715 1685.470 204.885 1685.640 ;
      LAYER li1 ;
        RECT 209.720 1685.415 210.325 1687.005 ;
        RECT 210.155 1685.325 210.325 1685.415 ;
      LAYER li1 ;
        RECT 204.715 1685.010 204.885 1685.180 ;
        RECT 210.155 1685.010 210.325 1685.180 ;
      LAYER li1 ;
        RECT 210.155 1684.780 210.325 1684.865 ;
      LAYER li1 ;
        RECT 204.715 1684.550 204.885 1684.720 ;
        RECT 204.715 1684.090 204.885 1684.260 ;
        RECT 204.715 1683.630 204.885 1683.800 ;
        RECT 204.715 1683.170 204.885 1683.340 ;
        RECT 204.715 1682.710 204.885 1682.880 ;
        RECT 204.715 1682.250 204.885 1682.420 ;
        RECT 204.715 1681.790 204.885 1681.960 ;
        RECT 204.715 1681.330 204.885 1681.500 ;
      LAYER li1 ;
        RECT 209.720 1681.375 210.325 1684.780 ;
      LAYER li1 ;
        RECT 204.715 1680.870 204.885 1681.040 ;
      LAYER li1 ;
        RECT 208.470 1681.025 210.325 1681.375 ;
      LAYER li1 ;
        RECT 204.715 1680.410 204.885 1680.580 ;
        RECT 204.715 1679.950 204.885 1680.120 ;
        RECT 204.715 1679.490 204.885 1679.660 ;
      LAYER li1 ;
        RECT 209.720 1679.435 210.325 1681.025 ;
        RECT 210.155 1679.345 210.325 1679.435 ;
      LAYER li1 ;
        RECT 204.715 1679.030 204.885 1679.200 ;
        RECT 210.155 1679.030 210.325 1679.200 ;
      LAYER li1 ;
        RECT 210.155 1678.800 210.325 1678.885 ;
      LAYER li1 ;
        RECT 204.715 1678.570 204.885 1678.740 ;
        RECT 204.715 1678.110 204.885 1678.280 ;
        RECT 204.715 1677.650 204.885 1677.820 ;
        RECT 204.715 1677.190 204.885 1677.360 ;
        RECT 204.715 1676.730 204.885 1676.900 ;
        RECT 204.715 1676.270 204.885 1676.440 ;
        RECT 204.715 1675.810 204.885 1675.980 ;
        RECT 204.715 1675.350 204.885 1675.520 ;
      LAYER li1 ;
        RECT 209.720 1675.395 210.325 1678.800 ;
      LAYER li1 ;
        RECT 204.715 1674.890 204.885 1675.060 ;
      LAYER li1 ;
        RECT 208.470 1675.045 210.325 1675.395 ;
      LAYER li1 ;
        RECT 204.715 1674.430 204.885 1674.600 ;
        RECT 204.715 1673.970 204.885 1674.140 ;
        RECT 204.715 1673.510 204.885 1673.680 ;
      LAYER li1 ;
        RECT 209.720 1673.455 210.325 1675.045 ;
        RECT 210.155 1673.365 210.325 1673.455 ;
      LAYER li1 ;
        RECT 204.715 1673.050 204.885 1673.220 ;
        RECT 210.155 1673.050 210.325 1673.220 ;
      LAYER mcon ;
        RECT 210.155 1761.830 210.325 1762.000 ;
        RECT 210.155 1761.370 210.325 1761.540 ;
        RECT 210.155 1760.910 210.325 1761.080 ;
        RECT 210.155 1760.450 210.325 1760.620 ;
        RECT 210.155 1759.990 210.325 1760.160 ;
        RECT 210.155 1759.530 210.325 1759.700 ;
        RECT 210.155 1759.070 210.325 1759.240 ;
        RECT 210.155 1758.610 210.325 1758.780 ;
        RECT 210.155 1758.150 210.325 1758.320 ;
        RECT 210.155 1757.690 210.325 1757.860 ;
        RECT 210.155 1757.230 210.325 1757.400 ;
        RECT 210.155 1755.850 210.325 1756.020 ;
        RECT 210.155 1755.390 210.325 1755.560 ;
        RECT 210.155 1754.930 210.325 1755.100 ;
        RECT 210.155 1754.470 210.325 1754.640 ;
        RECT 210.155 1754.010 210.325 1754.180 ;
        RECT 210.155 1753.550 210.325 1753.720 ;
        RECT 210.155 1753.090 210.325 1753.260 ;
        RECT 210.155 1752.630 210.325 1752.800 ;
        RECT 210.155 1752.170 210.325 1752.340 ;
        RECT 210.155 1751.710 210.325 1751.880 ;
        RECT 210.155 1751.250 210.325 1751.420 ;
        RECT 210.155 1743.890 210.325 1744.060 ;
        RECT 210.155 1743.430 210.325 1743.600 ;
        RECT 210.155 1742.970 210.325 1743.140 ;
        RECT 210.155 1742.510 210.325 1742.680 ;
        RECT 210.155 1742.050 210.325 1742.220 ;
        RECT 210.155 1741.590 210.325 1741.760 ;
        RECT 210.155 1741.130 210.325 1741.300 ;
        RECT 210.155 1740.670 210.325 1740.840 ;
        RECT 210.155 1740.210 210.325 1740.380 ;
        RECT 210.155 1739.750 210.325 1739.920 ;
        RECT 210.155 1739.290 210.325 1739.460 ;
        RECT 210.155 1737.910 210.325 1738.080 ;
        RECT 210.155 1737.450 210.325 1737.620 ;
        RECT 210.155 1736.990 210.325 1737.160 ;
        RECT 210.155 1736.530 210.325 1736.700 ;
        RECT 210.155 1736.070 210.325 1736.240 ;
        RECT 210.155 1735.610 210.325 1735.780 ;
        RECT 210.155 1735.150 210.325 1735.320 ;
        RECT 210.155 1734.690 210.325 1734.860 ;
        RECT 210.155 1734.230 210.325 1734.400 ;
        RECT 210.155 1733.770 210.325 1733.940 ;
        RECT 210.155 1733.310 210.325 1733.480 ;
        RECT 210.155 1731.930 210.325 1732.100 ;
        RECT 210.155 1731.470 210.325 1731.640 ;
        RECT 210.155 1731.010 210.325 1731.180 ;
        RECT 210.155 1730.550 210.325 1730.720 ;
        RECT 210.155 1730.090 210.325 1730.260 ;
        RECT 210.155 1729.630 210.325 1729.800 ;
        RECT 210.155 1729.170 210.325 1729.340 ;
        RECT 210.155 1728.710 210.325 1728.880 ;
        RECT 210.155 1728.250 210.325 1728.420 ;
        RECT 210.155 1727.790 210.325 1727.960 ;
        RECT 210.155 1727.330 210.325 1727.500 ;
        RECT 210.155 1725.950 210.325 1726.120 ;
        RECT 210.155 1725.490 210.325 1725.660 ;
        RECT 210.155 1725.030 210.325 1725.200 ;
        RECT 210.155 1724.570 210.325 1724.740 ;
        RECT 210.155 1724.110 210.325 1724.280 ;
        RECT 210.155 1723.650 210.325 1723.820 ;
        RECT 210.155 1723.190 210.325 1723.360 ;
        RECT 210.155 1722.730 210.325 1722.900 ;
        RECT 210.155 1722.270 210.325 1722.440 ;
        RECT 210.155 1721.810 210.325 1721.980 ;
        RECT 210.155 1721.350 210.325 1721.520 ;
        RECT 210.155 1719.970 210.325 1720.140 ;
        RECT 210.155 1719.510 210.325 1719.680 ;
        RECT 210.155 1719.050 210.325 1719.220 ;
        RECT 210.155 1718.590 210.325 1718.760 ;
        RECT 210.155 1718.130 210.325 1718.300 ;
        RECT 210.155 1717.670 210.325 1717.840 ;
        RECT 210.155 1717.210 210.325 1717.380 ;
        RECT 210.155 1716.750 210.325 1716.920 ;
        RECT 210.155 1716.290 210.325 1716.460 ;
        RECT 210.155 1715.830 210.325 1716.000 ;
        RECT 210.155 1715.370 210.325 1715.540 ;
        RECT 210.155 1713.990 210.325 1714.160 ;
        RECT 210.155 1713.530 210.325 1713.700 ;
        RECT 210.155 1713.070 210.325 1713.240 ;
        RECT 210.155 1712.610 210.325 1712.780 ;
        RECT 210.155 1712.150 210.325 1712.320 ;
        RECT 210.155 1711.690 210.325 1711.860 ;
        RECT 210.155 1711.230 210.325 1711.400 ;
        RECT 210.155 1710.770 210.325 1710.940 ;
        RECT 210.155 1710.310 210.325 1710.480 ;
        RECT 210.155 1709.850 210.325 1710.020 ;
        RECT 210.155 1709.390 210.325 1709.560 ;
        RECT 210.155 1708.010 210.325 1708.180 ;
        RECT 210.155 1707.550 210.325 1707.720 ;
        RECT 210.155 1707.090 210.325 1707.260 ;
        RECT 210.155 1706.630 210.325 1706.800 ;
        RECT 210.155 1706.170 210.325 1706.340 ;
        RECT 210.155 1705.710 210.325 1705.880 ;
        RECT 210.155 1705.250 210.325 1705.420 ;
        RECT 210.155 1704.790 210.325 1704.960 ;
        RECT 210.155 1704.330 210.325 1704.500 ;
        RECT 210.155 1703.870 210.325 1704.040 ;
        RECT 210.155 1703.410 210.325 1703.580 ;
        RECT 210.155 1702.030 210.325 1702.200 ;
        RECT 210.155 1701.570 210.325 1701.740 ;
        RECT 210.155 1701.110 210.325 1701.280 ;
        RECT 210.155 1700.650 210.325 1700.820 ;
        RECT 210.155 1700.190 210.325 1700.360 ;
        RECT 210.155 1699.730 210.325 1699.900 ;
        RECT 210.155 1699.270 210.325 1699.440 ;
        RECT 210.155 1698.810 210.325 1698.980 ;
        RECT 210.155 1698.350 210.325 1698.520 ;
        RECT 210.155 1697.890 210.325 1698.060 ;
        RECT 210.155 1697.430 210.325 1697.600 ;
        RECT 210.155 1696.050 210.325 1696.220 ;
        RECT 210.155 1695.590 210.325 1695.760 ;
        RECT 210.155 1695.130 210.325 1695.300 ;
        RECT 210.155 1694.670 210.325 1694.840 ;
        RECT 210.155 1694.210 210.325 1694.380 ;
        RECT 210.155 1693.750 210.325 1693.920 ;
        RECT 210.155 1693.290 210.325 1693.460 ;
        RECT 210.155 1692.830 210.325 1693.000 ;
        RECT 210.155 1692.370 210.325 1692.540 ;
        RECT 210.155 1691.910 210.325 1692.080 ;
        RECT 210.155 1691.450 210.325 1691.620 ;
        RECT 210.155 1690.070 210.325 1690.240 ;
        RECT 210.155 1689.610 210.325 1689.780 ;
        RECT 210.155 1689.150 210.325 1689.320 ;
        RECT 210.155 1688.690 210.325 1688.860 ;
        RECT 210.155 1688.230 210.325 1688.400 ;
        RECT 210.155 1687.770 210.325 1687.940 ;
        RECT 210.155 1687.310 210.325 1687.480 ;
        RECT 210.155 1686.850 210.325 1687.020 ;
        RECT 210.155 1686.390 210.325 1686.560 ;
        RECT 210.155 1685.930 210.325 1686.100 ;
        RECT 210.155 1685.470 210.325 1685.640 ;
        RECT 210.155 1684.090 210.325 1684.260 ;
        RECT 210.155 1683.630 210.325 1683.800 ;
        RECT 210.155 1683.170 210.325 1683.340 ;
        RECT 210.155 1682.710 210.325 1682.880 ;
        RECT 210.155 1682.250 210.325 1682.420 ;
        RECT 210.155 1681.790 210.325 1681.960 ;
        RECT 210.155 1681.330 210.325 1681.500 ;
        RECT 210.155 1680.870 210.325 1681.040 ;
        RECT 210.155 1680.410 210.325 1680.580 ;
        RECT 210.155 1679.950 210.325 1680.120 ;
        RECT 210.155 1679.490 210.325 1679.660 ;
        RECT 210.155 1678.110 210.325 1678.280 ;
        RECT 210.155 1677.650 210.325 1677.820 ;
        RECT 210.155 1677.190 210.325 1677.360 ;
        RECT 210.155 1676.730 210.325 1676.900 ;
        RECT 210.155 1676.270 210.325 1676.440 ;
        RECT 210.155 1675.810 210.325 1675.980 ;
        RECT 210.155 1675.350 210.325 1675.520 ;
        RECT 210.155 1674.890 210.325 1675.060 ;
        RECT 210.155 1674.430 210.325 1674.600 ;
        RECT 210.155 1673.970 210.325 1674.140 ;
        RECT 210.155 1673.510 210.325 1673.680 ;
      LAYER met1 ;
        RECT 204.560 1672.905 205.040 1763.065 ;
        RECT 210.000 1672.905 210.480 1763.065 ;
      LAYER via ;
        RECT 204.655 1728.815 204.955 1730.600 ;
        RECT 210.095 1728.815 210.395 1730.600 ;
      LAYER met2 ;
        RECT 204.595 1728.775 205.025 1730.640 ;
        RECT 210.035 1728.775 210.465 1730.640 ;
      LAYER via2 ;
        RECT 204.655 1728.815 204.955 1730.600 ;
        RECT 210.095 1728.815 210.395 1730.600 ;
      LAYER met3 ;
        RECT 200.210 1728.780 210.465 1730.630 ;
    END
    PORT
      LAYER li1 ;
        RECT 204.605 3050.655 204.775 3050.825 ;
        RECT 210.045 3050.655 210.215 3050.825 ;
      LAYER li1 ;
        RECT 210.045 3050.425 210.215 3050.510 ;
      LAYER li1 ;
        RECT 204.605 3050.195 204.775 3050.365 ;
        RECT 204.605 3049.735 204.775 3049.905 ;
        RECT 204.605 3049.275 204.775 3049.445 ;
        RECT 204.605 3048.815 204.775 3048.985 ;
        RECT 204.605 3048.355 204.775 3048.525 ;
        RECT 204.605 3047.895 204.775 3048.065 ;
        RECT 204.605 3047.435 204.775 3047.605 ;
        RECT 204.605 3046.975 204.775 3047.145 ;
      LAYER li1 ;
        RECT 209.610 3047.020 210.215 3050.425 ;
      LAYER li1 ;
        RECT 204.605 3046.515 204.775 3046.685 ;
      LAYER li1 ;
        RECT 208.360 3046.670 210.215 3047.020 ;
      LAYER li1 ;
        RECT 204.605 3046.055 204.775 3046.225 ;
        RECT 204.605 3045.595 204.775 3045.765 ;
        RECT 204.605 3045.135 204.775 3045.305 ;
      LAYER li1 ;
        RECT 209.610 3045.080 210.215 3046.670 ;
        RECT 210.045 3044.990 210.215 3045.080 ;
      LAYER li1 ;
        RECT 204.605 3044.675 204.775 3044.845 ;
        RECT 210.045 3044.675 210.215 3044.845 ;
      LAYER li1 ;
        RECT 210.045 3044.445 210.215 3044.530 ;
      LAYER li1 ;
        RECT 204.605 3044.215 204.775 3044.385 ;
        RECT 204.605 3043.755 204.775 3043.925 ;
        RECT 204.605 3043.295 204.775 3043.465 ;
        RECT 204.605 3042.835 204.775 3043.005 ;
        RECT 204.605 3042.375 204.775 3042.545 ;
        RECT 204.605 3041.915 204.775 3042.085 ;
        RECT 204.605 3041.455 204.775 3041.625 ;
        RECT 204.605 3040.995 204.775 3041.165 ;
      LAYER li1 ;
        RECT 209.610 3041.040 210.215 3044.445 ;
      LAYER li1 ;
        RECT 204.605 3040.535 204.775 3040.705 ;
      LAYER li1 ;
        RECT 208.360 3040.690 210.215 3041.040 ;
      LAYER li1 ;
        RECT 204.605 3040.075 204.775 3040.245 ;
        RECT 204.605 3039.615 204.775 3039.785 ;
        RECT 204.605 3039.155 204.775 3039.325 ;
      LAYER li1 ;
        RECT 209.610 3039.100 210.215 3040.690 ;
        RECT 210.045 3039.010 210.215 3039.100 ;
      LAYER li1 ;
        RECT 204.605 3038.695 204.775 3038.865 ;
        RECT 210.045 3038.695 210.215 3038.865 ;
      LAYER li1 ;
        RECT 210.045 3038.465 210.215 3038.550 ;
      LAYER li1 ;
        RECT 204.605 3038.235 204.775 3038.405 ;
        RECT 204.605 3037.775 204.775 3037.945 ;
        RECT 204.605 3037.315 204.775 3037.485 ;
        RECT 204.605 3036.855 204.775 3037.025 ;
        RECT 204.605 3036.395 204.775 3036.565 ;
        RECT 204.605 3035.935 204.775 3036.105 ;
        RECT 204.605 3035.475 204.775 3035.645 ;
        RECT 204.605 3035.015 204.775 3035.185 ;
      LAYER li1 ;
        RECT 209.610 3035.060 210.215 3038.465 ;
      LAYER li1 ;
        RECT 204.605 3034.555 204.775 3034.725 ;
      LAYER li1 ;
        RECT 208.360 3034.710 210.215 3035.060 ;
      LAYER li1 ;
        RECT 204.605 3034.095 204.775 3034.265 ;
        RECT 204.605 3033.635 204.775 3033.805 ;
        RECT 204.605 3033.175 204.775 3033.345 ;
      LAYER li1 ;
        RECT 209.610 3033.120 210.215 3034.710 ;
        RECT 210.045 3033.030 210.215 3033.120 ;
      LAYER li1 ;
        RECT 204.605 3032.715 204.775 3032.885 ;
        RECT 210.045 3032.715 210.215 3032.885 ;
      LAYER li1 ;
        RECT 210.045 3032.485 210.215 3032.570 ;
      LAYER li1 ;
        RECT 204.605 3032.255 204.775 3032.425 ;
        RECT 204.605 3031.795 204.775 3031.965 ;
        RECT 204.605 3031.335 204.775 3031.505 ;
        RECT 204.605 3030.875 204.775 3031.045 ;
        RECT 204.605 3030.415 204.775 3030.585 ;
        RECT 204.605 3029.955 204.775 3030.125 ;
        RECT 204.605 3029.495 204.775 3029.665 ;
        RECT 204.605 3029.035 204.775 3029.205 ;
      LAYER li1 ;
        RECT 209.610 3029.080 210.215 3032.485 ;
      LAYER li1 ;
        RECT 204.605 3028.575 204.775 3028.745 ;
      LAYER li1 ;
        RECT 208.360 3028.730 210.215 3029.080 ;
      LAYER li1 ;
        RECT 204.605 3028.115 204.775 3028.285 ;
        RECT 204.605 3027.655 204.775 3027.825 ;
        RECT 204.605 3027.195 204.775 3027.365 ;
      LAYER li1 ;
        RECT 209.610 3027.140 210.215 3028.730 ;
        RECT 210.045 3027.050 210.215 3027.140 ;
      LAYER li1 ;
        RECT 204.605 3026.735 204.775 3026.905 ;
        RECT 210.045 3026.735 210.215 3026.905 ;
      LAYER li1 ;
        RECT 210.045 3026.505 210.215 3026.590 ;
      LAYER li1 ;
        RECT 204.605 3026.275 204.775 3026.445 ;
        RECT 204.605 3025.815 204.775 3025.985 ;
        RECT 204.605 3025.355 204.775 3025.525 ;
        RECT 204.605 3024.895 204.775 3025.065 ;
        RECT 204.605 3024.435 204.775 3024.605 ;
        RECT 204.605 3023.975 204.775 3024.145 ;
        RECT 204.605 3023.515 204.775 3023.685 ;
        RECT 204.605 3023.055 204.775 3023.225 ;
      LAYER li1 ;
        RECT 209.610 3023.100 210.215 3026.505 ;
      LAYER li1 ;
        RECT 204.605 3022.595 204.775 3022.765 ;
      LAYER li1 ;
        RECT 208.360 3022.750 210.215 3023.100 ;
      LAYER li1 ;
        RECT 204.605 3022.135 204.775 3022.305 ;
        RECT 204.605 3021.675 204.775 3021.845 ;
        RECT 204.605 3021.215 204.775 3021.385 ;
      LAYER li1 ;
        RECT 209.610 3021.160 210.215 3022.750 ;
        RECT 210.045 3021.070 210.215 3021.160 ;
      LAYER li1 ;
        RECT 204.605 3020.755 204.775 3020.925 ;
        RECT 210.045 3020.755 210.215 3020.925 ;
      LAYER li1 ;
        RECT 210.045 3020.525 210.215 3020.610 ;
      LAYER li1 ;
        RECT 204.605 3020.295 204.775 3020.465 ;
        RECT 204.605 3019.835 204.775 3020.005 ;
        RECT 204.605 3019.375 204.775 3019.545 ;
        RECT 204.605 3018.915 204.775 3019.085 ;
        RECT 204.605 3018.455 204.775 3018.625 ;
        RECT 204.605 3017.995 204.775 3018.165 ;
        RECT 204.605 3017.535 204.775 3017.705 ;
        RECT 204.605 3017.075 204.775 3017.245 ;
      LAYER li1 ;
        RECT 209.610 3017.120 210.215 3020.525 ;
      LAYER li1 ;
        RECT 204.605 3016.615 204.775 3016.785 ;
      LAYER li1 ;
        RECT 208.360 3016.770 210.215 3017.120 ;
      LAYER li1 ;
        RECT 204.605 3016.155 204.775 3016.325 ;
        RECT 204.605 3015.695 204.775 3015.865 ;
        RECT 204.605 3015.235 204.775 3015.405 ;
      LAYER li1 ;
        RECT 209.610 3015.180 210.215 3016.770 ;
        RECT 210.045 3015.090 210.215 3015.180 ;
      LAYER li1 ;
        RECT 204.605 3014.775 204.775 3014.945 ;
        RECT 210.045 3014.775 210.215 3014.945 ;
      LAYER li1 ;
        RECT 210.045 3014.545 210.215 3014.630 ;
      LAYER li1 ;
        RECT 204.605 3014.315 204.775 3014.485 ;
        RECT 204.605 3013.855 204.775 3014.025 ;
        RECT 204.605 3013.395 204.775 3013.565 ;
        RECT 204.605 3012.935 204.775 3013.105 ;
        RECT 204.605 3012.475 204.775 3012.645 ;
        RECT 204.605 3012.015 204.775 3012.185 ;
        RECT 204.605 3011.555 204.775 3011.725 ;
        RECT 204.605 3011.095 204.775 3011.265 ;
      LAYER li1 ;
        RECT 209.610 3011.140 210.215 3014.545 ;
      LAYER li1 ;
        RECT 204.605 3010.635 204.775 3010.805 ;
      LAYER li1 ;
        RECT 208.360 3010.790 210.215 3011.140 ;
      LAYER li1 ;
        RECT 204.605 3010.175 204.775 3010.345 ;
        RECT 204.605 3009.715 204.775 3009.885 ;
        RECT 204.605 3009.255 204.775 3009.425 ;
      LAYER li1 ;
        RECT 209.610 3009.200 210.215 3010.790 ;
        RECT 210.045 3009.110 210.215 3009.200 ;
      LAYER li1 ;
        RECT 204.605 3008.795 204.775 3008.965 ;
        RECT 210.045 3008.795 210.215 3008.965 ;
      LAYER li1 ;
        RECT 210.045 3008.565 210.215 3008.650 ;
      LAYER li1 ;
        RECT 204.605 3008.335 204.775 3008.505 ;
        RECT 204.605 3007.875 204.775 3008.045 ;
        RECT 204.605 3007.415 204.775 3007.585 ;
        RECT 204.605 3006.955 204.775 3007.125 ;
        RECT 204.605 3006.495 204.775 3006.665 ;
        RECT 204.605 3006.035 204.775 3006.205 ;
        RECT 204.605 3005.575 204.775 3005.745 ;
        RECT 204.605 3005.115 204.775 3005.285 ;
      LAYER li1 ;
        RECT 209.610 3005.160 210.215 3008.565 ;
      LAYER li1 ;
        RECT 204.605 3004.655 204.775 3004.825 ;
      LAYER li1 ;
        RECT 208.360 3004.810 210.215 3005.160 ;
      LAYER li1 ;
        RECT 204.605 3004.195 204.775 3004.365 ;
        RECT 204.605 3003.735 204.775 3003.905 ;
        RECT 204.605 3003.275 204.775 3003.445 ;
      LAYER li1 ;
        RECT 209.610 3003.220 210.215 3004.810 ;
        RECT 210.045 3003.130 210.215 3003.220 ;
      LAYER li1 ;
        RECT 204.605 3002.815 204.775 3002.985 ;
        RECT 210.045 3002.815 210.215 3002.985 ;
      LAYER li1 ;
        RECT 210.045 3002.585 210.215 3002.670 ;
      LAYER li1 ;
        RECT 204.605 3002.355 204.775 3002.525 ;
        RECT 204.605 3001.895 204.775 3002.065 ;
        RECT 204.605 3001.435 204.775 3001.605 ;
        RECT 204.605 3000.975 204.775 3001.145 ;
        RECT 204.605 3000.515 204.775 3000.685 ;
        RECT 204.605 3000.055 204.775 3000.225 ;
        RECT 204.605 2999.595 204.775 2999.765 ;
        RECT 204.605 2999.135 204.775 2999.305 ;
      LAYER li1 ;
        RECT 209.610 2999.180 210.215 3002.585 ;
      LAYER li1 ;
        RECT 204.605 2998.675 204.775 2998.845 ;
      LAYER li1 ;
        RECT 208.360 2998.830 210.215 2999.180 ;
      LAYER li1 ;
        RECT 204.605 2998.215 204.775 2998.385 ;
        RECT 204.605 2997.755 204.775 2997.925 ;
        RECT 204.605 2997.295 204.775 2997.465 ;
      LAYER li1 ;
        RECT 209.610 2997.240 210.215 2998.830 ;
        RECT 210.045 2997.150 210.215 2997.240 ;
      LAYER li1 ;
        RECT 204.605 2996.835 204.775 2997.005 ;
        RECT 210.045 2996.835 210.215 2997.005 ;
      LAYER li1 ;
        RECT 210.045 2996.605 210.215 2996.690 ;
      LAYER li1 ;
        RECT 204.605 2996.375 204.775 2996.545 ;
        RECT 204.605 2995.915 204.775 2996.085 ;
        RECT 204.605 2995.455 204.775 2995.625 ;
        RECT 204.605 2994.995 204.775 2995.165 ;
        RECT 204.605 2994.535 204.775 2994.705 ;
        RECT 204.605 2994.075 204.775 2994.245 ;
        RECT 204.605 2993.615 204.775 2993.785 ;
        RECT 204.605 2993.155 204.775 2993.325 ;
      LAYER li1 ;
        RECT 209.610 2993.200 210.215 2996.605 ;
      LAYER li1 ;
        RECT 204.605 2992.695 204.775 2992.865 ;
      LAYER li1 ;
        RECT 208.360 2992.850 210.215 2993.200 ;
      LAYER li1 ;
        RECT 204.605 2992.235 204.775 2992.405 ;
        RECT 204.605 2991.775 204.775 2991.945 ;
        RECT 204.605 2991.315 204.775 2991.485 ;
      LAYER li1 ;
        RECT 209.610 2991.260 210.215 2992.850 ;
        RECT 210.045 2991.170 210.215 2991.260 ;
      LAYER li1 ;
        RECT 204.605 2990.855 204.775 2991.025 ;
        RECT 210.045 2990.855 210.215 2991.025 ;
      LAYER li1 ;
        RECT 210.045 2990.625 210.215 2990.710 ;
      LAYER li1 ;
        RECT 204.605 2990.395 204.775 2990.565 ;
        RECT 204.605 2989.935 204.775 2990.105 ;
        RECT 204.605 2989.475 204.775 2989.645 ;
        RECT 204.605 2989.015 204.775 2989.185 ;
        RECT 204.605 2988.555 204.775 2988.725 ;
        RECT 204.605 2988.095 204.775 2988.265 ;
        RECT 204.605 2987.635 204.775 2987.805 ;
        RECT 204.605 2987.175 204.775 2987.345 ;
      LAYER li1 ;
        RECT 209.610 2987.220 210.215 2990.625 ;
      LAYER li1 ;
        RECT 204.605 2986.715 204.775 2986.885 ;
      LAYER li1 ;
        RECT 208.360 2986.870 210.215 2987.220 ;
      LAYER li1 ;
        RECT 204.605 2986.255 204.775 2986.425 ;
        RECT 204.605 2985.795 204.775 2985.965 ;
        RECT 204.605 2985.335 204.775 2985.505 ;
      LAYER li1 ;
        RECT 209.610 2985.280 210.215 2986.870 ;
        RECT 210.045 2985.190 210.215 2985.280 ;
      LAYER li1 ;
        RECT 204.605 2984.875 204.775 2985.045 ;
        RECT 210.045 2984.875 210.215 2985.045 ;
      LAYER mcon ;
        RECT 210.045 3049.735 210.215 3049.905 ;
        RECT 210.045 3049.275 210.215 3049.445 ;
        RECT 210.045 3048.815 210.215 3048.985 ;
        RECT 210.045 3048.355 210.215 3048.525 ;
        RECT 210.045 3047.895 210.215 3048.065 ;
        RECT 210.045 3047.435 210.215 3047.605 ;
        RECT 210.045 3046.975 210.215 3047.145 ;
        RECT 210.045 3046.515 210.215 3046.685 ;
        RECT 210.045 3046.055 210.215 3046.225 ;
        RECT 210.045 3045.595 210.215 3045.765 ;
        RECT 210.045 3045.135 210.215 3045.305 ;
        RECT 210.045 3043.755 210.215 3043.925 ;
        RECT 210.045 3043.295 210.215 3043.465 ;
        RECT 210.045 3042.835 210.215 3043.005 ;
        RECT 210.045 3042.375 210.215 3042.545 ;
        RECT 210.045 3041.915 210.215 3042.085 ;
        RECT 210.045 3041.455 210.215 3041.625 ;
        RECT 210.045 3040.995 210.215 3041.165 ;
        RECT 210.045 3040.535 210.215 3040.705 ;
        RECT 210.045 3040.075 210.215 3040.245 ;
        RECT 210.045 3039.615 210.215 3039.785 ;
        RECT 210.045 3039.155 210.215 3039.325 ;
        RECT 210.045 3037.775 210.215 3037.945 ;
        RECT 210.045 3037.315 210.215 3037.485 ;
        RECT 210.045 3036.855 210.215 3037.025 ;
        RECT 210.045 3036.395 210.215 3036.565 ;
        RECT 210.045 3035.935 210.215 3036.105 ;
        RECT 210.045 3035.475 210.215 3035.645 ;
        RECT 210.045 3035.015 210.215 3035.185 ;
        RECT 210.045 3034.555 210.215 3034.725 ;
        RECT 210.045 3034.095 210.215 3034.265 ;
        RECT 210.045 3033.635 210.215 3033.805 ;
        RECT 210.045 3033.175 210.215 3033.345 ;
        RECT 210.045 3031.795 210.215 3031.965 ;
        RECT 210.045 3031.335 210.215 3031.505 ;
        RECT 210.045 3030.875 210.215 3031.045 ;
        RECT 210.045 3030.415 210.215 3030.585 ;
        RECT 210.045 3029.955 210.215 3030.125 ;
        RECT 210.045 3029.495 210.215 3029.665 ;
        RECT 210.045 3029.035 210.215 3029.205 ;
        RECT 210.045 3028.575 210.215 3028.745 ;
        RECT 210.045 3028.115 210.215 3028.285 ;
        RECT 210.045 3027.655 210.215 3027.825 ;
        RECT 210.045 3027.195 210.215 3027.365 ;
        RECT 210.045 3025.815 210.215 3025.985 ;
        RECT 210.045 3025.355 210.215 3025.525 ;
        RECT 210.045 3024.895 210.215 3025.065 ;
        RECT 210.045 3024.435 210.215 3024.605 ;
        RECT 210.045 3023.975 210.215 3024.145 ;
        RECT 210.045 3023.515 210.215 3023.685 ;
        RECT 210.045 3023.055 210.215 3023.225 ;
        RECT 210.045 3022.595 210.215 3022.765 ;
        RECT 210.045 3022.135 210.215 3022.305 ;
        RECT 210.045 3021.675 210.215 3021.845 ;
        RECT 210.045 3021.215 210.215 3021.385 ;
        RECT 210.045 3019.835 210.215 3020.005 ;
        RECT 210.045 3019.375 210.215 3019.545 ;
        RECT 210.045 3018.915 210.215 3019.085 ;
        RECT 210.045 3018.455 210.215 3018.625 ;
        RECT 210.045 3017.995 210.215 3018.165 ;
        RECT 210.045 3017.535 210.215 3017.705 ;
        RECT 210.045 3017.075 210.215 3017.245 ;
        RECT 210.045 3016.615 210.215 3016.785 ;
        RECT 210.045 3016.155 210.215 3016.325 ;
        RECT 210.045 3015.695 210.215 3015.865 ;
        RECT 210.045 3015.235 210.215 3015.405 ;
        RECT 210.045 3013.855 210.215 3014.025 ;
        RECT 210.045 3013.395 210.215 3013.565 ;
        RECT 210.045 3012.935 210.215 3013.105 ;
        RECT 210.045 3012.475 210.215 3012.645 ;
        RECT 210.045 3012.015 210.215 3012.185 ;
        RECT 210.045 3011.555 210.215 3011.725 ;
        RECT 210.045 3011.095 210.215 3011.265 ;
        RECT 210.045 3010.635 210.215 3010.805 ;
        RECT 210.045 3010.175 210.215 3010.345 ;
        RECT 210.045 3009.715 210.215 3009.885 ;
        RECT 210.045 3009.255 210.215 3009.425 ;
        RECT 210.045 3007.875 210.215 3008.045 ;
        RECT 210.045 3007.415 210.215 3007.585 ;
        RECT 210.045 3006.955 210.215 3007.125 ;
        RECT 210.045 3006.495 210.215 3006.665 ;
        RECT 210.045 3006.035 210.215 3006.205 ;
        RECT 210.045 3005.575 210.215 3005.745 ;
        RECT 210.045 3005.115 210.215 3005.285 ;
        RECT 210.045 3004.655 210.215 3004.825 ;
        RECT 210.045 3004.195 210.215 3004.365 ;
        RECT 210.045 3003.735 210.215 3003.905 ;
        RECT 210.045 3003.275 210.215 3003.445 ;
        RECT 210.045 3001.895 210.215 3002.065 ;
        RECT 210.045 3001.435 210.215 3001.605 ;
        RECT 210.045 3000.975 210.215 3001.145 ;
        RECT 210.045 3000.515 210.215 3000.685 ;
        RECT 210.045 3000.055 210.215 3000.225 ;
        RECT 210.045 2999.595 210.215 2999.765 ;
        RECT 210.045 2999.135 210.215 2999.305 ;
        RECT 210.045 2998.675 210.215 2998.845 ;
        RECT 210.045 2998.215 210.215 2998.385 ;
        RECT 210.045 2997.755 210.215 2997.925 ;
        RECT 210.045 2997.295 210.215 2997.465 ;
        RECT 210.045 2995.915 210.215 2996.085 ;
        RECT 210.045 2995.455 210.215 2995.625 ;
        RECT 210.045 2994.995 210.215 2995.165 ;
        RECT 210.045 2994.535 210.215 2994.705 ;
        RECT 210.045 2994.075 210.215 2994.245 ;
        RECT 210.045 2993.615 210.215 2993.785 ;
        RECT 210.045 2993.155 210.215 2993.325 ;
        RECT 210.045 2992.695 210.215 2992.865 ;
        RECT 210.045 2992.235 210.215 2992.405 ;
        RECT 210.045 2991.775 210.215 2991.945 ;
        RECT 210.045 2991.315 210.215 2991.485 ;
        RECT 210.045 2989.935 210.215 2990.105 ;
        RECT 210.045 2989.475 210.215 2989.645 ;
        RECT 210.045 2989.015 210.215 2989.185 ;
        RECT 210.045 2988.555 210.215 2988.725 ;
        RECT 210.045 2988.095 210.215 2988.265 ;
        RECT 210.045 2987.635 210.215 2987.805 ;
        RECT 210.045 2987.175 210.215 2987.345 ;
        RECT 210.045 2986.715 210.215 2986.885 ;
        RECT 210.045 2986.255 210.215 2986.425 ;
        RECT 210.045 2985.795 210.215 2985.965 ;
        RECT 210.045 2985.335 210.215 2985.505 ;
      LAYER met1 ;
        RECT 204.450 2984.730 204.930 3050.970 ;
        RECT 209.890 2984.730 210.370 3050.970 ;
      LAYER via ;
        RECT 204.560 3017.070 204.860 3018.855 ;
        RECT 210.000 3017.070 210.300 3018.855 ;
      LAYER met2 ;
        RECT 204.500 3017.030 204.930 3018.895 ;
        RECT 209.940 3017.030 210.370 3018.895 ;
      LAYER via2 ;
        RECT 204.560 3017.070 204.860 3018.855 ;
        RECT 210.000 3017.070 210.300 3018.855 ;
      LAYER met3 ;
        RECT 200.115 3017.035 210.370 3018.885 ;
    END
    PORT
      LAYER li1 ;
        RECT 204.480 4456.885 204.650 4457.055 ;
        RECT 209.920 4456.885 210.090 4457.055 ;
      LAYER li1 ;
        RECT 209.920 4456.655 210.090 4456.740 ;
      LAYER li1 ;
        RECT 204.480 4456.425 204.650 4456.595 ;
        RECT 204.480 4455.965 204.650 4456.135 ;
        RECT 204.480 4455.505 204.650 4455.675 ;
        RECT 204.480 4455.045 204.650 4455.215 ;
        RECT 204.480 4454.585 204.650 4454.755 ;
        RECT 204.480 4454.125 204.650 4454.295 ;
        RECT 204.480 4453.665 204.650 4453.835 ;
        RECT 204.480 4453.205 204.650 4453.375 ;
      LAYER li1 ;
        RECT 209.485 4453.250 210.090 4456.655 ;
      LAYER li1 ;
        RECT 204.480 4452.745 204.650 4452.915 ;
      LAYER li1 ;
        RECT 208.235 4452.900 210.090 4453.250 ;
      LAYER li1 ;
        RECT 204.480 4452.285 204.650 4452.455 ;
        RECT 204.480 4451.825 204.650 4451.995 ;
        RECT 204.480 4451.365 204.650 4451.535 ;
      LAYER li1 ;
        RECT 209.485 4451.310 210.090 4452.900 ;
        RECT 209.920 4451.220 210.090 4451.310 ;
      LAYER li1 ;
        RECT 204.480 4450.905 204.650 4451.075 ;
        RECT 209.920 4450.905 210.090 4451.075 ;
      LAYER li1 ;
        RECT 209.920 4450.675 210.090 4450.760 ;
      LAYER li1 ;
        RECT 204.480 4450.445 204.650 4450.615 ;
        RECT 204.480 4449.985 204.650 4450.155 ;
        RECT 204.480 4449.525 204.650 4449.695 ;
        RECT 204.480 4449.065 204.650 4449.235 ;
        RECT 204.480 4448.605 204.650 4448.775 ;
        RECT 204.480 4448.145 204.650 4448.315 ;
        RECT 204.480 4447.685 204.650 4447.855 ;
        RECT 204.480 4447.225 204.650 4447.395 ;
      LAYER li1 ;
        RECT 209.485 4447.270 210.090 4450.675 ;
      LAYER li1 ;
        RECT 204.480 4446.765 204.650 4446.935 ;
      LAYER li1 ;
        RECT 208.235 4446.920 210.090 4447.270 ;
      LAYER li1 ;
        RECT 204.480 4446.305 204.650 4446.475 ;
        RECT 204.480 4445.845 204.650 4446.015 ;
        RECT 204.480 4445.385 204.650 4445.555 ;
      LAYER li1 ;
        RECT 209.485 4445.330 210.090 4446.920 ;
        RECT 209.920 4445.240 210.090 4445.330 ;
      LAYER li1 ;
        RECT 204.480 4444.925 204.650 4445.095 ;
        RECT 209.920 4444.925 210.090 4445.095 ;
      LAYER li1 ;
        RECT 209.920 4444.695 210.090 4444.780 ;
      LAYER li1 ;
        RECT 204.480 4444.465 204.650 4444.635 ;
        RECT 204.480 4444.005 204.650 4444.175 ;
        RECT 204.480 4443.545 204.650 4443.715 ;
        RECT 204.480 4443.085 204.650 4443.255 ;
        RECT 204.480 4442.625 204.650 4442.795 ;
        RECT 204.480 4442.165 204.650 4442.335 ;
        RECT 204.480 4441.705 204.650 4441.875 ;
        RECT 204.480 4441.245 204.650 4441.415 ;
      LAYER li1 ;
        RECT 209.485 4441.290 210.090 4444.695 ;
      LAYER li1 ;
        RECT 204.480 4440.785 204.650 4440.955 ;
      LAYER li1 ;
        RECT 208.235 4440.940 210.090 4441.290 ;
      LAYER li1 ;
        RECT 204.480 4440.325 204.650 4440.495 ;
        RECT 204.480 4439.865 204.650 4440.035 ;
        RECT 204.480 4439.405 204.650 4439.575 ;
      LAYER li1 ;
        RECT 209.485 4439.350 210.090 4440.940 ;
        RECT 209.920 4439.260 210.090 4439.350 ;
      LAYER li1 ;
        RECT 204.480 4438.945 204.650 4439.115 ;
        RECT 209.920 4438.945 210.090 4439.115 ;
      LAYER li1 ;
        RECT 209.920 4438.715 210.090 4438.800 ;
      LAYER li1 ;
        RECT 204.480 4438.485 204.650 4438.655 ;
        RECT 204.480 4438.025 204.650 4438.195 ;
        RECT 204.480 4437.565 204.650 4437.735 ;
        RECT 204.480 4437.105 204.650 4437.275 ;
        RECT 204.480 4436.645 204.650 4436.815 ;
        RECT 204.480 4436.185 204.650 4436.355 ;
        RECT 204.480 4435.725 204.650 4435.895 ;
        RECT 204.480 4435.265 204.650 4435.435 ;
      LAYER li1 ;
        RECT 209.485 4435.310 210.090 4438.715 ;
      LAYER li1 ;
        RECT 204.480 4434.805 204.650 4434.975 ;
      LAYER li1 ;
        RECT 208.235 4434.960 210.090 4435.310 ;
      LAYER li1 ;
        RECT 204.480 4434.345 204.650 4434.515 ;
        RECT 204.480 4433.885 204.650 4434.055 ;
        RECT 204.480 4433.425 204.650 4433.595 ;
      LAYER li1 ;
        RECT 209.485 4433.370 210.090 4434.960 ;
        RECT 209.920 4433.280 210.090 4433.370 ;
      LAYER li1 ;
        RECT 204.480 4432.965 204.650 4433.135 ;
        RECT 209.920 4432.965 210.090 4433.135 ;
      LAYER li1 ;
        RECT 209.920 4432.735 210.090 4432.820 ;
      LAYER li1 ;
        RECT 204.480 4432.505 204.650 4432.675 ;
        RECT 204.480 4432.045 204.650 4432.215 ;
        RECT 204.480 4431.585 204.650 4431.755 ;
        RECT 204.480 4431.125 204.650 4431.295 ;
        RECT 204.480 4430.665 204.650 4430.835 ;
        RECT 204.480 4430.205 204.650 4430.375 ;
        RECT 204.480 4429.745 204.650 4429.915 ;
        RECT 204.480 4429.285 204.650 4429.455 ;
      LAYER li1 ;
        RECT 209.485 4429.330 210.090 4432.735 ;
      LAYER li1 ;
        RECT 204.480 4428.825 204.650 4428.995 ;
      LAYER li1 ;
        RECT 208.235 4428.980 210.090 4429.330 ;
      LAYER li1 ;
        RECT 204.480 4428.365 204.650 4428.535 ;
        RECT 204.480 4427.905 204.650 4428.075 ;
        RECT 204.480 4427.445 204.650 4427.615 ;
      LAYER li1 ;
        RECT 209.485 4427.390 210.090 4428.980 ;
        RECT 209.920 4427.300 210.090 4427.390 ;
      LAYER li1 ;
        RECT 204.480 4426.985 204.650 4427.155 ;
        RECT 209.920 4426.985 210.090 4427.155 ;
      LAYER mcon ;
        RECT 209.920 4455.965 210.090 4456.135 ;
        RECT 209.920 4455.505 210.090 4455.675 ;
        RECT 209.920 4455.045 210.090 4455.215 ;
        RECT 209.920 4454.585 210.090 4454.755 ;
        RECT 209.920 4454.125 210.090 4454.295 ;
        RECT 209.920 4453.665 210.090 4453.835 ;
        RECT 209.920 4453.205 210.090 4453.375 ;
        RECT 209.920 4452.745 210.090 4452.915 ;
        RECT 209.920 4452.285 210.090 4452.455 ;
        RECT 209.920 4451.825 210.090 4451.995 ;
        RECT 209.920 4451.365 210.090 4451.535 ;
        RECT 209.920 4449.985 210.090 4450.155 ;
        RECT 209.920 4449.525 210.090 4449.695 ;
        RECT 209.920 4449.065 210.090 4449.235 ;
        RECT 209.920 4448.605 210.090 4448.775 ;
        RECT 209.920 4448.145 210.090 4448.315 ;
        RECT 209.920 4447.685 210.090 4447.855 ;
        RECT 209.920 4447.225 210.090 4447.395 ;
        RECT 209.920 4446.765 210.090 4446.935 ;
        RECT 209.920 4446.305 210.090 4446.475 ;
        RECT 209.920 4445.845 210.090 4446.015 ;
        RECT 209.920 4445.385 210.090 4445.555 ;
        RECT 209.920 4444.005 210.090 4444.175 ;
        RECT 209.920 4443.545 210.090 4443.715 ;
        RECT 209.920 4443.085 210.090 4443.255 ;
        RECT 209.920 4442.625 210.090 4442.795 ;
        RECT 209.920 4442.165 210.090 4442.335 ;
        RECT 209.920 4441.705 210.090 4441.875 ;
        RECT 209.920 4441.245 210.090 4441.415 ;
        RECT 209.920 4440.785 210.090 4440.955 ;
        RECT 209.920 4440.325 210.090 4440.495 ;
        RECT 209.920 4439.865 210.090 4440.035 ;
        RECT 209.920 4439.405 210.090 4439.575 ;
        RECT 209.920 4438.025 210.090 4438.195 ;
        RECT 209.920 4437.565 210.090 4437.735 ;
        RECT 209.920 4437.105 210.090 4437.275 ;
        RECT 209.920 4436.645 210.090 4436.815 ;
        RECT 209.920 4436.185 210.090 4436.355 ;
        RECT 209.920 4435.725 210.090 4435.895 ;
        RECT 209.920 4435.265 210.090 4435.435 ;
        RECT 209.920 4434.805 210.090 4434.975 ;
        RECT 209.920 4434.345 210.090 4434.515 ;
        RECT 209.920 4433.885 210.090 4434.055 ;
        RECT 209.920 4433.425 210.090 4433.595 ;
        RECT 209.920 4432.045 210.090 4432.215 ;
        RECT 209.920 4431.585 210.090 4431.755 ;
        RECT 209.920 4431.125 210.090 4431.295 ;
        RECT 209.920 4430.665 210.090 4430.835 ;
        RECT 209.920 4430.205 210.090 4430.375 ;
        RECT 209.920 4429.745 210.090 4429.915 ;
        RECT 209.920 4429.285 210.090 4429.455 ;
        RECT 209.920 4428.825 210.090 4428.995 ;
        RECT 209.920 4428.365 210.090 4428.535 ;
        RECT 209.920 4427.905 210.090 4428.075 ;
        RECT 209.920 4427.445 210.090 4427.615 ;
      LAYER met1 ;
        RECT 204.325 4426.840 204.805 4457.200 ;
        RECT 209.765 4426.840 210.245 4457.200 ;
      LAYER via ;
        RECT 204.405 4440.940 204.705 4442.725 ;
        RECT 209.845 4440.940 210.145 4442.725 ;
      LAYER met2 ;
        RECT 204.345 4440.900 204.775 4442.765 ;
        RECT 209.785 4440.900 210.215 4442.765 ;
      LAYER via2 ;
        RECT 204.405 4440.940 204.705 4442.725 ;
        RECT 209.845 4440.940 210.145 4442.725 ;
      LAYER met3 ;
        RECT 199.960 4440.905 210.215 4442.755 ;
    END
  END vccd
  OBS
      LAYER pwell ;
        RECT 2088.490 4987.595 2088.660 4987.785 ;
        RECT 2082.845 4986.725 2083.275 4987.510 ;
        RECT 2083.675 4986.685 2088.805 4987.595 ;
        RECT 2088.825 4986.725 2089.255 4987.510 ;
        RECT 3315.495 4987.185 3315.665 4987.375 ;
        RECT 3321.475 4987.185 3321.645 4987.375 ;
        RECT 3327.455 4987.185 3327.625 4987.375 ;
        RECT 3333.435 4987.185 3333.605 4987.375 ;
        RECT 835.260 4985.970 835.430 4986.160 ;
        RECT 841.240 4985.970 841.410 4986.160 ;
        RECT 847.220 4985.970 847.390 4986.160 ;
        RECT 834.665 4985.100 835.095 4985.885 ;
        RECT 835.115 4985.060 840.245 4985.970 ;
        RECT 840.645 4985.100 841.075 4985.885 ;
        RECT 841.095 4985.060 846.225 4985.970 ;
        RECT 846.625 4985.100 847.055 4985.885 ;
        RECT 847.075 4985.060 852.205 4985.970 ;
        RECT 852.605 4985.100 853.035 4985.885 ;
      LAYER nwell ;
        RECT 834.460 4981.940 853.240 4984.770 ;
        RECT 2082.640 4983.565 2089.460 4986.395 ;
      LAYER pwell ;
        RECT 3309.850 4986.315 3310.280 4987.100 ;
        RECT 3310.680 4986.275 3315.810 4987.185 ;
        RECT 3315.830 4986.315 3316.260 4987.100 ;
        RECT 3316.660 4986.275 3321.790 4987.185 ;
        RECT 3321.810 4986.315 3322.240 4987.100 ;
        RECT 3322.640 4986.275 3327.770 4987.185 ;
        RECT 3327.790 4986.315 3328.220 4987.100 ;
        RECT 3328.620 4986.275 3333.750 4987.185 ;
        RECT 3333.770 4986.315 3334.200 4987.100 ;
        RECT 2082.845 4982.450 2083.275 4983.235 ;
        RECT 2083.295 4982.365 2088.425 4983.275 ;
        RECT 2088.825 4982.450 2089.255 4983.235 ;
      LAYER nwell ;
        RECT 3309.645 4983.155 3334.405 4985.985 ;
      LAYER pwell ;
        RECT 2083.440 4982.175 2083.610 4982.365 ;
        RECT 2088.450 4982.110 2088.730 4982.390 ;
        RECT 834.665 4980.825 835.095 4981.610 ;
        RECT 835.495 4980.740 840.625 4981.650 ;
        RECT 840.645 4980.825 841.075 4981.610 ;
        RECT 841.475 4980.740 846.605 4981.650 ;
        RECT 846.625 4980.825 847.055 4981.610 ;
        RECT 847.455 4980.740 852.585 4981.650 ;
        RECT 852.605 4980.825 853.035 4981.610 ;
        RECT 2082.845 4981.285 2083.275 4982.070 ;
        RECT 2088.825 4981.285 2089.255 4982.070 ;
        RECT 3309.850 4982.040 3310.280 4982.825 ;
        RECT 3310.300 4981.955 3315.430 4982.865 ;
        RECT 3315.830 4982.040 3316.260 4982.825 ;
        RECT 3310.445 4981.765 3310.615 4981.955 ;
        RECT 3315.455 4981.700 3315.735 4981.980 ;
        RECT 3316.280 4981.955 3321.410 4982.865 ;
        RECT 3321.810 4982.040 3322.240 4982.825 ;
        RECT 3316.425 4981.765 3316.595 4981.955 ;
        RECT 3321.435 4981.700 3321.715 4981.980 ;
        RECT 3322.260 4981.955 3327.390 4982.865 ;
        RECT 3327.790 4982.040 3328.220 4982.825 ;
        RECT 3322.405 4981.765 3322.575 4981.955 ;
        RECT 3327.415 4981.700 3327.695 4981.980 ;
        RECT 3328.240 4981.955 3333.370 4982.865 ;
        RECT 3333.770 4982.040 3334.200 4982.825 ;
        RECT 3328.385 4981.765 3328.555 4981.955 ;
        RECT 3333.395 4981.700 3333.675 4981.980 ;
        RECT 840.270 4980.485 840.550 4980.740 ;
        RECT 846.250 4980.485 846.530 4980.740 ;
        RECT 852.230 4980.485 852.510 4980.740 ;
        RECT 834.665 4979.660 835.095 4980.445 ;
        RECT 840.645 4979.660 841.075 4980.445 ;
        RECT 846.625 4979.660 847.055 4980.445 ;
        RECT 852.605 4979.660 853.035 4980.445 ;
      LAYER nwell ;
        RECT 2082.640 4979.350 2089.460 4980.955 ;
      LAYER pwell ;
        RECT 3309.850 4980.875 3310.280 4981.660 ;
        RECT 3315.830 4980.875 3316.260 4981.660 ;
        RECT 3321.810 4980.875 3322.240 4981.660 ;
        RECT 3327.790 4980.875 3328.220 4981.660 ;
        RECT 3333.770 4980.875 3334.200 4981.660 ;
      LAYER nwell ;
        RECT 834.460 4977.725 853.240 4979.330 ;
        RECT 3309.645 4978.940 3334.405 4980.545 ;
      LAYER pwell ;
        RECT 202.035 4456.755 202.820 4457.185 ;
        RECT 201.950 4451.540 202.860 4456.355 ;
        RECT 201.760 4451.370 202.860 4451.540 ;
        RECT 201.950 4451.225 202.860 4451.370 ;
        RECT 202.035 4450.775 202.820 4451.205 ;
        RECT 201.950 4445.560 202.860 4450.375 ;
        RECT 201.760 4445.390 202.860 4445.560 ;
        RECT 201.950 4445.245 202.860 4445.390 ;
        RECT 202.035 4444.795 202.820 4445.225 ;
        RECT 201.950 4439.580 202.860 4444.395 ;
        RECT 201.760 4439.410 202.860 4439.580 ;
        RECT 201.950 4439.265 202.860 4439.410 ;
        RECT 202.035 4438.815 202.820 4439.245 ;
        RECT 201.950 4433.600 202.860 4438.415 ;
        RECT 201.760 4433.430 202.860 4433.600 ;
        RECT 201.950 4433.285 202.860 4433.430 ;
        RECT 202.035 4432.835 202.820 4433.265 ;
        RECT 201.950 4427.620 202.860 4432.435 ;
        RECT 201.760 4427.450 202.860 4427.620 ;
        RECT 201.950 4427.305 202.860 4427.450 ;
        RECT 202.035 4426.855 202.820 4427.285 ;
      LAYER nwell ;
        RECT 203.150 4426.650 205.980 4457.390 ;
      LAYER pwell ;
        RECT 206.310 4456.755 207.095 4457.185 ;
        RECT 207.475 4456.755 208.260 4457.185 ;
        RECT 206.270 4456.660 207.180 4456.735 ;
        RECT 206.270 4456.380 207.435 4456.660 ;
        RECT 206.270 4451.605 207.180 4456.380 ;
        RECT 206.310 4450.775 207.095 4451.205 ;
        RECT 207.475 4450.775 208.260 4451.205 ;
        RECT 206.270 4450.680 207.180 4450.755 ;
        RECT 206.270 4450.400 207.435 4450.680 ;
        RECT 206.270 4445.625 207.180 4450.400 ;
        RECT 206.310 4444.795 207.095 4445.225 ;
        RECT 207.475 4444.795 208.260 4445.225 ;
        RECT 206.270 4444.700 207.180 4444.775 ;
        RECT 206.270 4444.420 207.435 4444.700 ;
        RECT 206.270 4439.645 207.180 4444.420 ;
        RECT 206.310 4438.815 207.095 4439.245 ;
        RECT 207.475 4438.815 208.260 4439.245 ;
        RECT 206.270 4438.720 207.180 4438.795 ;
        RECT 206.270 4438.440 207.435 4438.720 ;
        RECT 206.270 4433.665 207.180 4438.440 ;
        RECT 206.310 4432.835 207.095 4433.265 ;
        RECT 207.475 4432.835 208.260 4433.265 ;
        RECT 206.270 4432.740 207.180 4432.815 ;
        RECT 206.270 4432.460 207.435 4432.740 ;
        RECT 206.270 4427.685 207.180 4432.460 ;
        RECT 206.310 4426.855 207.095 4427.285 ;
        RECT 207.475 4426.855 208.260 4427.285 ;
      LAYER nwell ;
        RECT 208.590 4426.650 210.195 4457.390 ;
        RECT 3377.675 3601.870 3379.280 3638.590 ;
      LAYER pwell ;
        RECT 3379.610 3637.955 3380.395 3638.385 ;
        RECT 3380.775 3637.955 3381.560 3638.385 ;
        RECT 3380.690 3637.860 3381.600 3637.935 ;
        RECT 3380.435 3637.580 3381.600 3637.860 ;
        RECT 3380.690 3632.805 3381.600 3637.580 ;
        RECT 3379.610 3631.975 3380.395 3632.405 ;
        RECT 3380.775 3631.975 3381.560 3632.405 ;
        RECT 3380.690 3631.880 3381.600 3631.955 ;
        RECT 3380.435 3631.600 3381.600 3631.880 ;
        RECT 3380.690 3626.825 3381.600 3631.600 ;
        RECT 3379.610 3625.995 3380.395 3626.425 ;
        RECT 3380.775 3625.995 3381.560 3626.425 ;
        RECT 3380.690 3625.900 3381.600 3625.975 ;
        RECT 3380.435 3625.620 3381.600 3625.900 ;
        RECT 3380.690 3620.845 3381.600 3625.620 ;
        RECT 3379.610 3620.015 3380.395 3620.445 ;
        RECT 3380.775 3620.015 3381.560 3620.445 ;
        RECT 3380.690 3619.920 3381.600 3619.995 ;
        RECT 3380.435 3619.640 3381.600 3619.920 ;
        RECT 3380.690 3614.865 3381.600 3619.640 ;
        RECT 3379.610 3614.035 3380.395 3614.465 ;
        RECT 3380.775 3614.035 3381.560 3614.465 ;
        RECT 3380.690 3613.940 3381.600 3614.015 ;
        RECT 3380.435 3613.660 3381.600 3613.940 ;
        RECT 3380.690 3608.885 3381.600 3613.660 ;
        RECT 3379.610 3608.055 3380.395 3608.485 ;
        RECT 3380.775 3608.055 3381.560 3608.485 ;
        RECT 3380.690 3607.960 3381.600 3608.035 ;
        RECT 3380.435 3607.680 3381.600 3607.960 ;
        RECT 3380.690 3602.905 3381.600 3607.680 ;
        RECT 3379.610 3602.075 3380.395 3602.505 ;
        RECT 3380.775 3602.075 3381.560 3602.505 ;
      LAYER nwell ;
        RECT 3381.890 3601.870 3384.720 3638.590 ;
      LAYER pwell ;
        RECT 3385.050 3637.955 3385.835 3638.385 ;
        RECT 3385.010 3632.740 3385.920 3637.555 ;
        RECT 3385.010 3632.570 3386.110 3632.740 ;
        RECT 3385.010 3632.425 3385.920 3632.570 ;
        RECT 3385.050 3631.975 3385.835 3632.405 ;
        RECT 3385.010 3626.760 3385.920 3631.575 ;
        RECT 3385.010 3626.590 3386.110 3626.760 ;
        RECT 3385.010 3626.445 3385.920 3626.590 ;
        RECT 3385.050 3625.995 3385.835 3626.425 ;
        RECT 3385.010 3620.780 3385.920 3625.595 ;
        RECT 3385.010 3620.610 3386.110 3620.780 ;
        RECT 3385.010 3620.465 3385.920 3620.610 ;
        RECT 3385.050 3620.015 3385.835 3620.445 ;
        RECT 3385.010 3614.800 3385.920 3619.615 ;
        RECT 3385.010 3614.630 3386.110 3614.800 ;
        RECT 3385.010 3614.485 3385.920 3614.630 ;
        RECT 3385.050 3614.035 3385.835 3614.465 ;
        RECT 3385.010 3608.820 3385.920 3613.635 ;
        RECT 3385.010 3608.650 3386.110 3608.820 ;
        RECT 3385.010 3608.505 3385.920 3608.650 ;
        RECT 3385.050 3608.055 3385.835 3608.485 ;
        RECT 3385.010 3602.840 3385.920 3607.655 ;
        RECT 3385.010 3602.670 3386.110 3602.840 ;
        RECT 3385.010 3602.525 3385.920 3602.670 ;
        RECT 3385.050 3602.075 3385.835 3602.505 ;
        RECT 202.160 3050.525 202.945 3050.955 ;
        RECT 202.075 3045.310 202.985 3050.125 ;
        RECT 201.885 3045.140 202.985 3045.310 ;
        RECT 202.075 3044.995 202.985 3045.140 ;
        RECT 202.160 3044.545 202.945 3044.975 ;
        RECT 202.075 3039.330 202.985 3044.145 ;
        RECT 201.885 3039.160 202.985 3039.330 ;
        RECT 202.075 3039.015 202.985 3039.160 ;
        RECT 202.160 3038.565 202.945 3038.995 ;
        RECT 202.075 3033.350 202.985 3038.165 ;
        RECT 201.885 3033.180 202.985 3033.350 ;
        RECT 202.075 3033.035 202.985 3033.180 ;
        RECT 202.160 3032.585 202.945 3033.015 ;
        RECT 202.075 3027.370 202.985 3032.185 ;
        RECT 201.885 3027.200 202.985 3027.370 ;
        RECT 202.075 3027.055 202.985 3027.200 ;
        RECT 202.160 3026.605 202.945 3027.035 ;
        RECT 202.075 3021.390 202.985 3026.205 ;
        RECT 201.885 3021.220 202.985 3021.390 ;
        RECT 202.075 3021.075 202.985 3021.220 ;
        RECT 202.160 3020.625 202.945 3021.055 ;
        RECT 202.075 3015.410 202.985 3020.225 ;
        RECT 201.885 3015.240 202.985 3015.410 ;
        RECT 202.075 3015.095 202.985 3015.240 ;
        RECT 202.160 3014.645 202.945 3015.075 ;
        RECT 202.075 3009.430 202.985 3014.245 ;
        RECT 201.885 3009.260 202.985 3009.430 ;
        RECT 202.075 3009.115 202.985 3009.260 ;
        RECT 202.160 3008.665 202.945 3009.095 ;
        RECT 202.075 3003.450 202.985 3008.265 ;
        RECT 201.885 3003.280 202.985 3003.450 ;
        RECT 202.075 3003.135 202.985 3003.280 ;
        RECT 202.160 3002.685 202.945 3003.115 ;
        RECT 202.075 2997.470 202.985 3002.285 ;
        RECT 201.885 2997.300 202.985 2997.470 ;
        RECT 202.075 2997.155 202.985 2997.300 ;
        RECT 202.160 2996.705 202.945 2997.135 ;
        RECT 202.075 2991.490 202.985 2996.305 ;
        RECT 201.885 2991.320 202.985 2991.490 ;
        RECT 202.075 2991.175 202.985 2991.320 ;
        RECT 202.160 2990.725 202.945 2991.155 ;
        RECT 202.075 2985.510 202.985 2990.325 ;
        RECT 201.885 2985.340 202.985 2985.510 ;
        RECT 202.075 2985.195 202.985 2985.340 ;
        RECT 202.160 2984.745 202.945 2985.175 ;
      LAYER nwell ;
        RECT 203.275 2984.540 206.105 3051.160 ;
      LAYER pwell ;
        RECT 206.435 3050.525 207.220 3050.955 ;
        RECT 207.600 3050.525 208.385 3050.955 ;
        RECT 206.395 3050.430 207.305 3050.505 ;
        RECT 206.395 3050.150 207.560 3050.430 ;
        RECT 206.395 3045.375 207.305 3050.150 ;
        RECT 206.435 3044.545 207.220 3044.975 ;
        RECT 207.600 3044.545 208.385 3044.975 ;
        RECT 206.395 3044.450 207.305 3044.525 ;
        RECT 206.395 3044.170 207.560 3044.450 ;
        RECT 206.395 3039.395 207.305 3044.170 ;
        RECT 206.435 3038.565 207.220 3038.995 ;
        RECT 207.600 3038.565 208.385 3038.995 ;
        RECT 206.395 3038.470 207.305 3038.545 ;
        RECT 206.395 3038.190 207.560 3038.470 ;
        RECT 206.395 3033.415 207.305 3038.190 ;
        RECT 206.435 3032.585 207.220 3033.015 ;
        RECT 207.600 3032.585 208.385 3033.015 ;
        RECT 206.395 3032.490 207.305 3032.565 ;
        RECT 206.395 3032.210 207.560 3032.490 ;
        RECT 206.395 3027.435 207.305 3032.210 ;
        RECT 206.435 3026.605 207.220 3027.035 ;
        RECT 207.600 3026.605 208.385 3027.035 ;
        RECT 206.395 3026.510 207.305 3026.585 ;
        RECT 206.395 3026.230 207.560 3026.510 ;
        RECT 206.395 3021.455 207.305 3026.230 ;
        RECT 206.435 3020.625 207.220 3021.055 ;
        RECT 207.600 3020.625 208.385 3021.055 ;
        RECT 206.395 3020.530 207.305 3020.605 ;
        RECT 206.395 3020.250 207.560 3020.530 ;
        RECT 206.395 3015.475 207.305 3020.250 ;
        RECT 206.435 3014.645 207.220 3015.075 ;
        RECT 207.600 3014.645 208.385 3015.075 ;
        RECT 206.395 3014.550 207.305 3014.625 ;
        RECT 206.395 3014.270 207.560 3014.550 ;
        RECT 206.395 3009.495 207.305 3014.270 ;
        RECT 206.435 3008.665 207.220 3009.095 ;
        RECT 207.600 3008.665 208.385 3009.095 ;
        RECT 206.395 3008.570 207.305 3008.645 ;
        RECT 206.395 3008.290 207.560 3008.570 ;
        RECT 206.395 3003.515 207.305 3008.290 ;
        RECT 206.435 3002.685 207.220 3003.115 ;
        RECT 207.600 3002.685 208.385 3003.115 ;
        RECT 206.395 3002.590 207.305 3002.665 ;
        RECT 206.395 3002.310 207.560 3002.590 ;
        RECT 206.395 2997.535 207.305 3002.310 ;
        RECT 206.435 2996.705 207.220 2997.135 ;
        RECT 207.600 2996.705 208.385 2997.135 ;
        RECT 206.395 2996.610 207.305 2996.685 ;
        RECT 206.395 2996.330 207.560 2996.610 ;
        RECT 206.395 2991.555 207.305 2996.330 ;
        RECT 206.435 2990.725 207.220 2991.155 ;
        RECT 207.600 2990.725 208.385 2991.155 ;
        RECT 206.395 2990.630 207.305 2990.705 ;
        RECT 206.395 2990.350 207.560 2990.630 ;
        RECT 206.395 2985.575 207.305 2990.350 ;
        RECT 206.435 2984.745 207.220 2985.175 ;
        RECT 207.600 2984.745 208.385 2985.175 ;
      LAYER nwell ;
        RECT 208.715 2984.540 210.320 3051.160 ;
        RECT 3377.675 2195.870 3379.280 2268.470 ;
      LAYER pwell ;
        RECT 3379.610 2267.835 3380.395 2268.265 ;
        RECT 3380.775 2267.835 3381.560 2268.265 ;
        RECT 3380.690 2267.740 3381.600 2267.815 ;
        RECT 3380.435 2267.460 3381.600 2267.740 ;
        RECT 3380.690 2262.685 3381.600 2267.460 ;
        RECT 3379.610 2261.855 3380.395 2262.285 ;
        RECT 3380.775 2261.855 3381.560 2262.285 ;
        RECT 3380.690 2261.760 3381.600 2261.835 ;
        RECT 3380.435 2261.480 3381.600 2261.760 ;
        RECT 3380.690 2256.705 3381.600 2261.480 ;
        RECT 3379.610 2255.875 3380.395 2256.305 ;
        RECT 3380.775 2255.875 3381.560 2256.305 ;
        RECT 3380.690 2255.780 3381.600 2255.855 ;
        RECT 3380.435 2255.500 3381.600 2255.780 ;
        RECT 3380.690 2250.725 3381.600 2255.500 ;
        RECT 3379.610 2249.895 3380.395 2250.325 ;
        RECT 3380.775 2249.895 3381.560 2250.325 ;
        RECT 3380.690 2249.800 3381.600 2249.875 ;
        RECT 3380.435 2249.520 3381.600 2249.800 ;
        RECT 3380.690 2244.745 3381.600 2249.520 ;
        RECT 3379.610 2243.915 3380.395 2244.345 ;
        RECT 3380.775 2243.915 3381.560 2244.345 ;
        RECT 3380.690 2243.820 3381.600 2243.895 ;
        RECT 3380.435 2243.540 3381.600 2243.820 ;
        RECT 3380.690 2238.765 3381.600 2243.540 ;
        RECT 3379.610 2237.935 3380.395 2238.365 ;
        RECT 3380.775 2237.935 3381.560 2238.365 ;
        RECT 3380.690 2237.840 3381.600 2237.915 ;
        RECT 3380.435 2237.560 3381.600 2237.840 ;
        RECT 3380.690 2232.785 3381.600 2237.560 ;
        RECT 3379.610 2231.955 3380.395 2232.385 ;
        RECT 3380.775 2231.955 3381.560 2232.385 ;
        RECT 3380.690 2231.860 3381.600 2231.935 ;
        RECT 3380.435 2231.580 3381.600 2231.860 ;
        RECT 3380.690 2226.805 3381.600 2231.580 ;
        RECT 3379.610 2225.975 3380.395 2226.405 ;
        RECT 3380.775 2225.975 3381.560 2226.405 ;
        RECT 3380.690 2225.880 3381.600 2225.955 ;
        RECT 3380.435 2225.600 3381.600 2225.880 ;
        RECT 3380.690 2220.825 3381.600 2225.600 ;
        RECT 3379.610 2219.995 3380.395 2220.425 ;
        RECT 3380.775 2219.995 3381.560 2220.425 ;
        RECT 3380.690 2219.900 3381.600 2219.975 ;
        RECT 3380.435 2219.620 3381.600 2219.900 ;
        RECT 3380.690 2214.845 3381.600 2219.620 ;
        RECT 3379.610 2214.015 3380.395 2214.445 ;
        RECT 3380.775 2214.015 3381.560 2214.445 ;
        RECT 3380.690 2213.920 3381.600 2213.995 ;
        RECT 3380.435 2213.640 3381.600 2213.920 ;
        RECT 3380.690 2208.865 3381.600 2213.640 ;
        RECT 3379.610 2208.035 3380.395 2208.465 ;
        RECT 3380.775 2208.035 3381.560 2208.465 ;
        RECT 3380.690 2207.940 3381.600 2208.015 ;
        RECT 3380.435 2207.660 3381.600 2207.940 ;
        RECT 3380.690 2202.885 3381.600 2207.660 ;
        RECT 3379.610 2202.055 3380.395 2202.485 ;
        RECT 3380.775 2202.055 3381.560 2202.485 ;
        RECT 3380.690 2201.960 3381.600 2202.035 ;
        RECT 3380.435 2201.680 3381.600 2201.960 ;
        RECT 3380.690 2196.905 3381.600 2201.680 ;
        RECT 3379.610 2196.075 3380.395 2196.505 ;
        RECT 3380.775 2196.075 3381.560 2196.505 ;
      LAYER nwell ;
        RECT 3381.890 2195.870 3384.720 2268.470 ;
      LAYER pwell ;
        RECT 3385.050 2267.835 3385.835 2268.265 ;
        RECT 3385.010 2262.620 3385.920 2267.435 ;
        RECT 3385.010 2262.450 3386.110 2262.620 ;
        RECT 3385.010 2262.305 3385.920 2262.450 ;
        RECT 3385.050 2261.855 3385.835 2262.285 ;
        RECT 3385.010 2256.640 3385.920 2261.455 ;
        RECT 3385.010 2256.470 3386.110 2256.640 ;
        RECT 3385.010 2256.325 3385.920 2256.470 ;
        RECT 3385.050 2255.875 3385.835 2256.305 ;
        RECT 3385.010 2250.660 3385.920 2255.475 ;
        RECT 3385.010 2250.490 3386.110 2250.660 ;
        RECT 3385.010 2250.345 3385.920 2250.490 ;
        RECT 3385.050 2249.895 3385.835 2250.325 ;
        RECT 3385.010 2244.680 3385.920 2249.495 ;
        RECT 3385.010 2244.510 3386.110 2244.680 ;
        RECT 3385.010 2244.365 3385.920 2244.510 ;
        RECT 3385.050 2243.915 3385.835 2244.345 ;
        RECT 3385.010 2238.700 3385.920 2243.515 ;
        RECT 3385.010 2238.530 3386.110 2238.700 ;
        RECT 3385.010 2238.385 3385.920 2238.530 ;
        RECT 3385.050 2237.935 3385.835 2238.365 ;
        RECT 3385.010 2232.720 3385.920 2237.535 ;
        RECT 3385.010 2232.550 3386.110 2232.720 ;
        RECT 3385.010 2232.405 3385.920 2232.550 ;
        RECT 3385.050 2231.955 3385.835 2232.385 ;
        RECT 3385.010 2226.740 3385.920 2231.555 ;
        RECT 3385.010 2226.570 3386.110 2226.740 ;
        RECT 3385.010 2226.425 3385.920 2226.570 ;
        RECT 3385.050 2225.975 3385.835 2226.405 ;
        RECT 3385.010 2220.760 3385.920 2225.575 ;
        RECT 3385.010 2220.590 3386.110 2220.760 ;
        RECT 3385.010 2220.445 3385.920 2220.590 ;
        RECT 3385.050 2219.995 3385.835 2220.425 ;
        RECT 3385.010 2214.780 3385.920 2219.595 ;
        RECT 3385.010 2214.610 3386.110 2214.780 ;
        RECT 3385.010 2214.465 3385.920 2214.610 ;
        RECT 3385.050 2214.015 3385.835 2214.445 ;
        RECT 3385.010 2208.800 3385.920 2213.615 ;
        RECT 3385.010 2208.630 3386.110 2208.800 ;
        RECT 3385.010 2208.485 3385.920 2208.630 ;
        RECT 3385.050 2208.035 3385.835 2208.465 ;
        RECT 3385.010 2202.820 3385.920 2207.635 ;
        RECT 3385.010 2202.650 3386.110 2202.820 ;
        RECT 3385.010 2202.505 3385.920 2202.650 ;
        RECT 3385.050 2202.055 3385.835 2202.485 ;
        RECT 3385.010 2196.840 3385.920 2201.655 ;
        RECT 3385.010 2196.670 3386.110 2196.840 ;
        RECT 3385.010 2196.525 3385.920 2196.670 ;
        RECT 3385.050 2196.075 3385.835 2196.505 ;
        RECT 202.270 1762.620 203.055 1763.050 ;
        RECT 202.185 1757.405 203.095 1762.220 ;
        RECT 201.995 1757.235 203.095 1757.405 ;
        RECT 202.185 1757.090 203.095 1757.235 ;
        RECT 202.270 1756.640 203.055 1757.070 ;
        RECT 202.185 1751.425 203.095 1756.240 ;
        RECT 201.995 1751.255 203.095 1751.425 ;
        RECT 202.185 1751.110 203.095 1751.255 ;
        RECT 202.270 1750.660 203.055 1751.090 ;
        RECT 202.185 1745.445 203.095 1750.260 ;
        RECT 201.995 1745.275 203.095 1745.445 ;
        RECT 202.185 1745.130 203.095 1745.275 ;
        RECT 202.270 1744.680 203.055 1745.110 ;
        RECT 202.185 1739.465 203.095 1744.280 ;
        RECT 201.995 1739.295 203.095 1739.465 ;
        RECT 202.185 1739.150 203.095 1739.295 ;
        RECT 202.270 1738.700 203.055 1739.130 ;
        RECT 202.185 1733.485 203.095 1738.300 ;
        RECT 201.995 1733.315 203.095 1733.485 ;
        RECT 202.185 1733.170 203.095 1733.315 ;
        RECT 202.270 1732.720 203.055 1733.150 ;
        RECT 202.185 1727.505 203.095 1732.320 ;
        RECT 201.995 1727.335 203.095 1727.505 ;
        RECT 202.185 1727.190 203.095 1727.335 ;
        RECT 202.270 1726.740 203.055 1727.170 ;
        RECT 202.185 1721.525 203.095 1726.340 ;
        RECT 201.995 1721.355 203.095 1721.525 ;
        RECT 202.185 1721.210 203.095 1721.355 ;
        RECT 202.270 1720.760 203.055 1721.190 ;
        RECT 202.185 1715.545 203.095 1720.360 ;
        RECT 201.995 1715.375 203.095 1715.545 ;
        RECT 202.185 1715.230 203.095 1715.375 ;
        RECT 202.270 1714.780 203.055 1715.210 ;
        RECT 202.185 1709.565 203.095 1714.380 ;
        RECT 201.995 1709.395 203.095 1709.565 ;
        RECT 202.185 1709.250 203.095 1709.395 ;
        RECT 202.270 1708.800 203.055 1709.230 ;
        RECT 202.185 1703.585 203.095 1708.400 ;
        RECT 201.995 1703.415 203.095 1703.585 ;
        RECT 202.185 1703.270 203.095 1703.415 ;
        RECT 202.270 1702.820 203.055 1703.250 ;
        RECT 202.185 1697.605 203.095 1702.420 ;
        RECT 201.995 1697.435 203.095 1697.605 ;
        RECT 202.185 1697.290 203.095 1697.435 ;
        RECT 202.270 1696.840 203.055 1697.270 ;
        RECT 202.185 1691.625 203.095 1696.440 ;
        RECT 201.995 1691.455 203.095 1691.625 ;
        RECT 202.185 1691.310 203.095 1691.455 ;
        RECT 202.270 1690.860 203.055 1691.290 ;
        RECT 202.185 1685.645 203.095 1690.460 ;
        RECT 201.995 1685.475 203.095 1685.645 ;
        RECT 202.185 1685.330 203.095 1685.475 ;
        RECT 202.270 1684.880 203.055 1685.310 ;
        RECT 202.185 1679.665 203.095 1684.480 ;
        RECT 201.995 1679.495 203.095 1679.665 ;
        RECT 202.185 1679.350 203.095 1679.495 ;
        RECT 202.270 1678.900 203.055 1679.330 ;
        RECT 202.185 1673.685 203.095 1678.500 ;
        RECT 201.995 1673.515 203.095 1673.685 ;
        RECT 202.185 1673.370 203.095 1673.515 ;
        RECT 202.270 1672.920 203.055 1673.350 ;
      LAYER nwell ;
        RECT 203.385 1672.715 206.215 1763.255 ;
      LAYER pwell ;
        RECT 206.545 1762.620 207.330 1763.050 ;
        RECT 207.710 1762.620 208.495 1763.050 ;
        RECT 206.505 1762.525 207.415 1762.600 ;
        RECT 206.505 1762.245 207.670 1762.525 ;
        RECT 206.505 1757.470 207.415 1762.245 ;
        RECT 206.545 1756.640 207.330 1757.070 ;
        RECT 207.710 1756.640 208.495 1757.070 ;
        RECT 206.505 1756.545 207.415 1756.620 ;
        RECT 206.505 1756.265 207.670 1756.545 ;
        RECT 206.505 1751.490 207.415 1756.265 ;
        RECT 206.545 1750.660 207.330 1751.090 ;
        RECT 207.710 1750.660 208.495 1751.090 ;
        RECT 206.505 1750.495 207.415 1750.640 ;
        RECT 207.625 1750.495 208.535 1750.640 ;
        RECT 206.505 1750.325 208.535 1750.495 ;
        RECT 206.505 1745.510 207.415 1750.325 ;
        RECT 207.625 1745.510 208.535 1750.325 ;
        RECT 206.545 1744.680 207.330 1745.110 ;
        RECT 207.710 1744.680 208.495 1745.110 ;
        RECT 206.505 1744.585 207.415 1744.660 ;
        RECT 206.505 1744.305 207.670 1744.585 ;
        RECT 206.505 1739.530 207.415 1744.305 ;
        RECT 206.545 1738.700 207.330 1739.130 ;
        RECT 207.710 1738.700 208.495 1739.130 ;
        RECT 206.505 1738.605 207.415 1738.680 ;
        RECT 206.505 1738.325 207.670 1738.605 ;
        RECT 206.505 1733.550 207.415 1738.325 ;
        RECT 206.545 1732.720 207.330 1733.150 ;
        RECT 207.710 1732.720 208.495 1733.150 ;
        RECT 206.505 1732.625 207.415 1732.700 ;
        RECT 206.505 1732.345 207.670 1732.625 ;
        RECT 206.505 1727.570 207.415 1732.345 ;
        RECT 206.545 1726.740 207.330 1727.170 ;
        RECT 207.710 1726.740 208.495 1727.170 ;
        RECT 206.505 1726.645 207.415 1726.720 ;
        RECT 206.505 1726.365 207.670 1726.645 ;
        RECT 206.505 1721.590 207.415 1726.365 ;
        RECT 206.545 1720.760 207.330 1721.190 ;
        RECT 207.710 1720.760 208.495 1721.190 ;
        RECT 206.505 1720.665 207.415 1720.740 ;
        RECT 206.505 1720.385 207.670 1720.665 ;
        RECT 206.505 1715.610 207.415 1720.385 ;
        RECT 206.545 1714.780 207.330 1715.210 ;
        RECT 207.710 1714.780 208.495 1715.210 ;
        RECT 206.505 1714.685 207.415 1714.760 ;
        RECT 206.505 1714.405 207.670 1714.685 ;
        RECT 206.505 1709.630 207.415 1714.405 ;
        RECT 206.545 1708.800 207.330 1709.230 ;
        RECT 207.710 1708.800 208.495 1709.230 ;
        RECT 206.505 1708.705 207.415 1708.780 ;
        RECT 206.505 1708.425 207.670 1708.705 ;
        RECT 206.505 1703.650 207.415 1708.425 ;
        RECT 206.545 1702.820 207.330 1703.250 ;
        RECT 207.710 1702.820 208.495 1703.250 ;
        RECT 206.505 1702.725 207.415 1702.800 ;
        RECT 206.505 1702.445 207.670 1702.725 ;
        RECT 206.505 1697.670 207.415 1702.445 ;
        RECT 206.545 1696.840 207.330 1697.270 ;
        RECT 207.710 1696.840 208.495 1697.270 ;
        RECT 206.505 1696.745 207.415 1696.820 ;
        RECT 206.505 1696.465 207.670 1696.745 ;
        RECT 206.505 1691.690 207.415 1696.465 ;
        RECT 206.545 1690.860 207.330 1691.290 ;
        RECT 207.710 1690.860 208.495 1691.290 ;
        RECT 206.505 1690.765 207.415 1690.840 ;
        RECT 206.505 1690.485 207.670 1690.765 ;
        RECT 206.505 1685.710 207.415 1690.485 ;
        RECT 206.545 1684.880 207.330 1685.310 ;
        RECT 207.710 1684.880 208.495 1685.310 ;
        RECT 206.505 1684.785 207.415 1684.860 ;
        RECT 206.505 1684.505 207.670 1684.785 ;
        RECT 206.505 1679.730 207.415 1684.505 ;
        RECT 206.545 1678.900 207.330 1679.330 ;
        RECT 207.710 1678.900 208.495 1679.330 ;
        RECT 206.505 1678.805 207.415 1678.880 ;
        RECT 206.505 1678.525 207.670 1678.805 ;
        RECT 206.505 1673.750 207.415 1678.525 ;
        RECT 206.545 1672.920 207.330 1673.350 ;
        RECT 207.710 1672.920 208.495 1673.350 ;
      LAYER nwell ;
        RECT 208.825 1672.715 210.430 1763.255 ;
        RECT 668.810 218.430 795.230 220.035 ;
        RECT 2145.810 218.430 2272.230 220.035 ;
      LAYER pwell ;
        RECT 669.015 217.315 669.445 218.100 ;
        RECT 674.995 217.315 675.425 218.100 ;
        RECT 680.975 217.315 681.405 218.100 ;
        RECT 686.955 217.315 687.385 218.100 ;
        RECT 692.935 217.315 693.365 218.100 ;
        RECT 698.915 217.315 699.345 218.100 ;
        RECT 704.895 217.315 705.325 218.100 ;
        RECT 710.875 217.315 711.305 218.100 ;
        RECT 716.855 217.315 717.285 218.100 ;
        RECT 722.835 217.315 723.265 218.100 ;
        RECT 728.815 217.315 729.245 218.100 ;
        RECT 734.795 217.315 735.225 218.100 ;
        RECT 740.775 217.315 741.205 218.100 ;
        RECT 746.755 217.315 747.185 218.100 ;
        RECT 752.735 217.315 753.165 218.100 ;
        RECT 758.715 217.315 759.145 218.100 ;
        RECT 764.695 217.315 765.125 218.100 ;
        RECT 770.675 217.315 771.105 218.100 ;
        RECT 776.655 217.315 777.085 218.100 ;
        RECT 782.635 217.315 783.065 218.100 ;
        RECT 788.615 217.315 789.045 218.100 ;
        RECT 794.595 217.315 795.025 218.100 ;
        RECT 2146.015 217.315 2146.445 218.100 ;
        RECT 2151.995 217.315 2152.425 218.100 ;
        RECT 2157.975 217.315 2158.405 218.100 ;
        RECT 2163.955 217.315 2164.385 218.100 ;
        RECT 2169.935 217.315 2170.365 218.100 ;
        RECT 2175.915 217.315 2176.345 218.100 ;
        RECT 2181.895 217.315 2182.325 218.100 ;
        RECT 2187.875 217.315 2188.305 218.100 ;
        RECT 2193.855 217.315 2194.285 218.100 ;
        RECT 2199.835 217.315 2200.265 218.100 ;
        RECT 2205.815 217.315 2206.245 218.100 ;
        RECT 2211.795 217.315 2212.225 218.100 ;
        RECT 2217.775 217.315 2218.205 218.100 ;
        RECT 2223.755 217.315 2224.185 218.100 ;
        RECT 2229.735 217.315 2230.165 218.100 ;
        RECT 2235.715 217.315 2236.145 218.100 ;
        RECT 2241.695 217.315 2242.125 218.100 ;
        RECT 2247.675 217.315 2248.105 218.100 ;
        RECT 2253.655 217.315 2254.085 218.100 ;
        RECT 2259.635 217.315 2260.065 218.100 ;
        RECT 2265.615 217.315 2266.045 218.100 ;
        RECT 2271.595 217.315 2272.025 218.100 ;
        RECT 669.540 216.995 669.820 217.275 ;
        RECT 674.660 217.020 674.830 217.210 ;
        RECT 669.015 216.150 669.445 216.935 ;
        RECT 669.845 216.110 674.975 217.020 ;
        RECT 675.520 216.995 675.800 217.275 ;
        RECT 680.640 217.020 680.810 217.210 ;
        RECT 674.995 216.150 675.425 216.935 ;
        RECT 675.825 216.110 680.955 217.020 ;
        RECT 681.500 216.995 681.780 217.275 ;
        RECT 686.620 217.020 686.790 217.210 ;
        RECT 680.975 216.150 681.405 216.935 ;
        RECT 681.805 216.110 686.935 217.020 ;
        RECT 687.480 216.995 687.760 217.275 ;
        RECT 692.600 217.020 692.770 217.210 ;
        RECT 686.955 216.150 687.385 216.935 ;
        RECT 687.785 216.110 692.915 217.020 ;
        RECT 693.460 216.995 693.740 217.275 ;
        RECT 698.580 217.020 698.750 217.210 ;
        RECT 692.935 216.150 693.365 216.935 ;
        RECT 693.765 216.110 698.895 217.020 ;
        RECT 699.440 216.995 699.720 217.275 ;
        RECT 704.560 217.020 704.730 217.210 ;
        RECT 698.915 216.150 699.345 216.935 ;
        RECT 699.745 216.110 704.875 217.020 ;
        RECT 705.420 216.995 705.700 217.275 ;
        RECT 710.540 217.020 710.710 217.210 ;
        RECT 704.895 216.150 705.325 216.935 ;
        RECT 705.725 216.110 710.855 217.020 ;
        RECT 711.400 216.995 711.680 217.275 ;
        RECT 716.520 217.020 716.690 217.210 ;
        RECT 710.875 216.150 711.305 216.935 ;
        RECT 711.705 216.110 716.835 217.020 ;
        RECT 717.380 216.995 717.660 217.275 ;
        RECT 722.500 217.020 722.670 217.210 ;
        RECT 716.855 216.150 717.285 216.935 ;
        RECT 717.685 216.110 722.815 217.020 ;
        RECT 723.360 216.995 723.640 217.275 ;
        RECT 728.480 217.020 728.650 217.210 ;
        RECT 722.835 216.150 723.265 216.935 ;
        RECT 723.665 216.110 728.795 217.020 ;
        RECT 729.340 216.995 729.620 217.275 ;
        RECT 734.460 217.020 734.630 217.210 ;
        RECT 728.815 216.150 729.245 216.935 ;
        RECT 729.645 216.110 734.775 217.020 ;
        RECT 735.320 216.995 735.600 217.275 ;
        RECT 740.440 217.020 740.610 217.210 ;
        RECT 734.795 216.150 735.225 216.935 ;
        RECT 735.625 216.110 740.755 217.020 ;
        RECT 741.300 216.995 741.580 217.275 ;
        RECT 746.420 217.020 746.590 217.210 ;
        RECT 740.775 216.150 741.205 216.935 ;
        RECT 741.605 216.110 746.735 217.020 ;
        RECT 747.280 216.995 747.560 217.275 ;
        RECT 752.400 217.020 752.570 217.210 ;
        RECT 746.755 216.150 747.185 216.935 ;
        RECT 747.585 216.110 752.715 217.020 ;
        RECT 753.260 216.995 753.540 217.275 ;
        RECT 758.380 217.020 758.550 217.210 ;
        RECT 752.735 216.150 753.165 216.935 ;
        RECT 753.565 216.110 758.695 217.020 ;
        RECT 759.240 216.995 759.520 217.275 ;
        RECT 764.360 217.020 764.530 217.210 ;
        RECT 758.715 216.150 759.145 216.935 ;
        RECT 759.545 216.110 764.675 217.020 ;
        RECT 765.220 216.995 765.500 217.275 ;
        RECT 770.340 217.020 770.510 217.210 ;
        RECT 764.695 216.150 765.125 216.935 ;
        RECT 765.525 216.110 770.655 217.020 ;
        RECT 771.200 216.995 771.480 217.275 ;
        RECT 776.320 217.020 776.490 217.210 ;
        RECT 770.675 216.150 771.105 216.935 ;
        RECT 771.505 216.110 776.635 217.020 ;
        RECT 777.180 216.995 777.460 217.275 ;
        RECT 782.300 217.020 782.470 217.210 ;
        RECT 776.655 216.150 777.085 216.935 ;
        RECT 777.485 216.110 782.615 217.020 ;
        RECT 783.160 216.995 783.440 217.275 ;
        RECT 788.280 217.020 788.450 217.210 ;
        RECT 782.635 216.150 783.065 216.935 ;
        RECT 783.465 216.110 788.595 217.020 ;
        RECT 789.140 216.995 789.420 217.275 ;
        RECT 794.260 217.020 794.430 217.210 ;
        RECT 788.615 216.150 789.045 216.935 ;
        RECT 789.445 216.110 794.575 217.020 ;
        RECT 2146.540 216.995 2146.820 217.275 ;
        RECT 2151.660 217.020 2151.830 217.210 ;
        RECT 794.595 216.150 795.025 216.935 ;
        RECT 2146.015 216.150 2146.445 216.935 ;
        RECT 2146.845 216.110 2151.975 217.020 ;
        RECT 2152.520 216.995 2152.800 217.275 ;
        RECT 2157.640 217.020 2157.810 217.210 ;
        RECT 2151.995 216.150 2152.425 216.935 ;
        RECT 2152.825 216.110 2157.955 217.020 ;
        RECT 2158.500 216.995 2158.780 217.275 ;
        RECT 2163.620 217.020 2163.790 217.210 ;
        RECT 2157.975 216.150 2158.405 216.935 ;
        RECT 2158.805 216.110 2163.935 217.020 ;
        RECT 2164.480 216.995 2164.760 217.275 ;
        RECT 2169.600 217.020 2169.770 217.210 ;
        RECT 2163.955 216.150 2164.385 216.935 ;
        RECT 2164.785 216.110 2169.915 217.020 ;
        RECT 2170.460 216.995 2170.740 217.275 ;
        RECT 2175.580 217.020 2175.750 217.210 ;
        RECT 2169.935 216.150 2170.365 216.935 ;
        RECT 2170.765 216.110 2175.895 217.020 ;
        RECT 2176.440 216.995 2176.720 217.275 ;
        RECT 2181.560 217.020 2181.730 217.210 ;
        RECT 2175.915 216.150 2176.345 216.935 ;
        RECT 2176.745 216.110 2181.875 217.020 ;
        RECT 2182.420 216.995 2182.700 217.275 ;
        RECT 2187.540 217.020 2187.710 217.210 ;
        RECT 2181.895 216.150 2182.325 216.935 ;
        RECT 2182.725 216.110 2187.855 217.020 ;
        RECT 2188.400 216.995 2188.680 217.275 ;
        RECT 2193.520 217.020 2193.690 217.210 ;
        RECT 2187.875 216.150 2188.305 216.935 ;
        RECT 2188.705 216.110 2193.835 217.020 ;
        RECT 2194.380 216.995 2194.660 217.275 ;
        RECT 2199.500 217.020 2199.670 217.210 ;
        RECT 2193.855 216.150 2194.285 216.935 ;
        RECT 2194.685 216.110 2199.815 217.020 ;
        RECT 2200.360 216.995 2200.640 217.275 ;
        RECT 2205.480 217.020 2205.650 217.210 ;
        RECT 2199.835 216.150 2200.265 216.935 ;
        RECT 2200.665 216.110 2205.795 217.020 ;
        RECT 2206.340 216.995 2206.620 217.275 ;
        RECT 2211.460 217.020 2211.630 217.210 ;
        RECT 2205.815 216.150 2206.245 216.935 ;
        RECT 2206.645 216.110 2211.775 217.020 ;
        RECT 2212.320 216.995 2212.600 217.275 ;
        RECT 2217.440 217.020 2217.610 217.210 ;
        RECT 2211.795 216.150 2212.225 216.935 ;
        RECT 2212.625 216.110 2217.755 217.020 ;
        RECT 2218.300 216.995 2218.580 217.275 ;
        RECT 2223.420 217.020 2223.590 217.210 ;
        RECT 2217.775 216.150 2218.205 216.935 ;
        RECT 2218.605 216.110 2223.735 217.020 ;
        RECT 2224.280 216.995 2224.560 217.275 ;
        RECT 2229.400 217.020 2229.570 217.210 ;
        RECT 2223.755 216.150 2224.185 216.935 ;
        RECT 2224.585 216.110 2229.715 217.020 ;
        RECT 2230.260 216.995 2230.540 217.275 ;
        RECT 2235.380 217.020 2235.550 217.210 ;
        RECT 2229.735 216.150 2230.165 216.935 ;
        RECT 2230.565 216.110 2235.695 217.020 ;
        RECT 2236.240 216.995 2236.520 217.275 ;
        RECT 2241.360 217.020 2241.530 217.210 ;
        RECT 2235.715 216.150 2236.145 216.935 ;
        RECT 2236.545 216.110 2241.675 217.020 ;
        RECT 2242.220 216.995 2242.500 217.275 ;
        RECT 2247.340 217.020 2247.510 217.210 ;
        RECT 2241.695 216.150 2242.125 216.935 ;
        RECT 2242.525 216.110 2247.655 217.020 ;
        RECT 2248.200 216.995 2248.480 217.275 ;
        RECT 2253.320 217.020 2253.490 217.210 ;
        RECT 2247.675 216.150 2248.105 216.935 ;
        RECT 2248.505 216.110 2253.635 217.020 ;
        RECT 2254.180 216.995 2254.460 217.275 ;
        RECT 2259.300 217.020 2259.470 217.210 ;
        RECT 2253.655 216.150 2254.085 216.935 ;
        RECT 2254.485 216.110 2259.615 217.020 ;
        RECT 2260.160 216.995 2260.440 217.275 ;
        RECT 2265.280 217.020 2265.450 217.210 ;
        RECT 2259.635 216.150 2260.065 216.935 ;
        RECT 2260.465 216.110 2265.595 217.020 ;
        RECT 2266.140 216.995 2266.420 217.275 ;
        RECT 2271.260 217.020 2271.430 217.210 ;
        RECT 2265.615 216.150 2266.045 216.935 ;
        RECT 2266.445 216.110 2271.575 217.020 ;
        RECT 2271.595 216.150 2272.025 216.935 ;
      LAYER nwell ;
        RECT 668.810 212.990 795.230 215.820 ;
        RECT 2145.810 212.990 2272.230 215.820 ;
      LAYER pwell ;
        RECT 669.015 211.875 669.445 212.660 ;
        RECT 674.995 211.875 675.425 212.660 ;
        RECT 669.540 211.555 669.820 211.835 ;
        RECT 675.445 211.790 680.575 212.700 ;
        RECT 680.975 211.875 681.405 212.660 ;
        RECT 681.425 211.790 686.555 212.700 ;
        RECT 686.955 211.875 687.385 212.660 ;
        RECT 687.405 211.790 692.535 212.700 ;
        RECT 692.935 211.875 693.365 212.660 ;
        RECT 693.385 211.790 698.515 212.700 ;
        RECT 698.915 211.875 699.345 212.660 ;
        RECT 699.365 211.790 704.495 212.700 ;
        RECT 704.895 211.875 705.325 212.660 ;
        RECT 705.345 211.790 710.475 212.700 ;
        RECT 710.875 211.875 711.305 212.660 ;
        RECT 711.325 211.790 716.455 212.700 ;
        RECT 716.855 211.875 717.285 212.660 ;
        RECT 717.305 211.790 722.435 212.700 ;
        RECT 722.835 211.875 723.265 212.660 ;
        RECT 723.285 211.790 728.415 212.700 ;
        RECT 728.815 211.875 729.245 212.660 ;
        RECT 729.265 211.790 734.395 212.700 ;
        RECT 734.795 211.875 735.225 212.660 ;
        RECT 735.245 211.790 740.375 212.700 ;
        RECT 740.775 211.875 741.205 212.660 ;
        RECT 741.225 211.790 746.355 212.700 ;
        RECT 746.755 211.875 747.185 212.660 ;
        RECT 747.205 211.790 752.335 212.700 ;
        RECT 752.735 211.875 753.165 212.660 ;
        RECT 753.185 211.790 758.315 212.700 ;
        RECT 758.715 211.875 759.145 212.660 ;
        RECT 759.165 211.790 764.295 212.700 ;
        RECT 764.695 211.875 765.125 212.660 ;
        RECT 765.145 211.790 770.275 212.700 ;
        RECT 770.675 211.875 771.105 212.660 ;
        RECT 771.125 211.790 776.255 212.700 ;
        RECT 776.655 211.875 777.085 212.660 ;
        RECT 777.105 211.790 782.235 212.700 ;
        RECT 782.635 211.875 783.065 212.660 ;
        RECT 783.085 211.790 788.215 212.700 ;
        RECT 788.615 211.875 789.045 212.660 ;
        RECT 789.445 211.790 794.575 212.700 ;
        RECT 794.595 211.875 795.025 212.660 ;
        RECT 2146.015 211.875 2146.445 212.660 ;
        RECT 2151.995 211.875 2152.425 212.660 ;
        RECT 675.590 211.600 675.760 211.790 ;
        RECT 681.570 211.600 681.740 211.790 ;
        RECT 687.550 211.600 687.720 211.790 ;
        RECT 693.530 211.600 693.700 211.790 ;
        RECT 699.510 211.600 699.680 211.790 ;
        RECT 705.490 211.600 705.660 211.790 ;
        RECT 711.470 211.600 711.640 211.790 ;
        RECT 717.450 211.600 717.620 211.790 ;
        RECT 723.430 211.600 723.600 211.790 ;
        RECT 729.410 211.600 729.580 211.790 ;
        RECT 735.390 211.600 735.560 211.790 ;
        RECT 741.370 211.600 741.540 211.790 ;
        RECT 747.350 211.600 747.520 211.790 ;
        RECT 753.330 211.600 753.500 211.790 ;
        RECT 759.310 211.600 759.480 211.790 ;
        RECT 765.290 211.600 765.460 211.790 ;
        RECT 771.270 211.600 771.440 211.790 ;
        RECT 777.250 211.600 777.420 211.790 ;
        RECT 783.230 211.600 783.400 211.790 ;
        RECT 794.260 211.600 794.430 211.790 ;
        RECT 2146.540 211.555 2146.820 211.835 ;
        RECT 2152.445 211.790 2157.575 212.700 ;
        RECT 2157.975 211.875 2158.405 212.660 ;
        RECT 2158.425 211.790 2163.555 212.700 ;
        RECT 2163.955 211.875 2164.385 212.660 ;
        RECT 2164.405 211.790 2169.535 212.700 ;
        RECT 2169.935 211.875 2170.365 212.660 ;
        RECT 2170.385 211.790 2175.515 212.700 ;
        RECT 2175.915 211.875 2176.345 212.660 ;
        RECT 2176.365 211.790 2181.495 212.700 ;
        RECT 2181.895 211.875 2182.325 212.660 ;
        RECT 2182.345 211.790 2187.475 212.700 ;
        RECT 2187.875 211.875 2188.305 212.660 ;
        RECT 2188.325 211.790 2193.455 212.700 ;
        RECT 2193.855 211.875 2194.285 212.660 ;
        RECT 2194.305 211.790 2199.435 212.700 ;
        RECT 2199.835 211.875 2200.265 212.660 ;
        RECT 2200.285 211.790 2205.415 212.700 ;
        RECT 2205.815 211.875 2206.245 212.660 ;
        RECT 2206.265 211.790 2211.395 212.700 ;
        RECT 2211.795 211.875 2212.225 212.660 ;
        RECT 2212.245 211.790 2217.375 212.700 ;
        RECT 2217.775 211.875 2218.205 212.660 ;
        RECT 2218.225 211.790 2223.355 212.700 ;
        RECT 2223.755 211.875 2224.185 212.660 ;
        RECT 2224.205 211.790 2229.335 212.700 ;
        RECT 2229.735 211.875 2230.165 212.660 ;
        RECT 2230.185 211.790 2235.315 212.700 ;
        RECT 2235.715 211.875 2236.145 212.660 ;
        RECT 2236.165 211.790 2241.295 212.700 ;
        RECT 2241.695 211.875 2242.125 212.660 ;
        RECT 2242.145 211.790 2247.275 212.700 ;
        RECT 2247.675 211.875 2248.105 212.660 ;
        RECT 2248.125 211.790 2253.255 212.700 ;
        RECT 2253.655 211.875 2254.085 212.660 ;
        RECT 2254.105 211.790 2259.235 212.700 ;
        RECT 2259.635 211.875 2260.065 212.660 ;
        RECT 2260.085 211.790 2265.215 212.700 ;
        RECT 2265.615 211.875 2266.045 212.660 ;
        RECT 2266.445 211.790 2271.575 212.700 ;
        RECT 2271.595 211.875 2272.025 212.660 ;
        RECT 2152.590 211.600 2152.760 211.790 ;
        RECT 2158.570 211.600 2158.740 211.790 ;
        RECT 2164.550 211.600 2164.720 211.790 ;
        RECT 2170.530 211.600 2170.700 211.790 ;
        RECT 2176.510 211.600 2176.680 211.790 ;
        RECT 2182.490 211.600 2182.660 211.790 ;
        RECT 2188.470 211.600 2188.640 211.790 ;
        RECT 2194.450 211.600 2194.620 211.790 ;
        RECT 2200.430 211.600 2200.600 211.790 ;
        RECT 2206.410 211.600 2206.580 211.790 ;
        RECT 2212.390 211.600 2212.560 211.790 ;
        RECT 2218.370 211.600 2218.540 211.790 ;
        RECT 2224.350 211.600 2224.520 211.790 ;
        RECT 2230.330 211.600 2230.500 211.790 ;
        RECT 2236.310 211.600 2236.480 211.790 ;
        RECT 2242.290 211.600 2242.460 211.790 ;
        RECT 2248.270 211.600 2248.440 211.790 ;
        RECT 2254.250 211.600 2254.420 211.790 ;
        RECT 2260.230 211.600 2260.400 211.790 ;
        RECT 2271.260 211.600 2271.430 211.790 ;
      LAYER li1 ;
        RECT 2082.830 4987.615 2082.975 4987.785 ;
        RECT 2083.145 4987.615 2083.435 4987.785 ;
        RECT 2083.605 4987.615 2083.895 4987.785 ;
        RECT 2084.065 4987.615 2084.355 4987.785 ;
        RECT 2084.525 4987.615 2084.815 4987.785 ;
        RECT 2084.985 4987.615 2085.275 4987.785 ;
        RECT 2085.445 4987.615 2085.735 4987.785 ;
        RECT 2085.905 4987.615 2086.195 4987.785 ;
        RECT 2086.365 4987.615 2086.655 4987.785 ;
        RECT 2086.825 4987.615 2087.115 4987.785 ;
        RECT 2087.285 4987.615 2087.575 4987.785 ;
        RECT 2087.745 4987.615 2088.035 4987.785 ;
        RECT 2088.205 4987.615 2088.495 4987.785 ;
        RECT 2088.665 4987.615 2088.955 4987.785 ;
        RECT 2089.125 4987.615 2089.270 4987.785 ;
        RECT 2082.915 4986.890 2083.205 4987.615 ;
        RECT 2083.765 4986.815 2084.095 4987.615 ;
        RECT 2084.605 4987.135 2084.935 4987.615 ;
        RECT 2085.445 4987.135 2085.775 4987.615 ;
        RECT 2086.285 4987.135 2086.615 4987.615 ;
        RECT 2087.125 4987.135 2087.455 4987.615 ;
        RECT 2087.625 4986.965 2087.795 4987.440 ;
        RECT 2087.965 4987.135 2088.295 4987.615 ;
        RECT 2088.465 4986.965 2088.635 4987.445 ;
        RECT 2087.215 4986.795 2088.635 4986.965 ;
        RECT 2088.895 4986.890 2089.185 4987.615 ;
        RECT 3309.835 4987.205 3309.980 4987.375 ;
        RECT 3310.150 4987.205 3310.440 4987.375 ;
        RECT 3310.610 4987.205 3310.900 4987.375 ;
        RECT 3311.070 4987.205 3311.360 4987.375 ;
        RECT 3311.530 4987.205 3311.820 4987.375 ;
        RECT 3311.990 4987.205 3312.280 4987.375 ;
        RECT 3312.450 4987.205 3312.740 4987.375 ;
        RECT 3312.910 4987.205 3313.200 4987.375 ;
        RECT 3313.370 4987.205 3313.660 4987.375 ;
        RECT 3313.830 4987.205 3314.120 4987.375 ;
        RECT 3314.290 4987.205 3314.580 4987.375 ;
        RECT 3314.750 4987.205 3315.040 4987.375 ;
        RECT 3315.210 4987.205 3315.500 4987.375 ;
        RECT 3315.670 4987.205 3315.960 4987.375 ;
        RECT 3316.130 4987.205 3316.420 4987.375 ;
        RECT 3316.590 4987.205 3316.880 4987.375 ;
        RECT 3317.050 4987.205 3317.340 4987.375 ;
        RECT 3317.510 4987.205 3317.800 4987.375 ;
        RECT 3317.970 4987.205 3318.260 4987.375 ;
        RECT 3318.430 4987.205 3318.720 4987.375 ;
        RECT 3318.890 4987.205 3319.180 4987.375 ;
        RECT 3319.350 4987.205 3319.640 4987.375 ;
        RECT 3319.810 4987.205 3320.100 4987.375 ;
        RECT 3320.270 4987.205 3320.560 4987.375 ;
        RECT 3320.730 4987.205 3321.020 4987.375 ;
        RECT 3321.190 4987.205 3321.480 4987.375 ;
        RECT 3321.650 4987.205 3321.940 4987.375 ;
        RECT 3322.110 4987.205 3322.400 4987.375 ;
        RECT 3322.570 4987.205 3322.860 4987.375 ;
        RECT 3323.030 4987.205 3323.320 4987.375 ;
        RECT 3323.490 4987.205 3323.780 4987.375 ;
        RECT 3323.950 4987.205 3324.240 4987.375 ;
        RECT 3324.410 4987.205 3324.700 4987.375 ;
        RECT 3324.870 4987.205 3325.160 4987.375 ;
        RECT 3325.330 4987.205 3325.620 4987.375 ;
        RECT 3325.790 4987.205 3326.080 4987.375 ;
        RECT 3326.250 4987.205 3326.540 4987.375 ;
        RECT 3326.710 4987.205 3327.000 4987.375 ;
        RECT 3327.170 4987.205 3327.460 4987.375 ;
        RECT 3327.630 4987.205 3327.920 4987.375 ;
        RECT 3328.090 4987.205 3328.380 4987.375 ;
        RECT 3328.550 4987.205 3328.840 4987.375 ;
        RECT 3329.010 4987.205 3329.300 4987.375 ;
        RECT 3329.470 4987.205 3329.760 4987.375 ;
        RECT 3329.930 4987.205 3330.220 4987.375 ;
        RECT 3330.390 4987.205 3330.680 4987.375 ;
        RECT 3330.850 4987.205 3331.140 4987.375 ;
        RECT 3331.310 4987.205 3331.600 4987.375 ;
        RECT 3331.770 4987.205 3332.060 4987.375 ;
        RECT 3332.230 4987.205 3332.520 4987.375 ;
        RECT 3332.690 4987.205 3332.980 4987.375 ;
        RECT 3333.150 4987.205 3333.440 4987.375 ;
        RECT 3333.610 4987.205 3333.900 4987.375 ;
        RECT 3334.070 4987.205 3334.215 4987.375 ;
        RECT 2087.215 4986.625 2087.390 4986.795 ;
        RECT 2084.765 4986.455 2087.390 4986.625 ;
        RECT 2087.215 4986.255 2087.390 4986.455 ;
      LAYER li1 ;
        RECT 2087.570 4986.425 2088.670 4986.625 ;
      LAYER li1 ;
        RECT 3309.920 4986.480 3310.210 4987.205 ;
        RECT 3310.770 4986.405 3311.100 4987.205 ;
      LAYER li1 ;
        RECT 3311.270 4986.555 3311.440 4987.035 ;
      LAYER li1 ;
        RECT 3311.610 4986.725 3311.940 4987.205 ;
      LAYER li1 ;
        RECT 3312.110 4986.555 3312.280 4987.035 ;
      LAYER li1 ;
        RECT 3312.450 4986.725 3312.780 4987.205 ;
      LAYER li1 ;
        RECT 3312.950 4986.555 3313.120 4987.035 ;
      LAYER li1 ;
        RECT 3313.290 4986.725 3313.620 4987.205 ;
      LAYER li1 ;
        RECT 3313.790 4986.555 3313.960 4987.035 ;
      LAYER li1 ;
        RECT 3314.130 4986.725 3314.460 4987.205 ;
        RECT 3314.630 4986.555 3314.800 4987.030 ;
        RECT 3314.970 4986.725 3315.300 4987.205 ;
        RECT 3315.470 4986.555 3315.640 4987.035 ;
      LAYER li1 ;
        RECT 3311.270 4986.385 3313.960 4986.555 ;
      LAYER li1 ;
        RECT 3314.220 4986.385 3315.640 4986.555 ;
        RECT 3315.900 4986.480 3316.190 4987.205 ;
        RECT 3316.750 4986.405 3317.080 4987.205 ;
        RECT 3317.590 4986.725 3317.920 4987.205 ;
        RECT 3318.430 4986.725 3318.760 4987.205 ;
        RECT 3319.270 4986.725 3319.600 4987.205 ;
        RECT 3320.110 4986.725 3320.440 4987.205 ;
        RECT 3320.610 4986.555 3320.780 4987.030 ;
        RECT 3320.950 4986.725 3321.280 4987.205 ;
        RECT 3321.450 4986.555 3321.620 4987.035 ;
        RECT 3320.200 4986.385 3321.620 4986.555 ;
        RECT 3321.880 4986.480 3322.170 4987.205 ;
        RECT 3322.730 4986.405 3323.060 4987.205 ;
        RECT 3323.570 4986.725 3323.900 4987.205 ;
        RECT 3324.410 4986.725 3324.740 4987.205 ;
        RECT 3325.250 4986.725 3325.580 4987.205 ;
        RECT 3326.090 4986.725 3326.420 4987.205 ;
        RECT 3326.590 4986.555 3326.760 4987.030 ;
        RECT 3326.930 4986.725 3327.260 4987.205 ;
        RECT 3327.430 4986.555 3327.600 4987.035 ;
        RECT 3326.180 4986.385 3327.600 4986.555 ;
        RECT 3327.860 4986.480 3328.150 4987.205 ;
        RECT 3328.710 4986.405 3329.040 4987.205 ;
        RECT 3329.550 4986.725 3329.880 4987.205 ;
        RECT 3330.390 4986.725 3330.720 4987.205 ;
        RECT 3331.230 4986.725 3331.560 4987.205 ;
        RECT 3332.070 4986.725 3332.400 4987.205 ;
        RECT 3332.570 4986.555 3332.740 4987.030 ;
        RECT 3332.910 4986.725 3333.240 4987.205 ;
        RECT 3333.410 4986.555 3333.580 4987.035 ;
        RECT 3332.160 4986.385 3333.580 4986.555 ;
        RECT 3333.840 4986.480 3334.130 4987.205 ;
        RECT 834.650 4985.990 834.795 4986.160 ;
        RECT 834.965 4985.990 835.255 4986.160 ;
        RECT 835.425 4985.990 835.715 4986.160 ;
        RECT 835.885 4985.990 836.175 4986.160 ;
        RECT 836.345 4985.990 836.635 4986.160 ;
        RECT 836.805 4985.990 837.095 4986.160 ;
        RECT 837.265 4985.990 837.555 4986.160 ;
        RECT 837.725 4985.990 838.015 4986.160 ;
        RECT 838.185 4985.990 838.475 4986.160 ;
        RECT 838.645 4985.990 838.935 4986.160 ;
        RECT 839.105 4985.990 839.395 4986.160 ;
        RECT 839.565 4985.990 839.855 4986.160 ;
        RECT 840.025 4985.990 840.315 4986.160 ;
        RECT 840.485 4985.990 840.775 4986.160 ;
        RECT 840.945 4985.990 841.235 4986.160 ;
        RECT 841.405 4985.990 841.695 4986.160 ;
        RECT 841.865 4985.990 842.155 4986.160 ;
        RECT 842.325 4985.990 842.615 4986.160 ;
        RECT 842.785 4985.990 843.075 4986.160 ;
        RECT 843.245 4985.990 843.535 4986.160 ;
        RECT 843.705 4985.990 843.995 4986.160 ;
        RECT 844.165 4985.990 844.455 4986.160 ;
        RECT 844.625 4985.990 844.915 4986.160 ;
        RECT 845.085 4985.990 845.375 4986.160 ;
        RECT 845.545 4985.990 845.835 4986.160 ;
        RECT 846.005 4985.990 846.295 4986.160 ;
        RECT 846.465 4985.990 846.755 4986.160 ;
        RECT 846.925 4985.990 847.215 4986.160 ;
        RECT 847.385 4985.990 847.675 4986.160 ;
        RECT 847.845 4985.990 848.135 4986.160 ;
        RECT 848.305 4985.990 848.595 4986.160 ;
        RECT 848.765 4985.990 849.055 4986.160 ;
        RECT 849.225 4985.990 849.515 4986.160 ;
        RECT 849.685 4985.990 849.975 4986.160 ;
        RECT 850.145 4985.990 850.435 4986.160 ;
        RECT 850.605 4985.990 850.895 4986.160 ;
        RECT 851.065 4985.990 851.355 4986.160 ;
        RECT 851.525 4985.990 851.815 4986.160 ;
        RECT 851.985 4985.990 852.275 4986.160 ;
        RECT 852.445 4985.990 852.735 4986.160 ;
        RECT 852.905 4985.990 853.050 4986.160 ;
        RECT 834.735 4985.265 835.025 4985.990 ;
        RECT 835.285 4985.340 835.455 4985.820 ;
        RECT 835.625 4985.510 835.955 4985.990 ;
        RECT 836.125 4985.340 836.295 4985.815 ;
        RECT 836.465 4985.510 836.795 4985.990 ;
        RECT 837.305 4985.510 837.635 4985.990 ;
        RECT 838.145 4985.510 838.475 4985.990 ;
        RECT 838.985 4985.510 839.315 4985.990 ;
        RECT 835.285 4985.170 836.705 4985.340 ;
        RECT 839.825 4985.190 840.155 4985.990 ;
        RECT 840.715 4985.265 841.005 4985.990 ;
        RECT 841.265 4985.340 841.435 4985.820 ;
        RECT 841.605 4985.510 841.935 4985.990 ;
        RECT 842.105 4985.340 842.275 4985.815 ;
        RECT 842.445 4985.510 842.775 4985.990 ;
        RECT 843.285 4985.510 843.615 4985.990 ;
        RECT 844.125 4985.510 844.455 4985.990 ;
        RECT 844.965 4985.510 845.295 4985.990 ;
        RECT 841.265 4985.170 842.685 4985.340 ;
        RECT 845.805 4985.190 846.135 4985.990 ;
        RECT 846.695 4985.265 846.985 4985.990 ;
        RECT 847.245 4985.340 847.415 4985.820 ;
        RECT 847.585 4985.510 847.915 4985.990 ;
        RECT 848.085 4985.340 848.255 4985.815 ;
        RECT 848.425 4985.510 848.755 4985.990 ;
        RECT 849.265 4985.510 849.595 4985.990 ;
        RECT 850.105 4985.510 850.435 4985.990 ;
        RECT 850.945 4985.510 851.275 4985.990 ;
        RECT 847.245 4985.170 848.665 4985.340 ;
        RECT 851.785 4985.190 852.115 4985.990 ;
        RECT 852.675 4985.265 852.965 4985.990 ;
        RECT 836.530 4985.000 836.705 4985.170 ;
        RECT 842.510 4985.000 842.685 4985.170 ;
        RECT 848.490 4985.000 848.665 4985.170 ;
        RECT 2082.915 4985.065 2083.205 4986.230 ;
        RECT 2083.765 4985.065 2084.095 4986.215 ;
        RECT 2087.215 4986.085 2088.715 4986.255 ;
        RECT 2084.605 4985.065 2084.935 4985.865 ;
        RECT 2085.445 4985.065 2085.775 4985.865 ;
        RECT 2086.285 4985.065 2086.615 4985.865 ;
        RECT 2087.205 4985.065 2087.375 4985.865 ;
        RECT 2087.545 4985.235 2087.875 4986.085 ;
        RECT 2088.045 4985.065 2088.215 4985.865 ;
        RECT 2088.385 4985.235 2088.715 4986.085 ;
        RECT 2088.895 4985.065 2089.185 4986.230 ;
      LAYER li1 ;
        RECT 3311.270 4985.845 3311.525 4986.385 ;
      LAYER li1 ;
        RECT 3314.220 4986.215 3314.395 4986.385 ;
        RECT 3320.200 4986.215 3320.375 4986.385 ;
        RECT 3326.180 4986.215 3326.355 4986.385 ;
        RECT 3332.160 4986.215 3332.335 4986.385 ;
        RECT 3311.770 4986.045 3314.395 4986.215 ;
        RECT 3314.220 4985.845 3314.395 4986.045 ;
      LAYER li1 ;
        RECT 3314.575 4986.015 3315.675 4986.215 ;
      LAYER li1 ;
        RECT 3317.750 4986.045 3320.375 4986.215 ;
        RECT 3320.200 4985.845 3320.375 4986.045 ;
      LAYER li1 ;
        RECT 3320.555 4986.015 3321.655 4986.215 ;
      LAYER li1 ;
        RECT 3323.730 4986.045 3326.355 4986.215 ;
        RECT 3326.180 4985.845 3326.355 4986.045 ;
      LAYER li1 ;
        RECT 3326.535 4986.015 3327.635 4986.215 ;
      LAYER li1 ;
        RECT 3329.710 4986.045 3332.335 4986.215 ;
        RECT 3332.160 4985.845 3332.335 4986.045 ;
      LAYER li1 ;
        RECT 3332.515 4986.015 3333.615 4986.215 ;
        RECT 835.250 4984.800 836.350 4985.000 ;
      LAYER li1 ;
        RECT 836.530 4984.830 839.155 4985.000 ;
        RECT 836.530 4984.630 836.705 4984.830 ;
      LAYER li1 ;
        RECT 841.230 4984.800 842.330 4985.000 ;
      LAYER li1 ;
        RECT 842.510 4984.830 845.135 4985.000 ;
        RECT 842.510 4984.630 842.685 4984.830 ;
      LAYER li1 ;
        RECT 847.210 4984.800 848.310 4985.000 ;
      LAYER li1 ;
        RECT 848.490 4984.830 851.115 4985.000 ;
        RECT 2082.830 4984.895 2082.975 4985.065 ;
        RECT 2083.145 4984.895 2083.435 4985.065 ;
        RECT 2083.605 4984.895 2083.895 4985.065 ;
        RECT 2084.065 4984.895 2084.355 4985.065 ;
        RECT 2084.525 4984.895 2084.815 4985.065 ;
        RECT 2084.985 4984.895 2085.275 4985.065 ;
        RECT 2085.445 4984.895 2085.735 4985.065 ;
        RECT 2085.905 4984.895 2086.195 4985.065 ;
        RECT 2086.365 4984.895 2086.655 4985.065 ;
        RECT 2086.825 4984.895 2087.115 4985.065 ;
        RECT 2087.285 4984.895 2087.575 4985.065 ;
        RECT 2087.745 4984.895 2088.035 4985.065 ;
        RECT 2088.205 4984.895 2088.495 4985.065 ;
        RECT 2088.665 4984.895 2088.955 4985.065 ;
        RECT 2089.125 4984.895 2089.270 4985.065 ;
        RECT 848.490 4984.630 848.665 4984.830 ;
        RECT 834.735 4983.440 835.025 4984.605 ;
        RECT 835.205 4984.460 836.705 4984.630 ;
        RECT 835.205 4983.610 835.535 4984.460 ;
        RECT 835.705 4983.440 835.875 4984.240 ;
        RECT 836.045 4983.610 836.375 4984.460 ;
        RECT 836.545 4983.440 836.715 4984.240 ;
        RECT 837.305 4983.440 837.635 4984.240 ;
        RECT 838.145 4983.440 838.475 4984.240 ;
        RECT 838.985 4983.440 839.315 4984.240 ;
        RECT 839.825 4983.440 840.155 4984.590 ;
        RECT 840.715 4983.440 841.005 4984.605 ;
        RECT 841.185 4984.460 842.685 4984.630 ;
        RECT 841.185 4983.610 841.515 4984.460 ;
        RECT 841.685 4983.440 841.855 4984.240 ;
        RECT 842.025 4983.610 842.355 4984.460 ;
        RECT 842.525 4983.440 842.695 4984.240 ;
        RECT 843.285 4983.440 843.615 4984.240 ;
        RECT 844.125 4983.440 844.455 4984.240 ;
        RECT 844.965 4983.440 845.295 4984.240 ;
        RECT 845.805 4983.440 846.135 4984.590 ;
        RECT 846.695 4983.440 846.985 4984.605 ;
        RECT 847.165 4984.460 848.665 4984.630 ;
        RECT 847.165 4983.610 847.495 4984.460 ;
        RECT 847.665 4983.440 847.835 4984.240 ;
        RECT 848.005 4983.610 848.335 4984.460 ;
        RECT 848.505 4983.440 848.675 4984.240 ;
        RECT 849.265 4983.440 849.595 4984.240 ;
        RECT 850.105 4983.440 850.435 4984.240 ;
        RECT 850.945 4983.440 851.275 4984.240 ;
        RECT 851.785 4983.440 852.115 4984.590 ;
        RECT 852.675 4983.440 852.965 4984.605 ;
        RECT 2082.915 4983.730 2083.205 4984.895 ;
        RECT 2083.385 4983.875 2083.715 4984.725 ;
        RECT 2083.885 4984.095 2084.055 4984.895 ;
        RECT 2084.225 4983.875 2084.555 4984.725 ;
        RECT 2084.725 4984.095 2084.895 4984.895 ;
      LAYER li1 ;
        RECT 2085.145 4983.875 2085.315 4984.725 ;
      LAYER li1 ;
        RECT 2085.485 4984.095 2085.815 4984.895 ;
      LAYER li1 ;
        RECT 2085.985 4983.875 2086.155 4984.725 ;
      LAYER li1 ;
        RECT 2086.325 4984.095 2086.655 4984.895 ;
      LAYER li1 ;
        RECT 2086.825 4983.875 2086.995 4984.725 ;
      LAYER li1 ;
        RECT 2087.165 4984.095 2087.495 4984.895 ;
      LAYER li1 ;
        RECT 2087.665 4983.875 2087.835 4984.725 ;
      LAYER li1 ;
        RECT 2083.385 4983.705 2084.885 4983.875 ;
      LAYER li1 ;
        RECT 2085.145 4983.705 2087.835 4983.875 ;
      LAYER li1 ;
        RECT 2088.005 4983.745 2088.335 4984.895 ;
        RECT 2088.895 4983.730 2089.185 4984.895 ;
        RECT 3309.920 4984.655 3310.210 4985.820 ;
        RECT 3310.770 4984.655 3311.100 4985.805 ;
      LAYER li1 ;
        RECT 3311.270 4985.675 3313.960 4985.845 ;
      LAYER li1 ;
        RECT 3314.220 4985.675 3315.720 4985.845 ;
      LAYER li1 ;
        RECT 3311.270 4984.825 3311.440 4985.675 ;
      LAYER li1 ;
        RECT 3311.610 4984.655 3311.940 4985.455 ;
      LAYER li1 ;
        RECT 3312.110 4984.825 3312.280 4985.675 ;
      LAYER li1 ;
        RECT 3312.450 4984.655 3312.780 4985.455 ;
      LAYER li1 ;
        RECT 3312.950 4984.825 3313.120 4985.675 ;
      LAYER li1 ;
        RECT 3313.290 4984.655 3313.620 4985.455 ;
      LAYER li1 ;
        RECT 3313.790 4984.825 3313.960 4985.675 ;
      LAYER li1 ;
        RECT 3314.210 4984.655 3314.380 4985.455 ;
        RECT 3314.550 4984.825 3314.880 4985.675 ;
        RECT 3315.050 4984.655 3315.220 4985.455 ;
        RECT 3315.390 4984.825 3315.720 4985.675 ;
        RECT 3315.900 4984.655 3316.190 4985.820 ;
        RECT 3316.750 4984.655 3317.080 4985.805 ;
        RECT 3320.200 4985.675 3321.700 4985.845 ;
        RECT 3317.590 4984.655 3317.920 4985.455 ;
        RECT 3318.430 4984.655 3318.760 4985.455 ;
        RECT 3319.270 4984.655 3319.600 4985.455 ;
        RECT 3320.190 4984.655 3320.360 4985.455 ;
        RECT 3320.530 4984.825 3320.860 4985.675 ;
        RECT 3321.030 4984.655 3321.200 4985.455 ;
        RECT 3321.370 4984.825 3321.700 4985.675 ;
        RECT 3321.880 4984.655 3322.170 4985.820 ;
        RECT 3322.730 4984.655 3323.060 4985.805 ;
        RECT 3326.180 4985.675 3327.680 4985.845 ;
        RECT 3323.570 4984.655 3323.900 4985.455 ;
        RECT 3324.410 4984.655 3324.740 4985.455 ;
        RECT 3325.250 4984.655 3325.580 4985.455 ;
        RECT 3326.170 4984.655 3326.340 4985.455 ;
        RECT 3326.510 4984.825 3326.840 4985.675 ;
        RECT 3327.010 4984.655 3327.180 4985.455 ;
        RECT 3327.350 4984.825 3327.680 4985.675 ;
        RECT 3327.860 4984.655 3328.150 4985.820 ;
        RECT 3328.710 4984.655 3329.040 4985.805 ;
        RECT 3332.160 4985.675 3333.660 4985.845 ;
        RECT 3329.550 4984.655 3329.880 4985.455 ;
        RECT 3330.390 4984.655 3330.720 4985.455 ;
        RECT 3331.230 4984.655 3331.560 4985.455 ;
        RECT 3332.150 4984.655 3332.320 4985.455 ;
        RECT 3332.490 4984.825 3332.820 4985.675 ;
        RECT 3332.990 4984.655 3333.160 4985.455 ;
        RECT 3333.330 4984.825 3333.660 4985.675 ;
        RECT 3333.840 4984.655 3334.130 4985.820 ;
        RECT 3309.835 4984.485 3309.980 4984.655 ;
        RECT 3310.150 4984.485 3310.440 4984.655 ;
        RECT 3310.610 4984.485 3310.900 4984.655 ;
        RECT 3311.070 4984.485 3311.360 4984.655 ;
        RECT 3311.530 4984.485 3311.820 4984.655 ;
        RECT 3311.990 4984.485 3312.280 4984.655 ;
        RECT 3312.450 4984.485 3312.740 4984.655 ;
        RECT 3312.910 4984.485 3313.200 4984.655 ;
        RECT 3313.370 4984.485 3313.660 4984.655 ;
        RECT 3313.830 4984.485 3314.120 4984.655 ;
        RECT 3314.290 4984.485 3314.580 4984.655 ;
        RECT 3314.750 4984.485 3315.040 4984.655 ;
        RECT 3315.210 4984.485 3315.500 4984.655 ;
        RECT 3315.670 4984.485 3315.960 4984.655 ;
        RECT 3316.130 4984.485 3316.420 4984.655 ;
        RECT 3316.590 4984.485 3316.880 4984.655 ;
        RECT 3317.050 4984.485 3317.340 4984.655 ;
        RECT 3317.510 4984.485 3317.800 4984.655 ;
        RECT 3317.970 4984.485 3318.260 4984.655 ;
        RECT 3318.430 4984.485 3318.720 4984.655 ;
        RECT 3318.890 4984.485 3319.180 4984.655 ;
        RECT 3319.350 4984.485 3319.640 4984.655 ;
        RECT 3319.810 4984.485 3320.100 4984.655 ;
        RECT 3320.270 4984.485 3320.560 4984.655 ;
        RECT 3320.730 4984.485 3321.020 4984.655 ;
        RECT 3321.190 4984.485 3321.480 4984.655 ;
        RECT 3321.650 4984.485 3321.940 4984.655 ;
        RECT 3322.110 4984.485 3322.400 4984.655 ;
        RECT 3322.570 4984.485 3322.860 4984.655 ;
        RECT 3323.030 4984.485 3323.320 4984.655 ;
        RECT 3323.490 4984.485 3323.780 4984.655 ;
        RECT 3323.950 4984.485 3324.240 4984.655 ;
        RECT 3324.410 4984.485 3324.700 4984.655 ;
        RECT 3324.870 4984.485 3325.160 4984.655 ;
        RECT 3325.330 4984.485 3325.620 4984.655 ;
        RECT 3325.790 4984.485 3326.080 4984.655 ;
        RECT 3326.250 4984.485 3326.540 4984.655 ;
        RECT 3326.710 4984.485 3327.000 4984.655 ;
        RECT 3327.170 4984.485 3327.460 4984.655 ;
        RECT 3327.630 4984.485 3327.920 4984.655 ;
        RECT 3328.090 4984.485 3328.380 4984.655 ;
        RECT 3328.550 4984.485 3328.840 4984.655 ;
        RECT 3329.010 4984.485 3329.300 4984.655 ;
        RECT 3329.470 4984.485 3329.760 4984.655 ;
        RECT 3329.930 4984.485 3330.220 4984.655 ;
        RECT 3330.390 4984.485 3330.680 4984.655 ;
        RECT 3330.850 4984.485 3331.140 4984.655 ;
        RECT 3331.310 4984.485 3331.600 4984.655 ;
        RECT 3331.770 4984.485 3332.060 4984.655 ;
        RECT 3332.230 4984.485 3332.520 4984.655 ;
        RECT 3332.690 4984.485 3332.980 4984.655 ;
        RECT 3333.150 4984.485 3333.440 4984.655 ;
        RECT 3333.610 4984.485 3333.900 4984.655 ;
        RECT 3334.070 4984.485 3334.215 4984.655 ;
        RECT 2084.710 4983.505 2084.885 4983.705 ;
        RECT 834.650 4983.270 834.795 4983.440 ;
        RECT 834.965 4983.270 835.255 4983.440 ;
        RECT 835.425 4983.270 835.715 4983.440 ;
        RECT 835.885 4983.270 836.175 4983.440 ;
        RECT 836.345 4983.270 836.635 4983.440 ;
        RECT 836.805 4983.270 837.095 4983.440 ;
        RECT 837.265 4983.270 837.555 4983.440 ;
        RECT 837.725 4983.270 838.015 4983.440 ;
        RECT 838.185 4983.270 838.475 4983.440 ;
        RECT 838.645 4983.270 838.935 4983.440 ;
        RECT 839.105 4983.270 839.395 4983.440 ;
        RECT 839.565 4983.270 839.855 4983.440 ;
        RECT 840.025 4983.270 840.315 4983.440 ;
        RECT 840.485 4983.270 840.775 4983.440 ;
        RECT 840.945 4983.270 841.235 4983.440 ;
        RECT 841.405 4983.270 841.695 4983.440 ;
        RECT 841.865 4983.270 842.155 4983.440 ;
        RECT 842.325 4983.270 842.615 4983.440 ;
        RECT 842.785 4983.270 843.075 4983.440 ;
        RECT 843.245 4983.270 843.535 4983.440 ;
        RECT 843.705 4983.270 843.995 4983.440 ;
        RECT 844.165 4983.270 844.455 4983.440 ;
        RECT 844.625 4983.270 844.915 4983.440 ;
        RECT 845.085 4983.270 845.375 4983.440 ;
        RECT 845.545 4983.270 845.835 4983.440 ;
        RECT 846.005 4983.270 846.295 4983.440 ;
        RECT 846.465 4983.270 846.755 4983.440 ;
        RECT 846.925 4983.270 847.215 4983.440 ;
        RECT 847.385 4983.270 847.675 4983.440 ;
        RECT 847.845 4983.270 848.135 4983.440 ;
        RECT 848.305 4983.270 848.595 4983.440 ;
        RECT 848.765 4983.270 849.055 4983.440 ;
        RECT 849.225 4983.270 849.515 4983.440 ;
        RECT 849.685 4983.270 849.975 4983.440 ;
        RECT 850.145 4983.270 850.435 4983.440 ;
        RECT 850.605 4983.270 850.895 4983.440 ;
        RECT 851.065 4983.270 851.355 4983.440 ;
        RECT 851.525 4983.270 851.815 4983.440 ;
        RECT 851.985 4983.270 852.275 4983.440 ;
        RECT 852.445 4983.270 852.735 4983.440 ;
        RECT 852.905 4983.270 853.050 4983.440 ;
        RECT 2084.710 4983.335 2087.335 4983.505 ;
        RECT 834.735 4982.105 835.025 4983.270 ;
        RECT 835.585 4982.120 835.915 4983.270 ;
      LAYER li1 ;
        RECT 836.085 4982.250 836.255 4983.100 ;
      LAYER li1 ;
        RECT 836.425 4982.470 836.755 4983.270 ;
      LAYER li1 ;
        RECT 836.925 4982.250 837.095 4983.100 ;
      LAYER li1 ;
        RECT 837.265 4982.470 837.595 4983.270 ;
      LAYER li1 ;
        RECT 837.765 4982.250 837.935 4983.100 ;
      LAYER li1 ;
        RECT 838.105 4982.470 838.435 4983.270 ;
      LAYER li1 ;
        RECT 838.605 4982.250 838.775 4983.100 ;
      LAYER li1 ;
        RECT 839.025 4982.470 839.195 4983.270 ;
        RECT 839.365 4982.250 839.695 4983.100 ;
        RECT 839.865 4982.470 840.035 4983.270 ;
        RECT 840.205 4982.250 840.535 4983.100 ;
      LAYER li1 ;
        RECT 836.085 4982.080 838.775 4982.250 ;
      LAYER li1 ;
        RECT 839.035 4982.080 840.535 4982.250 ;
        RECT 840.715 4982.105 841.005 4983.270 ;
        RECT 841.565 4982.120 841.895 4983.270 ;
      LAYER li1 ;
        RECT 842.065 4982.250 842.235 4983.100 ;
      LAYER li1 ;
        RECT 842.405 4982.470 842.735 4983.270 ;
      LAYER li1 ;
        RECT 842.905 4982.250 843.075 4983.100 ;
      LAYER li1 ;
        RECT 843.245 4982.470 843.575 4983.270 ;
      LAYER li1 ;
        RECT 843.745 4982.250 843.915 4983.100 ;
      LAYER li1 ;
        RECT 844.085 4982.470 844.415 4983.270 ;
      LAYER li1 ;
        RECT 844.585 4982.250 844.755 4983.100 ;
      LAYER li1 ;
        RECT 845.005 4982.470 845.175 4983.270 ;
        RECT 845.345 4982.250 845.675 4983.100 ;
        RECT 845.845 4982.470 846.015 4983.270 ;
        RECT 846.185 4982.250 846.515 4983.100 ;
      LAYER li1 ;
        RECT 842.065 4982.080 844.755 4982.250 ;
      LAYER li1 ;
        RECT 845.015 4982.080 846.515 4982.250 ;
        RECT 846.695 4982.105 846.985 4983.270 ;
        RECT 847.545 4982.120 847.875 4983.270 ;
      LAYER li1 ;
        RECT 848.045 4982.250 848.215 4983.100 ;
      LAYER li1 ;
        RECT 848.385 4982.470 848.715 4983.270 ;
      LAYER li1 ;
        RECT 848.885 4982.250 849.055 4983.100 ;
      LAYER li1 ;
        RECT 849.225 4982.470 849.555 4983.270 ;
      LAYER li1 ;
        RECT 849.725 4982.250 849.895 4983.100 ;
      LAYER li1 ;
        RECT 850.065 4982.470 850.395 4983.270 ;
      LAYER li1 ;
        RECT 850.565 4982.250 850.735 4983.100 ;
      LAYER li1 ;
        RECT 850.985 4982.470 851.155 4983.270 ;
        RECT 851.325 4982.250 851.655 4983.100 ;
        RECT 851.825 4982.470 851.995 4983.270 ;
        RECT 852.165 4982.250 852.495 4983.100 ;
      LAYER li1 ;
        RECT 848.045 4982.080 850.735 4982.250 ;
      LAYER li1 ;
        RECT 850.995 4982.080 852.495 4982.250 ;
        RECT 852.675 4982.105 852.965 4983.270 ;
        RECT 2084.710 4983.165 2084.885 4983.335 ;
      LAYER li1 ;
        RECT 2087.580 4983.165 2087.835 4983.705 ;
      LAYER li1 ;
        RECT 3309.920 4983.320 3310.210 4984.485 ;
        RECT 3310.390 4983.465 3310.720 4984.315 ;
        RECT 3310.890 4983.685 3311.060 4984.485 ;
        RECT 3311.230 4983.465 3311.560 4984.315 ;
        RECT 3311.730 4983.685 3311.900 4984.485 ;
      LAYER li1 ;
        RECT 3312.150 4983.465 3312.320 4984.315 ;
      LAYER li1 ;
        RECT 3312.490 4983.685 3312.820 4984.485 ;
      LAYER li1 ;
        RECT 3312.990 4983.465 3313.160 4984.315 ;
      LAYER li1 ;
        RECT 3313.330 4983.685 3313.660 4984.485 ;
      LAYER li1 ;
        RECT 3313.830 4983.465 3314.000 4984.315 ;
      LAYER li1 ;
        RECT 3314.170 4983.685 3314.500 4984.485 ;
      LAYER li1 ;
        RECT 3314.670 4983.465 3314.840 4984.315 ;
      LAYER li1 ;
        RECT 3310.390 4983.295 3311.890 4983.465 ;
      LAYER li1 ;
        RECT 3312.150 4983.295 3314.840 4983.465 ;
      LAYER li1 ;
        RECT 3315.010 4983.335 3315.340 4984.485 ;
        RECT 3315.900 4983.320 3316.190 4984.485 ;
        RECT 3316.370 4983.465 3316.700 4984.315 ;
        RECT 3316.870 4983.685 3317.040 4984.485 ;
        RECT 3317.210 4983.465 3317.540 4984.315 ;
        RECT 3317.710 4983.685 3317.880 4984.485 ;
      LAYER li1 ;
        RECT 3318.130 4983.465 3318.300 4984.315 ;
      LAYER li1 ;
        RECT 3318.470 4983.685 3318.800 4984.485 ;
      LAYER li1 ;
        RECT 3318.970 4983.465 3319.140 4984.315 ;
      LAYER li1 ;
        RECT 3319.310 4983.685 3319.640 4984.485 ;
      LAYER li1 ;
        RECT 3319.810 4983.465 3319.980 4984.315 ;
      LAYER li1 ;
        RECT 3320.150 4983.685 3320.480 4984.485 ;
      LAYER li1 ;
        RECT 3320.650 4983.465 3320.820 4984.315 ;
      LAYER li1 ;
        RECT 3316.370 4983.295 3317.870 4983.465 ;
      LAYER li1 ;
        RECT 3318.130 4983.295 3320.820 4983.465 ;
      LAYER li1 ;
        RECT 3320.990 4983.335 3321.320 4984.485 ;
        RECT 3321.880 4983.320 3322.170 4984.485 ;
        RECT 3322.350 4983.465 3322.680 4984.315 ;
        RECT 3322.850 4983.685 3323.020 4984.485 ;
        RECT 3323.190 4983.465 3323.520 4984.315 ;
        RECT 3323.690 4983.685 3323.860 4984.485 ;
      LAYER li1 ;
        RECT 3324.110 4983.465 3324.280 4984.315 ;
      LAYER li1 ;
        RECT 3324.450 4983.685 3324.780 4984.485 ;
      LAYER li1 ;
        RECT 3324.950 4983.465 3325.120 4984.315 ;
      LAYER li1 ;
        RECT 3325.290 4983.685 3325.620 4984.485 ;
      LAYER li1 ;
        RECT 3325.790 4983.465 3325.960 4984.315 ;
      LAYER li1 ;
        RECT 3326.130 4983.685 3326.460 4984.485 ;
      LAYER li1 ;
        RECT 3326.630 4983.465 3326.800 4984.315 ;
      LAYER li1 ;
        RECT 3322.350 4983.295 3323.850 4983.465 ;
      LAYER li1 ;
        RECT 3324.110 4983.295 3326.800 4983.465 ;
      LAYER li1 ;
        RECT 3326.970 4983.335 3327.300 4984.485 ;
        RECT 3327.860 4983.320 3328.150 4984.485 ;
        RECT 3328.330 4983.465 3328.660 4984.315 ;
        RECT 3328.830 4983.685 3329.000 4984.485 ;
        RECT 3329.170 4983.465 3329.500 4984.315 ;
        RECT 3329.670 4983.685 3329.840 4984.485 ;
      LAYER li1 ;
        RECT 3330.090 4983.465 3330.260 4984.315 ;
      LAYER li1 ;
        RECT 3330.430 4983.685 3330.760 4984.485 ;
      LAYER li1 ;
        RECT 3330.930 4983.465 3331.100 4984.315 ;
      LAYER li1 ;
        RECT 3331.270 4983.685 3331.600 4984.485 ;
      LAYER li1 ;
        RECT 3331.770 4983.465 3331.940 4984.315 ;
      LAYER li1 ;
        RECT 3332.110 4983.685 3332.440 4984.485 ;
      LAYER li1 ;
        RECT 3332.610 4983.465 3332.780 4984.315 ;
      LAYER li1 ;
        RECT 3328.330 4983.295 3329.830 4983.465 ;
      LAYER li1 ;
        RECT 3330.090 4983.295 3332.780 4983.465 ;
      LAYER li1 ;
        RECT 3332.950 4983.335 3333.280 4984.485 ;
        RECT 3333.840 4983.320 3334.130 4984.485 ;
        RECT 2082.915 4982.345 2083.205 4983.070 ;
        RECT 2083.465 4982.995 2084.885 4983.165 ;
      LAYER li1 ;
        RECT 2085.145 4982.995 2087.835 4983.165 ;
      LAYER li1 ;
        RECT 2083.465 4982.515 2083.635 4982.995 ;
        RECT 2083.805 4982.345 2084.135 4982.825 ;
        RECT 2084.305 4982.520 2084.475 4982.995 ;
        RECT 2084.645 4982.345 2084.975 4982.825 ;
      LAYER li1 ;
        RECT 2085.145 4982.515 2085.315 4982.995 ;
      LAYER li1 ;
        RECT 2085.485 4982.345 2085.815 4982.825 ;
      LAYER li1 ;
        RECT 2085.985 4982.515 2086.155 4982.995 ;
      LAYER li1 ;
        RECT 2086.325 4982.345 2086.655 4982.825 ;
      LAYER li1 ;
        RECT 2086.825 4982.515 2086.995 4982.995 ;
      LAYER li1 ;
        RECT 2087.165 4982.345 2087.495 4982.825 ;
      LAYER li1 ;
        RECT 2087.665 4982.515 2087.835 4982.995 ;
      LAYER li1 ;
        RECT 2088.005 4982.345 2088.335 4983.145 ;
        RECT 2088.895 4982.345 2089.185 4983.070 ;
      LAYER li1 ;
        RECT 3309.945 4982.925 3311.535 4983.125 ;
      LAYER li1 ;
        RECT 3311.715 4983.095 3311.890 4983.295 ;
        RECT 3311.715 4982.925 3314.340 4983.095 ;
        RECT 3311.715 4982.755 3311.890 4982.925 ;
      LAYER li1 ;
        RECT 3314.585 4982.755 3314.840 4983.295 ;
      LAYER li1 ;
        RECT 3317.695 4983.095 3317.870 4983.295 ;
        RECT 3317.695 4982.925 3320.320 4983.095 ;
        RECT 3317.695 4982.755 3317.870 4982.925 ;
      LAYER li1 ;
        RECT 3320.565 4982.755 3320.820 4983.295 ;
      LAYER li1 ;
        RECT 3323.675 4983.095 3323.850 4983.295 ;
        RECT 3323.675 4982.925 3326.300 4983.095 ;
        RECT 3323.675 4982.755 3323.850 4982.925 ;
      LAYER li1 ;
        RECT 3326.545 4982.755 3326.800 4983.295 ;
      LAYER li1 ;
        RECT 3329.655 4983.095 3329.830 4983.295 ;
        RECT 3329.655 4982.925 3332.280 4983.095 ;
        RECT 3329.655 4982.755 3329.830 4982.925 ;
      LAYER li1 ;
        RECT 3332.525 4982.755 3332.780 4983.295 ;
      LAYER li1 ;
        RECT 2082.830 4982.175 2082.975 4982.345 ;
        RECT 2083.145 4982.175 2083.435 4982.345 ;
        RECT 2083.605 4982.175 2083.895 4982.345 ;
        RECT 2084.065 4982.175 2084.355 4982.345 ;
        RECT 2084.525 4982.175 2084.815 4982.345 ;
        RECT 2084.985 4982.175 2085.275 4982.345 ;
        RECT 2085.445 4982.175 2085.735 4982.345 ;
        RECT 2085.905 4982.175 2086.195 4982.345 ;
        RECT 2086.365 4982.175 2086.655 4982.345 ;
        RECT 2086.825 4982.175 2087.115 4982.345 ;
        RECT 2087.285 4982.175 2087.575 4982.345 ;
        RECT 2087.745 4982.175 2088.035 4982.345 ;
        RECT 2088.205 4982.175 2088.495 4982.345 ;
        RECT 2088.665 4982.175 2088.955 4982.345 ;
        RECT 2089.125 4982.175 2089.270 4982.345 ;
      LAYER li1 ;
        RECT 836.085 4981.540 836.340 4982.080 ;
      LAYER li1 ;
        RECT 839.035 4981.880 839.210 4982.080 ;
        RECT 836.585 4981.710 839.210 4981.880 ;
        RECT 839.035 4981.540 839.210 4981.710 ;
      LAYER li1 ;
        RECT 842.065 4981.540 842.320 4982.080 ;
      LAYER li1 ;
        RECT 845.015 4981.880 845.190 4982.080 ;
        RECT 842.565 4981.710 845.190 4981.880 ;
        RECT 845.015 4981.540 845.190 4981.710 ;
      LAYER li1 ;
        RECT 848.045 4981.540 848.300 4982.080 ;
      LAYER li1 ;
        RECT 850.995 4981.880 851.170 4982.080 ;
        RECT 848.545 4981.710 851.170 4981.880 ;
        RECT 850.995 4981.540 851.170 4981.710 ;
        RECT 834.735 4980.720 835.025 4981.445 ;
        RECT 835.585 4980.720 835.915 4981.520 ;
      LAYER li1 ;
        RECT 836.085 4981.370 838.775 4981.540 ;
      LAYER li1 ;
        RECT 839.035 4981.370 840.455 4981.540 ;
      LAYER li1 ;
        RECT 836.085 4980.890 836.255 4981.370 ;
      LAYER li1 ;
        RECT 836.425 4980.720 836.755 4981.200 ;
      LAYER li1 ;
        RECT 836.925 4980.890 837.095 4981.370 ;
      LAYER li1 ;
        RECT 837.265 4980.720 837.595 4981.200 ;
      LAYER li1 ;
        RECT 837.765 4980.890 837.935 4981.370 ;
      LAYER li1 ;
        RECT 838.105 4980.720 838.435 4981.200 ;
      LAYER li1 ;
        RECT 838.605 4980.890 838.775 4981.370 ;
      LAYER li1 ;
        RECT 838.945 4980.720 839.275 4981.200 ;
        RECT 839.445 4980.895 839.615 4981.370 ;
        RECT 839.785 4980.720 840.115 4981.200 ;
        RECT 840.285 4980.890 840.455 4981.370 ;
        RECT 840.715 4980.720 841.005 4981.445 ;
        RECT 841.565 4980.720 841.895 4981.520 ;
      LAYER li1 ;
        RECT 842.065 4981.370 844.755 4981.540 ;
      LAYER li1 ;
        RECT 845.015 4981.370 846.435 4981.540 ;
      LAYER li1 ;
        RECT 842.065 4980.890 842.235 4981.370 ;
      LAYER li1 ;
        RECT 842.405 4980.720 842.735 4981.200 ;
      LAYER li1 ;
        RECT 842.905 4980.890 843.075 4981.370 ;
      LAYER li1 ;
        RECT 843.245 4980.720 843.575 4981.200 ;
      LAYER li1 ;
        RECT 843.745 4980.890 843.915 4981.370 ;
      LAYER li1 ;
        RECT 844.085 4980.720 844.415 4981.200 ;
      LAYER li1 ;
        RECT 844.585 4980.890 844.755 4981.370 ;
      LAYER li1 ;
        RECT 844.925 4980.720 845.255 4981.200 ;
        RECT 845.425 4980.895 845.595 4981.370 ;
        RECT 845.765 4980.720 846.095 4981.200 ;
        RECT 846.265 4980.890 846.435 4981.370 ;
        RECT 846.695 4980.720 846.985 4981.445 ;
        RECT 847.545 4980.720 847.875 4981.520 ;
      LAYER li1 ;
        RECT 848.045 4981.370 850.735 4981.540 ;
      LAYER li1 ;
        RECT 850.995 4981.370 852.415 4981.540 ;
        RECT 2082.915 4981.450 2083.205 4982.175 ;
      LAYER li1 ;
        RECT 2083.380 4981.630 2088.725 4982.175 ;
        RECT 848.045 4980.890 848.215 4981.370 ;
      LAYER li1 ;
        RECT 848.385 4980.720 848.715 4981.200 ;
      LAYER li1 ;
        RECT 848.885 4980.890 849.055 4981.370 ;
      LAYER li1 ;
        RECT 849.225 4980.720 849.555 4981.200 ;
      LAYER li1 ;
        RECT 849.725 4980.890 849.895 4981.370 ;
      LAYER li1 ;
        RECT 850.065 4980.720 850.395 4981.200 ;
      LAYER li1 ;
        RECT 850.565 4980.890 850.735 4981.370 ;
      LAYER li1 ;
        RECT 850.905 4980.720 851.235 4981.200 ;
        RECT 851.405 4980.895 851.575 4981.370 ;
        RECT 851.745 4980.720 852.075 4981.200 ;
        RECT 852.245 4980.890 852.415 4981.370 ;
        RECT 852.675 4980.720 852.965 4981.445 ;
      LAYER li1 ;
        RECT 2086.800 4980.800 2087.140 4981.630 ;
      LAYER li1 ;
        RECT 2088.895 4981.450 2089.185 4982.175 ;
        RECT 3309.920 4981.935 3310.210 4982.660 ;
        RECT 3310.470 4982.585 3311.890 4982.755 ;
      LAYER li1 ;
        RECT 3312.150 4982.585 3314.840 4982.755 ;
      LAYER li1 ;
        RECT 3310.470 4982.105 3310.640 4982.585 ;
        RECT 3310.810 4981.935 3311.140 4982.415 ;
        RECT 3311.310 4982.110 3311.480 4982.585 ;
        RECT 3311.650 4981.935 3311.980 4982.415 ;
      LAYER li1 ;
        RECT 3312.150 4982.105 3312.320 4982.585 ;
      LAYER li1 ;
        RECT 3312.490 4981.935 3312.820 4982.415 ;
      LAYER li1 ;
        RECT 3312.990 4982.105 3313.160 4982.585 ;
      LAYER li1 ;
        RECT 3313.330 4981.935 3313.660 4982.415 ;
      LAYER li1 ;
        RECT 3313.830 4982.105 3314.000 4982.585 ;
      LAYER li1 ;
        RECT 3314.170 4981.935 3314.500 4982.415 ;
      LAYER li1 ;
        RECT 3314.670 4982.105 3314.840 4982.585 ;
      LAYER li1 ;
        RECT 3315.010 4981.935 3315.340 4982.735 ;
        RECT 3315.900 4981.935 3316.190 4982.660 ;
        RECT 3316.450 4982.585 3317.870 4982.755 ;
      LAYER li1 ;
        RECT 3318.130 4982.585 3320.820 4982.755 ;
      LAYER li1 ;
        RECT 3316.450 4982.105 3316.620 4982.585 ;
        RECT 3316.790 4981.935 3317.120 4982.415 ;
        RECT 3317.290 4982.110 3317.460 4982.585 ;
        RECT 3317.630 4981.935 3317.960 4982.415 ;
      LAYER li1 ;
        RECT 3318.130 4982.105 3318.300 4982.585 ;
      LAYER li1 ;
        RECT 3318.470 4981.935 3318.800 4982.415 ;
      LAYER li1 ;
        RECT 3318.970 4982.105 3319.140 4982.585 ;
      LAYER li1 ;
        RECT 3319.310 4981.935 3319.640 4982.415 ;
      LAYER li1 ;
        RECT 3319.810 4982.105 3319.980 4982.585 ;
      LAYER li1 ;
        RECT 3320.150 4981.935 3320.480 4982.415 ;
      LAYER li1 ;
        RECT 3320.650 4982.105 3320.820 4982.585 ;
      LAYER li1 ;
        RECT 3320.990 4981.935 3321.320 4982.735 ;
        RECT 3321.880 4981.935 3322.170 4982.660 ;
        RECT 3322.430 4982.585 3323.850 4982.755 ;
      LAYER li1 ;
        RECT 3324.110 4982.585 3326.800 4982.755 ;
      LAYER li1 ;
        RECT 3322.430 4982.105 3322.600 4982.585 ;
        RECT 3322.770 4981.935 3323.100 4982.415 ;
        RECT 3323.270 4982.110 3323.440 4982.585 ;
        RECT 3323.610 4981.935 3323.940 4982.415 ;
      LAYER li1 ;
        RECT 3324.110 4982.105 3324.280 4982.585 ;
      LAYER li1 ;
        RECT 3324.450 4981.935 3324.780 4982.415 ;
      LAYER li1 ;
        RECT 3324.950 4982.105 3325.120 4982.585 ;
      LAYER li1 ;
        RECT 3325.290 4981.935 3325.620 4982.415 ;
      LAYER li1 ;
        RECT 3325.790 4982.105 3325.960 4982.585 ;
      LAYER li1 ;
        RECT 3326.130 4981.935 3326.460 4982.415 ;
      LAYER li1 ;
        RECT 3326.630 4982.105 3326.800 4982.585 ;
      LAYER li1 ;
        RECT 3326.970 4981.935 3327.300 4982.735 ;
        RECT 3327.860 4981.935 3328.150 4982.660 ;
        RECT 3328.410 4982.585 3329.830 4982.755 ;
      LAYER li1 ;
        RECT 3330.090 4982.585 3332.780 4982.755 ;
      LAYER li1 ;
        RECT 3328.410 4982.105 3328.580 4982.585 ;
        RECT 3328.750 4981.935 3329.080 4982.415 ;
        RECT 3329.250 4982.110 3329.420 4982.585 ;
        RECT 3329.590 4981.935 3329.920 4982.415 ;
      LAYER li1 ;
        RECT 3330.090 4982.105 3330.260 4982.585 ;
      LAYER li1 ;
        RECT 3330.430 4981.935 3330.760 4982.415 ;
      LAYER li1 ;
        RECT 3330.930 4982.105 3331.100 4982.585 ;
      LAYER li1 ;
        RECT 3331.270 4981.935 3331.600 4982.415 ;
      LAYER li1 ;
        RECT 3331.770 4982.105 3331.940 4982.585 ;
      LAYER li1 ;
        RECT 3332.110 4981.935 3332.440 4982.415 ;
      LAYER li1 ;
        RECT 3332.610 4982.105 3332.780 4982.585 ;
      LAYER li1 ;
        RECT 3332.950 4981.935 3333.280 4982.735 ;
        RECT 3333.840 4981.935 3334.130 4982.660 ;
        RECT 3309.835 4981.765 3309.980 4981.935 ;
        RECT 3310.150 4981.765 3310.295 4981.935 ;
        RECT 3315.815 4981.765 3315.960 4981.935 ;
        RECT 3316.130 4981.765 3316.420 4981.935 ;
        RECT 3316.590 4981.765 3316.880 4981.935 ;
        RECT 3317.050 4981.765 3317.340 4981.935 ;
        RECT 3317.510 4981.765 3317.800 4981.935 ;
        RECT 3317.970 4981.765 3318.260 4981.935 ;
        RECT 3318.430 4981.765 3318.720 4981.935 ;
        RECT 3318.890 4981.765 3319.180 4981.935 ;
        RECT 3319.350 4981.765 3319.640 4981.935 ;
        RECT 3319.810 4981.765 3320.100 4981.935 ;
        RECT 3320.270 4981.765 3320.560 4981.935 ;
        RECT 3320.730 4981.765 3321.020 4981.935 ;
        RECT 3321.190 4981.765 3321.480 4981.935 ;
        RECT 3321.650 4981.765 3321.940 4981.935 ;
        RECT 3322.110 4981.765 3322.400 4981.935 ;
        RECT 3322.570 4981.765 3322.860 4981.935 ;
        RECT 3323.030 4981.765 3323.320 4981.935 ;
        RECT 3323.490 4981.765 3323.780 4981.935 ;
        RECT 3323.950 4981.765 3324.240 4981.935 ;
        RECT 3324.410 4981.765 3324.700 4981.935 ;
        RECT 3324.870 4981.765 3325.160 4981.935 ;
        RECT 3325.330 4981.765 3325.620 4981.935 ;
        RECT 3325.790 4981.765 3326.080 4981.935 ;
        RECT 3326.250 4981.765 3326.540 4981.935 ;
        RECT 3326.710 4981.765 3327.000 4981.935 ;
        RECT 3327.170 4981.765 3327.460 4981.935 ;
        RECT 3327.630 4981.765 3327.920 4981.935 ;
        RECT 3328.090 4981.765 3328.380 4981.935 ;
        RECT 3328.550 4981.765 3328.840 4981.935 ;
        RECT 3329.010 4981.765 3329.300 4981.935 ;
        RECT 3329.470 4981.765 3329.760 4981.935 ;
        RECT 3329.930 4981.765 3330.220 4981.935 ;
        RECT 3330.390 4981.765 3330.680 4981.935 ;
        RECT 3330.850 4981.765 3331.140 4981.935 ;
        RECT 3331.310 4981.765 3331.600 4981.935 ;
        RECT 3331.770 4981.765 3332.060 4981.935 ;
        RECT 3332.230 4981.765 3332.520 4981.935 ;
        RECT 3332.690 4981.765 3332.980 4981.935 ;
        RECT 3333.150 4981.765 3333.440 4981.935 ;
        RECT 3333.610 4981.765 3333.900 4981.935 ;
        RECT 3334.070 4981.765 3334.215 4981.935 ;
        RECT 3309.920 4981.040 3310.210 4981.765 ;
        RECT 3315.900 4981.040 3316.190 4981.765 ;
      LAYER li1 ;
        RECT 3316.365 4981.220 3321.710 4981.765 ;
      LAYER li1 ;
        RECT 834.650 4980.550 834.795 4980.720 ;
        RECT 834.965 4980.550 835.255 4980.720 ;
        RECT 835.425 4980.550 835.715 4980.720 ;
        RECT 835.885 4980.550 836.175 4980.720 ;
        RECT 836.345 4980.550 836.635 4980.720 ;
        RECT 836.805 4980.550 837.095 4980.720 ;
        RECT 837.265 4980.550 837.555 4980.720 ;
        RECT 837.725 4980.550 838.015 4980.720 ;
        RECT 838.185 4980.550 838.475 4980.720 ;
        RECT 838.645 4980.550 838.935 4980.720 ;
        RECT 839.105 4980.550 839.395 4980.720 ;
        RECT 839.565 4980.550 839.855 4980.720 ;
        RECT 840.025 4980.550 840.315 4980.720 ;
        RECT 840.485 4980.550 840.775 4980.720 ;
        RECT 840.945 4980.550 841.235 4980.720 ;
        RECT 841.405 4980.550 841.695 4980.720 ;
        RECT 841.865 4980.550 842.155 4980.720 ;
        RECT 842.325 4980.550 842.615 4980.720 ;
        RECT 842.785 4980.550 843.075 4980.720 ;
        RECT 843.245 4980.550 843.535 4980.720 ;
        RECT 843.705 4980.550 843.995 4980.720 ;
        RECT 844.165 4980.550 844.455 4980.720 ;
        RECT 844.625 4980.550 844.915 4980.720 ;
        RECT 845.085 4980.550 845.375 4980.720 ;
        RECT 845.545 4980.550 845.835 4980.720 ;
        RECT 846.005 4980.550 846.295 4980.720 ;
        RECT 846.465 4980.550 846.755 4980.720 ;
        RECT 846.925 4980.550 847.215 4980.720 ;
        RECT 847.385 4980.550 847.675 4980.720 ;
        RECT 847.845 4980.550 848.135 4980.720 ;
        RECT 848.305 4980.550 848.595 4980.720 ;
        RECT 848.765 4980.550 849.055 4980.720 ;
        RECT 849.225 4980.550 849.515 4980.720 ;
        RECT 849.685 4980.550 849.975 4980.720 ;
        RECT 850.145 4980.550 850.435 4980.720 ;
        RECT 850.605 4980.550 850.895 4980.720 ;
        RECT 851.065 4980.550 851.355 4980.720 ;
        RECT 851.525 4980.550 851.815 4980.720 ;
        RECT 851.985 4980.550 852.275 4980.720 ;
        RECT 852.445 4980.550 852.735 4980.720 ;
        RECT 852.905 4980.550 853.050 4980.720 ;
        RECT 834.735 4979.825 835.025 4980.550 ;
      LAYER li1 ;
        RECT 835.200 4980.005 840.545 4980.550 ;
        RECT 838.620 4979.175 838.960 4980.005 ;
      LAYER li1 ;
        RECT 840.715 4979.825 841.005 4980.550 ;
      LAYER li1 ;
        RECT 841.180 4980.005 846.525 4980.550 ;
        RECT 844.600 4979.175 844.940 4980.005 ;
      LAYER li1 ;
        RECT 846.695 4979.825 846.985 4980.550 ;
      LAYER li1 ;
        RECT 847.160 4980.005 852.505 4980.550 ;
        RECT 850.580 4979.175 850.920 4980.005 ;
      LAYER li1 ;
        RECT 852.675 4979.825 852.965 4980.550 ;
        RECT 2082.915 4979.625 2083.205 4980.790 ;
        RECT 2088.895 4979.625 2089.185 4980.790 ;
      LAYER li1 ;
        RECT 3319.785 4980.390 3320.125 4981.220 ;
      LAYER li1 ;
        RECT 3321.880 4981.040 3322.170 4981.765 ;
      LAYER li1 ;
        RECT 3322.345 4981.220 3327.690 4981.765 ;
        RECT 3325.765 4980.390 3326.105 4981.220 ;
      LAYER li1 ;
        RECT 3327.860 4981.040 3328.150 4981.765 ;
      LAYER li1 ;
        RECT 3328.325 4981.220 3333.670 4981.765 ;
        RECT 3331.745 4980.390 3332.085 4981.220 ;
      LAYER li1 ;
        RECT 3333.840 4981.040 3334.130 4981.765 ;
        RECT 2082.830 4979.455 2082.975 4979.625 ;
        RECT 2083.145 4979.455 2083.290 4979.625 ;
        RECT 2088.810 4979.455 2088.955 4979.625 ;
        RECT 2089.125 4979.455 2089.270 4979.625 ;
        RECT 3309.920 4979.215 3310.210 4980.380 ;
        RECT 3315.900 4979.215 3316.190 4980.380 ;
        RECT 3321.880 4979.215 3322.170 4980.380 ;
        RECT 3327.860 4979.215 3328.150 4980.380 ;
        RECT 3333.840 4979.215 3334.130 4980.380 ;
        RECT 834.735 4978.000 835.025 4979.165 ;
        RECT 840.715 4978.000 841.005 4979.165 ;
        RECT 846.695 4978.000 846.985 4979.165 ;
        RECT 852.675 4978.000 852.965 4979.165 ;
        RECT 3309.835 4979.045 3309.980 4979.215 ;
        RECT 3310.150 4979.045 3310.295 4979.215 ;
        RECT 3315.815 4979.045 3315.960 4979.215 ;
        RECT 3316.130 4979.045 3316.275 4979.215 ;
        RECT 3321.795 4979.045 3321.940 4979.215 ;
        RECT 3322.110 4979.045 3322.255 4979.215 ;
        RECT 3327.775 4979.045 3327.920 4979.215 ;
        RECT 3328.090 4979.045 3328.235 4979.215 ;
        RECT 3333.755 4979.045 3333.900 4979.215 ;
        RECT 3334.070 4979.045 3334.215 4979.215 ;
        RECT 834.650 4977.830 834.795 4978.000 ;
        RECT 834.965 4977.830 835.110 4978.000 ;
        RECT 840.630 4977.830 840.775 4978.000 ;
        RECT 840.945 4977.830 841.090 4978.000 ;
        RECT 846.610 4977.830 846.755 4978.000 ;
        RECT 846.925 4977.830 847.070 4978.000 ;
        RECT 852.590 4977.830 852.735 4978.000 ;
        RECT 852.905 4977.830 853.050 4978.000 ;
        RECT 201.760 4457.115 201.930 4457.200 ;
        RECT 204.480 4457.115 204.650 4457.200 ;
        RECT 207.200 4457.115 207.370 4457.200 ;
        RECT 209.920 4457.115 210.090 4457.200 ;
        RECT 201.760 4457.055 202.655 4457.115 ;
        RECT 201.930 4456.885 202.655 4457.055 ;
        RECT 201.760 4456.825 202.655 4456.885 ;
        RECT 203.315 4457.055 205.815 4457.115 ;
        RECT 203.315 4456.885 204.480 4457.055 ;
        RECT 204.650 4456.885 205.815 4457.055 ;
        RECT 203.315 4456.825 205.815 4456.885 ;
        RECT 201.760 4456.595 201.930 4456.825 ;
        RECT 204.480 4456.595 204.650 4456.825 ;
        RECT 201.760 4456.265 201.930 4456.425 ;
        RECT 204.480 4456.265 204.650 4456.425 ;
        RECT 204.820 4456.315 205.840 4456.645 ;
        RECT 201.760 4456.135 202.730 4456.265 ;
        RECT 201.930 4455.965 202.730 4456.135 ;
        RECT 201.760 4455.935 202.730 4455.965 ;
        RECT 203.330 4456.145 204.650 4456.265 ;
        RECT 203.330 4456.135 205.450 4456.145 ;
        RECT 203.330 4455.965 204.480 4456.135 ;
        RECT 204.650 4455.975 205.450 4456.135 ;
        RECT 203.330 4455.935 204.650 4455.965 ;
        RECT 201.760 4455.675 201.930 4455.935 ;
      LAYER li1 ;
        RECT 202.100 4455.595 204.310 4455.765 ;
      LAYER li1 ;
        RECT 204.480 4455.675 204.650 4455.935 ;
        RECT 205.670 4455.805 205.840 4456.315 ;
      LAYER li1 ;
        RECT 202.580 4455.510 203.460 4455.595 ;
      LAYER li1 ;
        RECT 201.760 4455.425 201.930 4455.505 ;
        RECT 201.760 4455.215 202.410 4455.425 ;
        RECT 201.930 4455.095 202.410 4455.215 ;
        RECT 201.760 4454.755 201.930 4455.045 ;
      LAYER li1 ;
        RECT 202.580 4454.925 202.750 4455.510 ;
        RECT 202.100 4454.755 202.750 4454.925 ;
      LAYER li1 ;
        RECT 201.760 4454.295 202.410 4454.585 ;
        RECT 201.930 4454.255 202.410 4454.295 ;
        RECT 201.760 4453.835 201.930 4454.125 ;
      LAYER li1 ;
        RECT 202.580 4454.085 202.750 4454.755 ;
        RECT 202.100 4453.915 202.750 4454.085 ;
      LAYER li1 ;
        RECT 201.930 4453.665 202.410 4453.745 ;
        RECT 201.760 4453.415 202.410 4453.665 ;
        RECT 201.760 4453.375 201.930 4453.415 ;
      LAYER li1 ;
        RECT 202.580 4453.245 202.750 4453.915 ;
      LAYER li1 ;
        RECT 201.760 4452.915 201.930 4453.205 ;
      LAYER li1 ;
        RECT 202.100 4453.075 202.750 4453.245 ;
      LAYER li1 ;
        RECT 201.930 4452.745 202.410 4452.905 ;
        RECT 202.920 4452.815 203.090 4455.265 ;
      LAYER li1 ;
        RECT 203.290 4454.925 203.460 4455.510 ;
      LAYER li1 ;
        RECT 204.480 4455.425 204.650 4455.505 ;
        RECT 204.820 4455.475 205.840 4455.805 ;
      LAYER li1 ;
        RECT 206.010 4455.500 206.210 4457.090 ;
      LAYER li1 ;
        RECT 206.475 4457.055 208.095 4457.115 ;
        RECT 206.475 4456.885 207.200 4457.055 ;
        RECT 207.370 4456.885 208.095 4457.055 ;
        RECT 206.475 4456.825 208.095 4456.885 ;
        RECT 208.755 4457.055 210.090 4457.115 ;
        RECT 208.755 4456.885 209.920 4457.055 ;
        RECT 208.755 4456.825 210.090 4456.885 ;
        RECT 207.200 4456.595 207.370 4456.825 ;
        RECT 209.920 4456.740 210.090 4456.825 ;
        RECT 206.380 4456.395 207.030 4456.565 ;
        RECT 206.380 4455.725 206.550 4456.395 ;
        RECT 207.200 4456.225 207.370 4456.425 ;
        RECT 206.720 4456.135 207.370 4456.225 ;
        RECT 206.720 4455.965 207.200 4456.135 ;
        RECT 206.720 4455.895 207.370 4455.965 ;
        RECT 206.380 4455.555 207.025 4455.725 ;
        RECT 207.200 4455.675 207.370 4455.895 ;
        RECT 203.680 4455.305 204.650 4455.425 ;
        RECT 205.670 4455.320 205.840 4455.475 ;
        RECT 206.380 4455.320 206.550 4455.555 ;
        RECT 207.200 4455.385 207.370 4455.505 ;
        RECT 203.680 4455.215 205.450 4455.305 ;
        RECT 203.680 4455.095 204.480 4455.215 ;
        RECT 204.650 4455.135 205.450 4455.215 ;
        RECT 205.670 4455.145 206.550 4455.320 ;
        RECT 206.720 4455.215 207.370 4455.385 ;
      LAYER li1 ;
        RECT 203.290 4454.755 204.310 4454.925 ;
      LAYER li1 ;
        RECT 204.480 4454.755 204.650 4455.045 ;
      LAYER li1 ;
        RECT 203.290 4454.085 203.460 4454.755 ;
        RECT 204.820 4454.715 205.840 4454.885 ;
      LAYER li1 ;
        RECT 203.680 4454.545 204.650 4454.585 ;
        RECT 203.680 4454.295 205.450 4454.545 ;
        RECT 203.680 4454.255 204.480 4454.295 ;
        RECT 204.650 4454.215 205.450 4454.295 ;
      LAYER li1 ;
        RECT 203.290 4453.915 204.310 4454.085 ;
        RECT 203.290 4453.245 203.460 4453.915 ;
      LAYER li1 ;
        RECT 204.480 4453.835 204.650 4454.125 ;
      LAYER li1 ;
        RECT 205.670 4454.045 205.840 4454.715 ;
        RECT 204.820 4453.875 205.840 4454.045 ;
      LAYER li1 ;
        RECT 203.680 4453.665 204.480 4453.745 ;
        RECT 204.650 4453.665 205.450 4453.705 ;
        RECT 203.680 4453.415 205.450 4453.665 ;
        RECT 204.480 4453.375 205.450 4453.415 ;
      LAYER li1 ;
        RECT 203.290 4453.075 204.310 4453.245 ;
        RECT 205.670 4453.205 205.840 4453.875 ;
      LAYER li1 ;
        RECT 204.480 4452.915 204.650 4453.205 ;
      LAYER li1 ;
        RECT 204.820 4453.035 205.840 4453.205 ;
      LAYER li1 ;
        RECT 201.760 4452.575 202.410 4452.745 ;
        RECT 202.580 4452.640 203.460 4452.815 ;
        RECT 203.680 4452.745 204.480 4452.825 ;
        RECT 204.650 4452.745 205.450 4452.865 ;
        RECT 203.680 4452.655 205.450 4452.745 ;
        RECT 201.760 4452.455 201.930 4452.575 ;
        RECT 202.580 4452.405 202.750 4452.640 ;
        RECT 203.290 4452.485 203.460 4452.640 ;
        RECT 204.480 4452.535 205.450 4452.655 ;
        RECT 201.760 4452.065 201.930 4452.285 ;
        RECT 202.105 4452.235 202.750 4452.405 ;
        RECT 201.760 4451.995 202.410 4452.065 ;
        RECT 201.930 4451.825 202.410 4451.995 ;
        RECT 201.760 4451.735 202.410 4451.825 ;
        RECT 201.760 4451.535 201.930 4451.735 ;
        RECT 202.580 4451.565 202.750 4452.235 ;
        RECT 202.100 4451.395 202.750 4451.565 ;
        RECT 201.760 4451.135 201.930 4451.365 ;
      LAYER li1 ;
        RECT 202.920 4451.360 203.120 4452.460 ;
      LAYER li1 ;
        RECT 203.290 4452.155 204.310 4452.485 ;
        RECT 204.480 4452.455 204.650 4452.535 ;
      LAYER li1 ;
        RECT 205.670 4452.450 205.840 4453.035 ;
      LAYER li1 ;
        RECT 206.040 4452.695 206.210 4455.145 ;
        RECT 206.720 4455.055 207.200 4455.215 ;
      LAYER li1 ;
        RECT 207.370 4455.070 207.915 4456.655 ;
        RECT 206.380 4454.715 207.030 4454.885 ;
      LAYER li1 ;
        RECT 207.200 4454.755 207.370 4455.045 ;
      LAYER li1 ;
        RECT 207.370 4454.730 208.745 4455.070 ;
        RECT 206.380 4454.045 206.550 4454.715 ;
      LAYER li1 ;
        RECT 207.200 4454.545 207.370 4454.585 ;
        RECT 206.720 4454.295 207.370 4454.545 ;
        RECT 206.720 4454.215 207.200 4454.295 ;
      LAYER li1 ;
        RECT 206.380 4453.875 207.030 4454.045 ;
        RECT 206.380 4453.205 206.550 4453.875 ;
      LAYER li1 ;
        RECT 207.200 4453.835 207.370 4454.125 ;
        RECT 206.720 4453.665 207.200 4453.705 ;
        RECT 206.720 4453.375 207.370 4453.665 ;
      LAYER li1 ;
        RECT 206.380 4453.035 207.030 4453.205 ;
        RECT 206.380 4452.450 206.550 4453.035 ;
      LAYER li1 ;
        RECT 207.200 4452.915 207.370 4453.205 ;
        RECT 206.720 4452.745 207.200 4452.865 ;
        RECT 206.720 4452.535 207.370 4452.745 ;
        RECT 207.200 4452.455 207.370 4452.535 ;
      LAYER li1 ;
        RECT 205.670 4452.365 206.550 4452.450 ;
      LAYER li1 ;
        RECT 203.290 4451.645 203.460 4452.155 ;
        RECT 204.480 4452.025 204.650 4452.285 ;
      LAYER li1 ;
        RECT 204.820 4452.195 207.030 4452.365 ;
      LAYER li1 ;
        RECT 207.200 4452.025 207.370 4452.285 ;
        RECT 204.480 4451.995 205.800 4452.025 ;
        RECT 203.680 4451.825 204.480 4451.985 ;
        RECT 204.650 4451.825 205.800 4451.995 ;
        RECT 203.680 4451.815 205.800 4451.825 ;
        RECT 204.480 4451.695 205.800 4451.815 ;
        RECT 206.400 4451.995 207.370 4452.025 ;
        RECT 206.400 4451.825 207.200 4451.995 ;
        RECT 206.400 4451.695 207.370 4451.825 ;
        RECT 203.290 4451.315 204.310 4451.645 ;
        RECT 204.480 4451.535 204.650 4451.695 ;
        RECT 207.200 4451.535 207.370 4451.695 ;
        RECT 204.480 4451.135 204.650 4451.365 ;
        RECT 207.200 4451.135 207.370 4451.365 ;
      LAYER li1 ;
        RECT 207.370 4451.310 207.915 4454.730 ;
      LAYER li1 ;
        RECT 209.920 4451.135 210.090 4451.220 ;
        RECT 201.760 4451.075 202.655 4451.135 ;
        RECT 201.930 4450.905 202.655 4451.075 ;
        RECT 201.760 4450.845 202.655 4450.905 ;
        RECT 203.315 4451.075 205.815 4451.135 ;
        RECT 203.315 4450.905 204.480 4451.075 ;
        RECT 204.650 4450.905 205.815 4451.075 ;
        RECT 203.315 4450.845 205.815 4450.905 ;
        RECT 201.760 4450.615 201.930 4450.845 ;
        RECT 204.480 4450.615 204.650 4450.845 ;
        RECT 201.760 4450.285 201.930 4450.445 ;
        RECT 204.480 4450.285 204.650 4450.445 ;
        RECT 204.820 4450.335 205.840 4450.665 ;
        RECT 201.760 4450.155 202.730 4450.285 ;
        RECT 201.930 4449.985 202.730 4450.155 ;
        RECT 201.760 4449.955 202.730 4449.985 ;
        RECT 203.330 4450.165 204.650 4450.285 ;
        RECT 203.330 4450.155 205.450 4450.165 ;
        RECT 203.330 4449.985 204.480 4450.155 ;
        RECT 204.650 4449.995 205.450 4450.155 ;
        RECT 203.330 4449.955 204.650 4449.985 ;
        RECT 201.760 4449.695 201.930 4449.955 ;
      LAYER li1 ;
        RECT 202.100 4449.615 204.310 4449.785 ;
      LAYER li1 ;
        RECT 204.480 4449.695 204.650 4449.955 ;
        RECT 205.670 4449.825 205.840 4450.335 ;
      LAYER li1 ;
        RECT 202.580 4449.530 203.460 4449.615 ;
      LAYER li1 ;
        RECT 201.760 4449.445 201.930 4449.525 ;
        RECT 201.760 4449.235 202.410 4449.445 ;
        RECT 201.930 4449.115 202.410 4449.235 ;
        RECT 201.760 4448.775 201.930 4449.065 ;
      LAYER li1 ;
        RECT 202.580 4448.945 202.750 4449.530 ;
        RECT 202.100 4448.775 202.750 4448.945 ;
      LAYER li1 ;
        RECT 201.760 4448.315 202.410 4448.605 ;
        RECT 201.930 4448.275 202.410 4448.315 ;
        RECT 201.760 4447.855 201.930 4448.145 ;
      LAYER li1 ;
        RECT 202.580 4448.105 202.750 4448.775 ;
        RECT 202.100 4447.935 202.750 4448.105 ;
      LAYER li1 ;
        RECT 201.930 4447.685 202.410 4447.765 ;
        RECT 201.760 4447.435 202.410 4447.685 ;
        RECT 201.760 4447.395 201.930 4447.435 ;
      LAYER li1 ;
        RECT 202.580 4447.265 202.750 4447.935 ;
      LAYER li1 ;
        RECT 201.760 4446.935 201.930 4447.225 ;
      LAYER li1 ;
        RECT 202.100 4447.095 202.750 4447.265 ;
      LAYER li1 ;
        RECT 201.930 4446.765 202.410 4446.925 ;
        RECT 202.920 4446.835 203.090 4449.285 ;
      LAYER li1 ;
        RECT 203.290 4448.945 203.460 4449.530 ;
      LAYER li1 ;
        RECT 204.480 4449.445 204.650 4449.525 ;
        RECT 204.820 4449.495 205.840 4449.825 ;
      LAYER li1 ;
        RECT 206.010 4449.520 206.210 4451.110 ;
      LAYER li1 ;
        RECT 206.475 4451.075 208.095 4451.135 ;
        RECT 206.475 4450.905 207.200 4451.075 ;
        RECT 207.370 4450.905 208.095 4451.075 ;
        RECT 206.475 4450.845 208.095 4450.905 ;
        RECT 208.755 4451.075 210.090 4451.135 ;
        RECT 208.755 4450.905 209.920 4451.075 ;
        RECT 208.755 4450.845 210.090 4450.905 ;
        RECT 207.200 4450.615 207.370 4450.845 ;
        RECT 209.920 4450.760 210.090 4450.845 ;
        RECT 206.380 4450.415 207.030 4450.585 ;
        RECT 206.380 4449.745 206.550 4450.415 ;
        RECT 207.200 4450.245 207.370 4450.445 ;
        RECT 206.720 4450.155 207.370 4450.245 ;
        RECT 206.720 4449.985 207.200 4450.155 ;
        RECT 206.720 4449.915 207.370 4449.985 ;
        RECT 206.380 4449.575 207.025 4449.745 ;
        RECT 207.200 4449.695 207.370 4449.915 ;
        RECT 203.680 4449.325 204.650 4449.445 ;
        RECT 205.670 4449.340 205.840 4449.495 ;
        RECT 206.380 4449.340 206.550 4449.575 ;
        RECT 207.200 4449.405 207.370 4449.525 ;
        RECT 203.680 4449.235 205.450 4449.325 ;
        RECT 203.680 4449.115 204.480 4449.235 ;
        RECT 204.650 4449.155 205.450 4449.235 ;
        RECT 205.670 4449.165 206.550 4449.340 ;
        RECT 206.720 4449.235 207.370 4449.405 ;
      LAYER li1 ;
        RECT 203.290 4448.775 204.310 4448.945 ;
      LAYER li1 ;
        RECT 204.480 4448.775 204.650 4449.065 ;
      LAYER li1 ;
        RECT 203.290 4448.105 203.460 4448.775 ;
        RECT 204.820 4448.735 205.840 4448.905 ;
      LAYER li1 ;
        RECT 203.680 4448.565 204.650 4448.605 ;
        RECT 203.680 4448.315 205.450 4448.565 ;
        RECT 203.680 4448.275 204.480 4448.315 ;
        RECT 204.650 4448.235 205.450 4448.315 ;
      LAYER li1 ;
        RECT 203.290 4447.935 204.310 4448.105 ;
        RECT 203.290 4447.265 203.460 4447.935 ;
      LAYER li1 ;
        RECT 204.480 4447.855 204.650 4448.145 ;
      LAYER li1 ;
        RECT 205.670 4448.065 205.840 4448.735 ;
        RECT 204.820 4447.895 205.840 4448.065 ;
      LAYER li1 ;
        RECT 203.680 4447.685 204.480 4447.765 ;
        RECT 204.650 4447.685 205.450 4447.725 ;
        RECT 203.680 4447.435 205.450 4447.685 ;
        RECT 204.480 4447.395 205.450 4447.435 ;
      LAYER li1 ;
        RECT 203.290 4447.095 204.310 4447.265 ;
        RECT 205.670 4447.225 205.840 4447.895 ;
      LAYER li1 ;
        RECT 204.480 4446.935 204.650 4447.225 ;
      LAYER li1 ;
        RECT 204.820 4447.055 205.840 4447.225 ;
      LAYER li1 ;
        RECT 201.760 4446.595 202.410 4446.765 ;
        RECT 202.580 4446.660 203.460 4446.835 ;
        RECT 203.680 4446.765 204.480 4446.845 ;
        RECT 204.650 4446.765 205.450 4446.885 ;
        RECT 203.680 4446.675 205.450 4446.765 ;
        RECT 201.760 4446.475 201.930 4446.595 ;
        RECT 202.580 4446.425 202.750 4446.660 ;
        RECT 203.290 4446.505 203.460 4446.660 ;
        RECT 204.480 4446.555 205.450 4446.675 ;
        RECT 201.760 4446.085 201.930 4446.305 ;
        RECT 202.105 4446.255 202.750 4446.425 ;
        RECT 201.760 4446.015 202.410 4446.085 ;
        RECT 201.930 4445.845 202.410 4446.015 ;
        RECT 201.760 4445.755 202.410 4445.845 ;
        RECT 201.760 4445.555 201.930 4445.755 ;
        RECT 202.580 4445.585 202.750 4446.255 ;
        RECT 202.100 4445.415 202.750 4445.585 ;
        RECT 201.760 4445.155 201.930 4445.385 ;
      LAYER li1 ;
        RECT 202.920 4445.380 203.120 4446.480 ;
      LAYER li1 ;
        RECT 203.290 4446.175 204.310 4446.505 ;
        RECT 204.480 4446.475 204.650 4446.555 ;
      LAYER li1 ;
        RECT 205.670 4446.470 205.840 4447.055 ;
      LAYER li1 ;
        RECT 206.040 4446.715 206.210 4449.165 ;
        RECT 206.720 4449.075 207.200 4449.235 ;
      LAYER li1 ;
        RECT 207.370 4449.090 207.915 4450.675 ;
        RECT 206.380 4448.735 207.030 4448.905 ;
      LAYER li1 ;
        RECT 207.200 4448.775 207.370 4449.065 ;
      LAYER li1 ;
        RECT 207.370 4448.750 208.745 4449.090 ;
        RECT 206.380 4448.065 206.550 4448.735 ;
      LAYER li1 ;
        RECT 207.200 4448.565 207.370 4448.605 ;
        RECT 206.720 4448.315 207.370 4448.565 ;
        RECT 206.720 4448.235 207.200 4448.315 ;
      LAYER li1 ;
        RECT 206.380 4447.895 207.030 4448.065 ;
        RECT 206.380 4447.225 206.550 4447.895 ;
      LAYER li1 ;
        RECT 207.200 4447.855 207.370 4448.145 ;
        RECT 206.720 4447.685 207.200 4447.725 ;
        RECT 206.720 4447.395 207.370 4447.685 ;
      LAYER li1 ;
        RECT 206.380 4447.055 207.030 4447.225 ;
        RECT 206.380 4446.470 206.550 4447.055 ;
      LAYER li1 ;
        RECT 207.200 4446.935 207.370 4447.225 ;
        RECT 206.720 4446.765 207.200 4446.885 ;
        RECT 206.720 4446.555 207.370 4446.765 ;
        RECT 207.200 4446.475 207.370 4446.555 ;
      LAYER li1 ;
        RECT 205.670 4446.385 206.550 4446.470 ;
      LAYER li1 ;
        RECT 203.290 4445.665 203.460 4446.175 ;
        RECT 204.480 4446.045 204.650 4446.305 ;
      LAYER li1 ;
        RECT 204.820 4446.215 207.030 4446.385 ;
      LAYER li1 ;
        RECT 207.200 4446.045 207.370 4446.305 ;
        RECT 204.480 4446.015 205.800 4446.045 ;
        RECT 203.680 4445.845 204.480 4446.005 ;
        RECT 204.650 4445.845 205.800 4446.015 ;
        RECT 203.680 4445.835 205.800 4445.845 ;
        RECT 204.480 4445.715 205.800 4445.835 ;
        RECT 206.400 4446.015 207.370 4446.045 ;
        RECT 206.400 4445.845 207.200 4446.015 ;
        RECT 206.400 4445.715 207.370 4445.845 ;
        RECT 203.290 4445.335 204.310 4445.665 ;
        RECT 204.480 4445.555 204.650 4445.715 ;
        RECT 207.200 4445.555 207.370 4445.715 ;
        RECT 204.480 4445.155 204.650 4445.385 ;
        RECT 207.200 4445.155 207.370 4445.385 ;
      LAYER li1 ;
        RECT 207.370 4445.330 207.915 4448.750 ;
      LAYER li1 ;
        RECT 209.920 4445.155 210.090 4445.240 ;
        RECT 201.760 4445.095 202.655 4445.155 ;
        RECT 201.930 4444.925 202.655 4445.095 ;
        RECT 201.760 4444.865 202.655 4444.925 ;
        RECT 203.315 4445.095 205.815 4445.155 ;
        RECT 203.315 4444.925 204.480 4445.095 ;
        RECT 204.650 4444.925 205.815 4445.095 ;
        RECT 203.315 4444.865 205.815 4444.925 ;
        RECT 201.760 4444.635 201.930 4444.865 ;
        RECT 204.480 4444.635 204.650 4444.865 ;
        RECT 201.760 4444.305 201.930 4444.465 ;
        RECT 204.480 4444.305 204.650 4444.465 ;
        RECT 204.820 4444.355 205.840 4444.685 ;
        RECT 201.760 4444.175 202.730 4444.305 ;
        RECT 201.930 4444.005 202.730 4444.175 ;
        RECT 201.760 4443.975 202.730 4444.005 ;
        RECT 203.330 4444.185 204.650 4444.305 ;
        RECT 203.330 4444.175 205.450 4444.185 ;
        RECT 203.330 4444.005 204.480 4444.175 ;
        RECT 204.650 4444.015 205.450 4444.175 ;
        RECT 203.330 4443.975 204.650 4444.005 ;
        RECT 201.760 4443.715 201.930 4443.975 ;
      LAYER li1 ;
        RECT 202.100 4443.635 204.310 4443.805 ;
      LAYER li1 ;
        RECT 204.480 4443.715 204.650 4443.975 ;
        RECT 205.670 4443.845 205.840 4444.355 ;
      LAYER li1 ;
        RECT 202.580 4443.550 203.460 4443.635 ;
      LAYER li1 ;
        RECT 201.760 4443.465 201.930 4443.545 ;
        RECT 201.760 4443.255 202.410 4443.465 ;
        RECT 201.930 4443.135 202.410 4443.255 ;
        RECT 201.760 4442.795 201.930 4443.085 ;
      LAYER li1 ;
        RECT 202.580 4442.965 202.750 4443.550 ;
        RECT 202.100 4442.795 202.750 4442.965 ;
      LAYER li1 ;
        RECT 201.760 4442.335 202.410 4442.625 ;
        RECT 201.930 4442.295 202.410 4442.335 ;
        RECT 201.760 4441.875 201.930 4442.165 ;
      LAYER li1 ;
        RECT 202.580 4442.125 202.750 4442.795 ;
        RECT 202.100 4441.955 202.750 4442.125 ;
      LAYER li1 ;
        RECT 201.930 4441.705 202.410 4441.785 ;
        RECT 201.760 4441.455 202.410 4441.705 ;
        RECT 201.760 4441.415 201.930 4441.455 ;
      LAYER li1 ;
        RECT 202.580 4441.285 202.750 4441.955 ;
      LAYER li1 ;
        RECT 201.760 4440.955 201.930 4441.245 ;
      LAYER li1 ;
        RECT 202.100 4441.115 202.750 4441.285 ;
      LAYER li1 ;
        RECT 201.930 4440.785 202.410 4440.945 ;
        RECT 202.920 4440.855 203.090 4443.305 ;
      LAYER li1 ;
        RECT 203.290 4442.965 203.460 4443.550 ;
      LAYER li1 ;
        RECT 204.480 4443.465 204.650 4443.545 ;
        RECT 204.820 4443.515 205.840 4443.845 ;
      LAYER li1 ;
        RECT 206.010 4443.540 206.210 4445.130 ;
      LAYER li1 ;
        RECT 206.475 4445.095 208.095 4445.155 ;
        RECT 206.475 4444.925 207.200 4445.095 ;
        RECT 207.370 4444.925 208.095 4445.095 ;
        RECT 206.475 4444.865 208.095 4444.925 ;
        RECT 208.755 4445.095 210.090 4445.155 ;
        RECT 208.755 4444.925 209.920 4445.095 ;
        RECT 208.755 4444.865 210.090 4444.925 ;
        RECT 207.200 4444.635 207.370 4444.865 ;
        RECT 209.920 4444.780 210.090 4444.865 ;
        RECT 206.380 4444.435 207.030 4444.605 ;
        RECT 206.380 4443.765 206.550 4444.435 ;
        RECT 207.200 4444.265 207.370 4444.465 ;
        RECT 206.720 4444.175 207.370 4444.265 ;
        RECT 206.720 4444.005 207.200 4444.175 ;
        RECT 206.720 4443.935 207.370 4444.005 ;
        RECT 206.380 4443.595 207.025 4443.765 ;
        RECT 207.200 4443.715 207.370 4443.935 ;
        RECT 203.680 4443.345 204.650 4443.465 ;
        RECT 205.670 4443.360 205.840 4443.515 ;
        RECT 206.380 4443.360 206.550 4443.595 ;
        RECT 207.200 4443.425 207.370 4443.545 ;
        RECT 203.680 4443.255 205.450 4443.345 ;
        RECT 203.680 4443.135 204.480 4443.255 ;
        RECT 204.650 4443.175 205.450 4443.255 ;
        RECT 205.670 4443.185 206.550 4443.360 ;
        RECT 206.720 4443.255 207.370 4443.425 ;
      LAYER li1 ;
        RECT 203.290 4442.795 204.310 4442.965 ;
      LAYER li1 ;
        RECT 204.480 4442.795 204.650 4443.085 ;
      LAYER li1 ;
        RECT 203.290 4442.125 203.460 4442.795 ;
        RECT 204.820 4442.755 205.840 4442.925 ;
      LAYER li1 ;
        RECT 203.680 4442.585 204.650 4442.625 ;
        RECT 203.680 4442.335 205.450 4442.585 ;
        RECT 203.680 4442.295 204.480 4442.335 ;
        RECT 204.650 4442.255 205.450 4442.335 ;
      LAYER li1 ;
        RECT 203.290 4441.955 204.310 4442.125 ;
        RECT 203.290 4441.285 203.460 4441.955 ;
      LAYER li1 ;
        RECT 204.480 4441.875 204.650 4442.165 ;
      LAYER li1 ;
        RECT 205.670 4442.085 205.840 4442.755 ;
        RECT 204.820 4441.915 205.840 4442.085 ;
      LAYER li1 ;
        RECT 203.680 4441.705 204.480 4441.785 ;
        RECT 204.650 4441.705 205.450 4441.745 ;
        RECT 203.680 4441.455 205.450 4441.705 ;
        RECT 204.480 4441.415 205.450 4441.455 ;
      LAYER li1 ;
        RECT 203.290 4441.115 204.310 4441.285 ;
        RECT 205.670 4441.245 205.840 4441.915 ;
      LAYER li1 ;
        RECT 204.480 4440.955 204.650 4441.245 ;
      LAYER li1 ;
        RECT 204.820 4441.075 205.840 4441.245 ;
      LAYER li1 ;
        RECT 201.760 4440.615 202.410 4440.785 ;
        RECT 202.580 4440.680 203.460 4440.855 ;
        RECT 203.680 4440.785 204.480 4440.865 ;
        RECT 204.650 4440.785 205.450 4440.905 ;
        RECT 203.680 4440.695 205.450 4440.785 ;
        RECT 201.760 4440.495 201.930 4440.615 ;
        RECT 202.580 4440.445 202.750 4440.680 ;
        RECT 203.290 4440.525 203.460 4440.680 ;
        RECT 204.480 4440.575 205.450 4440.695 ;
        RECT 201.760 4440.105 201.930 4440.325 ;
        RECT 202.105 4440.275 202.750 4440.445 ;
        RECT 201.760 4440.035 202.410 4440.105 ;
        RECT 201.930 4439.865 202.410 4440.035 ;
        RECT 201.760 4439.775 202.410 4439.865 ;
        RECT 201.760 4439.575 201.930 4439.775 ;
        RECT 202.580 4439.605 202.750 4440.275 ;
        RECT 202.100 4439.435 202.750 4439.605 ;
        RECT 201.760 4439.175 201.930 4439.405 ;
      LAYER li1 ;
        RECT 202.920 4439.400 203.120 4440.500 ;
      LAYER li1 ;
        RECT 203.290 4440.195 204.310 4440.525 ;
        RECT 204.480 4440.495 204.650 4440.575 ;
      LAYER li1 ;
        RECT 205.670 4440.490 205.840 4441.075 ;
      LAYER li1 ;
        RECT 206.040 4440.735 206.210 4443.185 ;
        RECT 206.720 4443.095 207.200 4443.255 ;
      LAYER li1 ;
        RECT 207.370 4443.110 207.915 4444.695 ;
        RECT 206.380 4442.755 207.030 4442.925 ;
      LAYER li1 ;
        RECT 207.200 4442.795 207.370 4443.085 ;
      LAYER li1 ;
        RECT 207.370 4442.770 208.745 4443.110 ;
        RECT 206.380 4442.085 206.550 4442.755 ;
      LAYER li1 ;
        RECT 207.200 4442.585 207.370 4442.625 ;
        RECT 206.720 4442.335 207.370 4442.585 ;
        RECT 206.720 4442.255 207.200 4442.335 ;
      LAYER li1 ;
        RECT 206.380 4441.915 207.030 4442.085 ;
        RECT 206.380 4441.245 206.550 4441.915 ;
      LAYER li1 ;
        RECT 207.200 4441.875 207.370 4442.165 ;
        RECT 206.720 4441.705 207.200 4441.745 ;
        RECT 206.720 4441.415 207.370 4441.705 ;
      LAYER li1 ;
        RECT 206.380 4441.075 207.030 4441.245 ;
        RECT 206.380 4440.490 206.550 4441.075 ;
      LAYER li1 ;
        RECT 207.200 4440.955 207.370 4441.245 ;
        RECT 206.720 4440.785 207.200 4440.905 ;
        RECT 206.720 4440.575 207.370 4440.785 ;
        RECT 207.200 4440.495 207.370 4440.575 ;
      LAYER li1 ;
        RECT 205.670 4440.405 206.550 4440.490 ;
      LAYER li1 ;
        RECT 203.290 4439.685 203.460 4440.195 ;
        RECT 204.480 4440.065 204.650 4440.325 ;
      LAYER li1 ;
        RECT 204.820 4440.235 207.030 4440.405 ;
      LAYER li1 ;
        RECT 207.200 4440.065 207.370 4440.325 ;
        RECT 204.480 4440.035 205.800 4440.065 ;
        RECT 203.680 4439.865 204.480 4440.025 ;
        RECT 204.650 4439.865 205.800 4440.035 ;
        RECT 203.680 4439.855 205.800 4439.865 ;
        RECT 204.480 4439.735 205.800 4439.855 ;
        RECT 206.400 4440.035 207.370 4440.065 ;
        RECT 206.400 4439.865 207.200 4440.035 ;
        RECT 206.400 4439.735 207.370 4439.865 ;
        RECT 203.290 4439.355 204.310 4439.685 ;
        RECT 204.480 4439.575 204.650 4439.735 ;
        RECT 207.200 4439.575 207.370 4439.735 ;
        RECT 204.480 4439.175 204.650 4439.405 ;
        RECT 207.200 4439.175 207.370 4439.405 ;
      LAYER li1 ;
        RECT 207.370 4439.350 207.915 4442.770 ;
      LAYER li1 ;
        RECT 209.920 4439.175 210.090 4439.260 ;
        RECT 201.760 4439.115 202.655 4439.175 ;
        RECT 201.930 4438.945 202.655 4439.115 ;
        RECT 201.760 4438.885 202.655 4438.945 ;
        RECT 203.315 4439.115 205.815 4439.175 ;
        RECT 203.315 4438.945 204.480 4439.115 ;
        RECT 204.650 4438.945 205.815 4439.115 ;
        RECT 203.315 4438.885 205.815 4438.945 ;
        RECT 206.475 4439.115 208.095 4439.175 ;
        RECT 206.475 4438.945 207.200 4439.115 ;
        RECT 207.370 4438.945 208.095 4439.115 ;
        RECT 206.475 4438.885 208.095 4438.945 ;
        RECT 208.755 4439.115 210.090 4439.175 ;
        RECT 208.755 4438.945 209.920 4439.115 ;
        RECT 208.755 4438.885 210.090 4438.945 ;
        RECT 201.760 4438.655 201.930 4438.885 ;
        RECT 204.480 4438.655 204.650 4438.885 ;
        RECT 201.760 4438.325 201.930 4438.485 ;
        RECT 204.480 4438.325 204.650 4438.485 ;
        RECT 204.820 4438.375 205.840 4438.705 ;
        RECT 207.200 4438.655 207.370 4438.885 ;
        RECT 209.920 4438.800 210.090 4438.885 ;
        RECT 201.760 4438.195 202.730 4438.325 ;
        RECT 201.930 4438.025 202.730 4438.195 ;
        RECT 201.760 4437.995 202.730 4438.025 ;
        RECT 203.330 4438.205 204.650 4438.325 ;
        RECT 203.330 4438.195 205.450 4438.205 ;
        RECT 203.330 4438.025 204.480 4438.195 ;
        RECT 204.650 4438.035 205.450 4438.195 ;
        RECT 203.330 4437.995 204.650 4438.025 ;
        RECT 201.760 4437.735 201.930 4437.995 ;
        RECT 204.480 4437.735 204.650 4437.995 ;
        RECT 205.670 4437.865 205.840 4438.375 ;
        RECT 201.760 4437.485 201.930 4437.565 ;
        RECT 204.480 4437.485 204.650 4437.565 ;
        RECT 204.820 4437.535 205.840 4437.865 ;
        RECT 201.760 4437.275 202.410 4437.485 ;
        RECT 203.680 4437.365 204.650 4437.485 ;
        RECT 205.670 4437.380 205.840 4437.535 ;
        RECT 206.380 4438.455 207.030 4438.625 ;
        RECT 206.380 4437.785 206.550 4438.455 ;
        RECT 207.200 4438.285 207.370 4438.485 ;
        RECT 206.720 4438.195 207.370 4438.285 ;
        RECT 206.720 4438.025 207.200 4438.195 ;
        RECT 206.720 4437.955 207.370 4438.025 ;
        RECT 206.380 4437.615 207.025 4437.785 ;
        RECT 207.200 4437.735 207.370 4437.955 ;
        RECT 206.380 4437.380 206.550 4437.615 ;
        RECT 207.200 4437.445 207.370 4437.565 ;
        RECT 201.930 4437.155 202.410 4437.275 ;
        RECT 201.760 4436.815 201.930 4437.105 ;
        RECT 201.760 4436.355 202.410 4436.645 ;
        RECT 201.930 4436.315 202.410 4436.355 ;
        RECT 201.760 4435.895 201.930 4436.185 ;
        RECT 201.930 4435.725 202.410 4435.805 ;
        RECT 201.760 4435.475 202.410 4435.725 ;
        RECT 201.760 4435.435 201.930 4435.475 ;
        RECT 201.760 4434.975 201.930 4435.265 ;
        RECT 201.930 4434.805 202.410 4434.965 ;
        RECT 202.920 4434.875 203.090 4437.325 ;
        RECT 203.680 4437.275 205.450 4437.365 ;
        RECT 203.680 4437.155 204.480 4437.275 ;
        RECT 204.650 4437.195 205.450 4437.275 ;
        RECT 205.670 4437.205 206.550 4437.380 ;
        RECT 206.720 4437.275 207.370 4437.445 ;
        RECT 204.480 4436.815 204.650 4437.105 ;
      LAYER li1 ;
        RECT 204.820 4436.775 205.840 4436.945 ;
      LAYER li1 ;
        RECT 203.680 4436.605 204.650 4436.645 ;
        RECT 203.680 4436.355 205.450 4436.605 ;
        RECT 203.680 4436.315 204.480 4436.355 ;
        RECT 204.650 4436.275 205.450 4436.355 ;
        RECT 204.480 4435.895 204.650 4436.185 ;
      LAYER li1 ;
        RECT 205.670 4436.105 205.840 4436.775 ;
        RECT 204.820 4435.935 205.840 4436.105 ;
      LAYER li1 ;
        RECT 203.680 4435.725 204.480 4435.805 ;
        RECT 204.650 4435.725 205.450 4435.765 ;
        RECT 203.680 4435.475 205.450 4435.725 ;
        RECT 204.480 4435.435 205.450 4435.475 ;
      LAYER li1 ;
        RECT 205.670 4435.265 205.840 4435.935 ;
      LAYER li1 ;
        RECT 204.480 4434.975 204.650 4435.265 ;
      LAYER li1 ;
        RECT 204.820 4435.095 205.840 4435.265 ;
      LAYER li1 ;
        RECT 201.760 4434.635 202.410 4434.805 ;
        RECT 202.580 4434.700 203.460 4434.875 ;
        RECT 203.680 4434.805 204.480 4434.885 ;
        RECT 204.650 4434.805 205.450 4434.925 ;
        RECT 203.680 4434.715 205.450 4434.805 ;
        RECT 201.760 4434.515 201.930 4434.635 ;
        RECT 202.580 4434.465 202.750 4434.700 ;
        RECT 203.290 4434.545 203.460 4434.700 ;
        RECT 204.480 4434.595 205.450 4434.715 ;
        RECT 201.760 4434.125 201.930 4434.345 ;
        RECT 202.105 4434.295 202.750 4434.465 ;
        RECT 201.760 4434.055 202.410 4434.125 ;
        RECT 201.930 4433.885 202.410 4434.055 ;
        RECT 201.760 4433.795 202.410 4433.885 ;
        RECT 201.760 4433.595 201.930 4433.795 ;
        RECT 202.580 4433.625 202.750 4434.295 ;
        RECT 202.100 4433.455 202.750 4433.625 ;
        RECT 201.760 4433.195 201.930 4433.425 ;
      LAYER li1 ;
        RECT 202.920 4433.420 203.120 4434.520 ;
      LAYER li1 ;
        RECT 203.290 4434.215 204.310 4434.545 ;
        RECT 204.480 4434.515 204.650 4434.595 ;
      LAYER li1 ;
        RECT 205.670 4434.510 205.840 4435.095 ;
      LAYER li1 ;
        RECT 206.040 4434.755 206.210 4437.205 ;
        RECT 206.720 4437.115 207.200 4437.275 ;
      LAYER li1 ;
        RECT 207.370 4437.130 207.915 4438.715 ;
        RECT 206.380 4436.775 207.030 4436.945 ;
      LAYER li1 ;
        RECT 207.200 4436.815 207.370 4437.105 ;
      LAYER li1 ;
        RECT 207.370 4436.790 208.745 4437.130 ;
        RECT 206.380 4436.105 206.550 4436.775 ;
      LAYER li1 ;
        RECT 207.200 4436.605 207.370 4436.645 ;
        RECT 206.720 4436.355 207.370 4436.605 ;
        RECT 206.720 4436.275 207.200 4436.355 ;
      LAYER li1 ;
        RECT 206.380 4435.935 207.030 4436.105 ;
        RECT 206.380 4435.265 206.550 4435.935 ;
      LAYER li1 ;
        RECT 207.200 4435.895 207.370 4436.185 ;
        RECT 206.720 4435.725 207.200 4435.765 ;
        RECT 206.720 4435.435 207.370 4435.725 ;
      LAYER li1 ;
        RECT 206.380 4435.095 207.030 4435.265 ;
        RECT 206.380 4434.510 206.550 4435.095 ;
      LAYER li1 ;
        RECT 207.200 4434.975 207.370 4435.265 ;
        RECT 206.720 4434.805 207.200 4434.925 ;
        RECT 206.720 4434.595 207.370 4434.805 ;
        RECT 207.200 4434.515 207.370 4434.595 ;
      LAYER li1 ;
        RECT 205.670 4434.425 206.550 4434.510 ;
      LAYER li1 ;
        RECT 203.290 4433.705 203.460 4434.215 ;
        RECT 204.480 4434.085 204.650 4434.345 ;
      LAYER li1 ;
        RECT 204.820 4434.255 207.030 4434.425 ;
      LAYER li1 ;
        RECT 207.200 4434.085 207.370 4434.345 ;
        RECT 204.480 4434.055 205.800 4434.085 ;
        RECT 203.680 4433.885 204.480 4434.045 ;
        RECT 204.650 4433.885 205.800 4434.055 ;
        RECT 203.680 4433.875 205.800 4433.885 ;
        RECT 204.480 4433.755 205.800 4433.875 ;
        RECT 206.400 4434.055 207.370 4434.085 ;
        RECT 206.400 4433.885 207.200 4434.055 ;
        RECT 206.400 4433.755 207.370 4433.885 ;
        RECT 203.290 4433.375 204.310 4433.705 ;
        RECT 204.480 4433.595 204.650 4433.755 ;
        RECT 207.200 4433.595 207.370 4433.755 ;
        RECT 204.480 4433.195 204.650 4433.425 ;
        RECT 207.200 4433.195 207.370 4433.425 ;
      LAYER li1 ;
        RECT 207.370 4433.370 207.915 4436.790 ;
      LAYER li1 ;
        RECT 209.920 4433.195 210.090 4433.280 ;
        RECT 201.760 4433.135 202.655 4433.195 ;
        RECT 201.930 4432.965 202.655 4433.135 ;
        RECT 201.760 4432.905 202.655 4432.965 ;
        RECT 203.315 4433.135 205.815 4433.195 ;
        RECT 203.315 4432.965 204.480 4433.135 ;
        RECT 204.650 4432.965 205.815 4433.135 ;
        RECT 203.315 4432.905 205.815 4432.965 ;
        RECT 206.475 4433.135 208.095 4433.195 ;
        RECT 206.475 4432.965 207.200 4433.135 ;
        RECT 207.370 4432.965 208.095 4433.135 ;
        RECT 206.475 4432.905 208.095 4432.965 ;
        RECT 208.755 4433.135 210.090 4433.195 ;
        RECT 208.755 4432.965 209.920 4433.135 ;
        RECT 208.755 4432.905 210.090 4432.965 ;
        RECT 201.760 4432.675 201.930 4432.905 ;
        RECT 204.480 4432.675 204.650 4432.905 ;
        RECT 201.760 4432.345 201.930 4432.505 ;
        RECT 204.480 4432.345 204.650 4432.505 ;
        RECT 204.820 4432.395 205.840 4432.725 ;
        RECT 207.200 4432.675 207.370 4432.905 ;
        RECT 209.920 4432.820 210.090 4432.905 ;
        RECT 201.760 4432.215 202.730 4432.345 ;
        RECT 201.930 4432.045 202.730 4432.215 ;
        RECT 201.760 4432.015 202.730 4432.045 ;
        RECT 203.330 4432.225 204.650 4432.345 ;
        RECT 203.330 4432.215 205.450 4432.225 ;
        RECT 203.330 4432.045 204.480 4432.215 ;
        RECT 204.650 4432.055 205.450 4432.215 ;
        RECT 203.330 4432.015 204.650 4432.045 ;
        RECT 201.760 4431.755 201.930 4432.015 ;
        RECT 204.480 4431.755 204.650 4432.015 ;
        RECT 205.670 4431.885 205.840 4432.395 ;
        RECT 201.760 4431.505 201.930 4431.585 ;
        RECT 204.480 4431.505 204.650 4431.585 ;
        RECT 204.820 4431.555 205.840 4431.885 ;
        RECT 201.760 4431.295 202.410 4431.505 ;
        RECT 203.680 4431.385 204.650 4431.505 ;
        RECT 205.670 4431.400 205.840 4431.555 ;
        RECT 206.380 4432.475 207.030 4432.645 ;
        RECT 206.380 4431.805 206.550 4432.475 ;
        RECT 207.200 4432.305 207.370 4432.505 ;
        RECT 206.720 4432.215 207.370 4432.305 ;
        RECT 206.720 4432.045 207.200 4432.215 ;
        RECT 206.720 4431.975 207.370 4432.045 ;
        RECT 206.380 4431.635 207.025 4431.805 ;
        RECT 207.200 4431.755 207.370 4431.975 ;
        RECT 206.380 4431.400 206.550 4431.635 ;
        RECT 207.200 4431.465 207.370 4431.585 ;
        RECT 201.930 4431.175 202.410 4431.295 ;
        RECT 201.760 4430.835 201.930 4431.125 ;
        RECT 201.760 4430.375 202.410 4430.665 ;
        RECT 201.930 4430.335 202.410 4430.375 ;
        RECT 201.760 4429.915 201.930 4430.205 ;
        RECT 201.930 4429.745 202.410 4429.825 ;
        RECT 201.760 4429.495 202.410 4429.745 ;
        RECT 201.760 4429.455 201.930 4429.495 ;
        RECT 201.760 4428.995 201.930 4429.285 ;
        RECT 201.930 4428.825 202.410 4428.985 ;
        RECT 202.920 4428.895 203.090 4431.345 ;
        RECT 203.680 4431.295 205.450 4431.385 ;
        RECT 203.680 4431.175 204.480 4431.295 ;
        RECT 204.650 4431.215 205.450 4431.295 ;
        RECT 205.670 4431.225 206.550 4431.400 ;
        RECT 206.720 4431.295 207.370 4431.465 ;
        RECT 204.480 4430.835 204.650 4431.125 ;
      LAYER li1 ;
        RECT 204.820 4430.795 205.840 4430.965 ;
      LAYER li1 ;
        RECT 203.680 4430.625 204.650 4430.665 ;
        RECT 203.680 4430.375 205.450 4430.625 ;
        RECT 203.680 4430.335 204.480 4430.375 ;
        RECT 204.650 4430.295 205.450 4430.375 ;
        RECT 204.480 4429.915 204.650 4430.205 ;
      LAYER li1 ;
        RECT 205.670 4430.125 205.840 4430.795 ;
        RECT 204.820 4429.955 205.840 4430.125 ;
      LAYER li1 ;
        RECT 203.680 4429.745 204.480 4429.825 ;
        RECT 204.650 4429.745 205.450 4429.785 ;
        RECT 203.680 4429.495 205.450 4429.745 ;
        RECT 204.480 4429.455 205.450 4429.495 ;
      LAYER li1 ;
        RECT 205.670 4429.285 205.840 4429.955 ;
      LAYER li1 ;
        RECT 204.480 4428.995 204.650 4429.285 ;
      LAYER li1 ;
        RECT 204.820 4429.115 205.840 4429.285 ;
      LAYER li1 ;
        RECT 201.760 4428.655 202.410 4428.825 ;
        RECT 202.580 4428.720 203.460 4428.895 ;
        RECT 203.680 4428.825 204.480 4428.905 ;
        RECT 204.650 4428.825 205.450 4428.945 ;
        RECT 203.680 4428.735 205.450 4428.825 ;
        RECT 201.760 4428.535 201.930 4428.655 ;
        RECT 202.580 4428.485 202.750 4428.720 ;
        RECT 203.290 4428.565 203.460 4428.720 ;
        RECT 204.480 4428.615 205.450 4428.735 ;
        RECT 201.760 4428.145 201.930 4428.365 ;
        RECT 202.105 4428.315 202.750 4428.485 ;
        RECT 201.760 4428.075 202.410 4428.145 ;
        RECT 201.930 4427.905 202.410 4428.075 ;
        RECT 201.760 4427.815 202.410 4427.905 ;
        RECT 201.760 4427.615 201.930 4427.815 ;
        RECT 202.580 4427.645 202.750 4428.315 ;
        RECT 202.100 4427.475 202.750 4427.645 ;
        RECT 201.760 4427.215 201.930 4427.445 ;
      LAYER li1 ;
        RECT 202.920 4427.440 203.120 4428.540 ;
      LAYER li1 ;
        RECT 203.290 4428.235 204.310 4428.565 ;
        RECT 204.480 4428.535 204.650 4428.615 ;
      LAYER li1 ;
        RECT 205.670 4428.530 205.840 4429.115 ;
      LAYER li1 ;
        RECT 206.040 4428.775 206.210 4431.225 ;
        RECT 206.720 4431.135 207.200 4431.295 ;
      LAYER li1 ;
        RECT 207.370 4431.150 207.915 4432.735 ;
        RECT 206.380 4430.795 207.030 4430.965 ;
      LAYER li1 ;
        RECT 207.200 4430.835 207.370 4431.125 ;
      LAYER li1 ;
        RECT 207.370 4430.810 208.745 4431.150 ;
        RECT 206.380 4430.125 206.550 4430.795 ;
      LAYER li1 ;
        RECT 207.200 4430.625 207.370 4430.665 ;
        RECT 206.720 4430.375 207.370 4430.625 ;
        RECT 206.720 4430.295 207.200 4430.375 ;
      LAYER li1 ;
        RECT 206.380 4429.955 207.030 4430.125 ;
        RECT 206.380 4429.285 206.550 4429.955 ;
      LAYER li1 ;
        RECT 207.200 4429.915 207.370 4430.205 ;
        RECT 206.720 4429.745 207.200 4429.785 ;
        RECT 206.720 4429.455 207.370 4429.745 ;
      LAYER li1 ;
        RECT 206.380 4429.115 207.030 4429.285 ;
        RECT 206.380 4428.530 206.550 4429.115 ;
      LAYER li1 ;
        RECT 207.200 4428.995 207.370 4429.285 ;
        RECT 206.720 4428.825 207.200 4428.945 ;
        RECT 206.720 4428.615 207.370 4428.825 ;
        RECT 207.200 4428.535 207.370 4428.615 ;
      LAYER li1 ;
        RECT 205.670 4428.445 206.550 4428.530 ;
      LAYER li1 ;
        RECT 203.290 4427.725 203.460 4428.235 ;
        RECT 204.480 4428.105 204.650 4428.365 ;
      LAYER li1 ;
        RECT 204.820 4428.275 207.030 4428.445 ;
      LAYER li1 ;
        RECT 207.200 4428.105 207.370 4428.365 ;
        RECT 204.480 4428.075 205.800 4428.105 ;
        RECT 203.680 4427.905 204.480 4428.065 ;
        RECT 204.650 4427.905 205.800 4428.075 ;
        RECT 203.680 4427.895 205.800 4427.905 ;
        RECT 204.480 4427.775 205.800 4427.895 ;
        RECT 206.400 4428.075 207.370 4428.105 ;
        RECT 206.400 4427.905 207.200 4428.075 ;
        RECT 206.400 4427.775 207.370 4427.905 ;
        RECT 203.290 4427.395 204.310 4427.725 ;
        RECT 204.480 4427.615 204.650 4427.775 ;
        RECT 207.200 4427.615 207.370 4427.775 ;
        RECT 204.480 4427.215 204.650 4427.445 ;
        RECT 207.200 4427.215 207.370 4427.445 ;
      LAYER li1 ;
        RECT 207.370 4427.390 207.915 4430.810 ;
      LAYER li1 ;
        RECT 209.920 4427.215 210.090 4427.300 ;
        RECT 201.760 4427.155 202.655 4427.215 ;
        RECT 201.930 4426.985 202.655 4427.155 ;
        RECT 201.760 4426.925 202.655 4426.985 ;
        RECT 203.315 4427.155 205.815 4427.215 ;
        RECT 203.315 4426.985 204.480 4427.155 ;
        RECT 204.650 4426.985 205.815 4427.155 ;
        RECT 203.315 4426.925 205.815 4426.985 ;
        RECT 206.475 4427.155 208.095 4427.215 ;
        RECT 206.475 4426.985 207.200 4427.155 ;
        RECT 207.370 4426.985 208.095 4427.155 ;
        RECT 206.475 4426.925 208.095 4426.985 ;
        RECT 208.755 4427.155 210.090 4427.215 ;
        RECT 208.755 4426.985 209.920 4427.155 ;
        RECT 208.755 4426.925 210.090 4426.985 ;
        RECT 201.760 4426.840 201.930 4426.925 ;
        RECT 204.480 4426.840 204.650 4426.925 ;
        RECT 207.200 4426.840 207.370 4426.925 ;
        RECT 209.920 4426.840 210.090 4426.925 ;
        RECT 3377.780 3638.315 3377.950 3638.400 ;
        RECT 3380.500 3638.315 3380.670 3638.400 ;
        RECT 3383.220 3638.315 3383.390 3638.400 ;
        RECT 3385.940 3638.315 3386.110 3638.400 ;
        RECT 3377.780 3638.255 3379.115 3638.315 ;
        RECT 3377.950 3638.085 3379.115 3638.255 ;
        RECT 3377.780 3638.025 3379.115 3638.085 ;
        RECT 3379.775 3638.255 3381.395 3638.315 ;
        RECT 3379.775 3638.085 3380.500 3638.255 ;
        RECT 3380.670 3638.085 3381.395 3638.255 ;
        RECT 3379.775 3638.025 3381.395 3638.085 ;
        RECT 3377.780 3637.940 3377.950 3638.025 ;
      LAYER li1 ;
        RECT 3379.955 3636.270 3380.500 3637.855 ;
      LAYER li1 ;
        RECT 3380.500 3637.795 3380.670 3638.025 ;
        RECT 3380.500 3637.425 3380.670 3637.625 ;
        RECT 3380.840 3637.595 3381.490 3637.765 ;
        RECT 3380.500 3637.335 3381.150 3637.425 ;
        RECT 3380.670 3637.165 3381.150 3637.335 ;
        RECT 3380.500 3637.095 3381.150 3637.165 ;
        RECT 3380.500 3636.875 3380.670 3637.095 ;
        RECT 3381.320 3636.925 3381.490 3637.595 ;
        RECT 3380.845 3636.755 3381.490 3636.925 ;
        RECT 3380.500 3636.585 3380.670 3636.705 ;
        RECT 3380.500 3636.415 3381.150 3636.585 ;
      LAYER li1 ;
        RECT 3379.125 3635.930 3380.500 3636.270 ;
      LAYER li1 ;
        RECT 3380.670 3636.255 3381.150 3636.415 ;
        RECT 3381.320 3636.520 3381.490 3636.755 ;
      LAYER li1 ;
        RECT 3381.660 3636.700 3381.860 3638.290 ;
      LAYER li1 ;
        RECT 3382.055 3638.255 3384.555 3638.315 ;
        RECT 3382.055 3638.085 3383.220 3638.255 ;
        RECT 3383.390 3638.085 3384.555 3638.255 ;
        RECT 3382.055 3638.025 3384.555 3638.085 ;
        RECT 3385.215 3638.255 3386.110 3638.315 ;
        RECT 3385.215 3638.085 3385.940 3638.255 ;
        RECT 3385.215 3638.025 3386.110 3638.085 ;
        RECT 3382.030 3637.515 3383.050 3637.845 ;
        RECT 3383.220 3637.795 3383.390 3638.025 ;
        RECT 3385.940 3637.795 3386.110 3638.025 ;
        RECT 3382.030 3637.005 3382.200 3637.515 ;
        RECT 3383.220 3637.465 3383.390 3637.625 ;
        RECT 3385.940 3637.465 3386.110 3637.625 ;
        RECT 3383.220 3637.345 3384.540 3637.465 ;
        RECT 3382.420 3637.335 3384.540 3637.345 ;
        RECT 3382.420 3637.175 3383.220 3637.335 ;
        RECT 3383.390 3637.165 3384.540 3637.335 ;
        RECT 3383.220 3637.135 3384.540 3637.165 ;
        RECT 3385.140 3637.335 3386.110 3637.465 ;
        RECT 3385.140 3637.165 3385.940 3637.335 ;
        RECT 3385.140 3637.135 3386.110 3637.165 ;
        RECT 3382.030 3636.675 3383.050 3637.005 ;
        RECT 3383.220 3636.875 3383.390 3637.135 ;
      LAYER li1 ;
        RECT 3383.560 3636.795 3385.770 3636.965 ;
      LAYER li1 ;
        RECT 3385.940 3636.875 3386.110 3637.135 ;
      LAYER li1 ;
        RECT 3384.410 3636.710 3385.290 3636.795 ;
      LAYER li1 ;
        RECT 3382.030 3636.520 3382.200 3636.675 ;
        RECT 3381.320 3636.345 3382.200 3636.520 ;
        RECT 3383.220 3636.625 3383.390 3636.705 ;
        RECT 3383.220 3636.505 3384.190 3636.625 ;
        RECT 3382.420 3636.415 3384.190 3636.505 ;
        RECT 3380.500 3635.955 3380.670 3636.245 ;
      LAYER li1 ;
        RECT 3379.955 3632.510 3380.500 3635.930 ;
        RECT 3380.840 3635.915 3381.490 3636.085 ;
      LAYER li1 ;
        RECT 3380.500 3635.745 3380.670 3635.785 ;
        RECT 3380.500 3635.495 3381.150 3635.745 ;
        RECT 3380.670 3635.415 3381.150 3635.495 ;
        RECT 3380.500 3635.035 3380.670 3635.325 ;
      LAYER li1 ;
        RECT 3381.320 3635.245 3381.490 3635.915 ;
        RECT 3380.840 3635.075 3381.490 3635.245 ;
      LAYER li1 ;
        RECT 3380.670 3634.865 3381.150 3634.905 ;
        RECT 3380.500 3634.575 3381.150 3634.865 ;
      LAYER li1 ;
        RECT 3381.320 3634.405 3381.490 3635.075 ;
      LAYER li1 ;
        RECT 3380.500 3634.115 3380.670 3634.405 ;
      LAYER li1 ;
        RECT 3380.840 3634.235 3381.490 3634.405 ;
      LAYER li1 ;
        RECT 3380.670 3633.945 3381.150 3634.065 ;
        RECT 3380.500 3633.735 3381.150 3633.945 ;
        RECT 3380.500 3633.655 3380.670 3633.735 ;
      LAYER li1 ;
        RECT 3381.320 3633.650 3381.490 3634.235 ;
      LAYER li1 ;
        RECT 3381.660 3633.895 3381.830 3636.345 ;
        RECT 3382.420 3636.335 3383.220 3636.415 ;
        RECT 3383.390 3636.295 3384.190 3636.415 ;
      LAYER li1 ;
        RECT 3382.030 3635.915 3383.050 3636.085 ;
      LAYER li1 ;
        RECT 3383.220 3635.955 3383.390 3636.245 ;
      LAYER li1 ;
        RECT 3384.410 3636.125 3384.580 3636.710 ;
        RECT 3383.560 3635.955 3384.580 3636.125 ;
        RECT 3382.030 3635.245 3382.200 3635.915 ;
      LAYER li1 ;
        RECT 3383.220 3635.745 3384.190 3635.785 ;
        RECT 3382.420 3635.495 3384.190 3635.745 ;
        RECT 3382.420 3635.415 3383.220 3635.495 ;
        RECT 3383.390 3635.455 3384.190 3635.495 ;
      LAYER li1 ;
        RECT 3382.030 3635.075 3383.050 3635.245 ;
        RECT 3382.030 3634.405 3382.200 3635.075 ;
      LAYER li1 ;
        RECT 3383.220 3635.035 3383.390 3635.325 ;
      LAYER li1 ;
        RECT 3384.410 3635.285 3384.580 3635.955 ;
        RECT 3383.560 3635.115 3384.580 3635.285 ;
      LAYER li1 ;
        RECT 3382.420 3634.865 3383.220 3634.905 ;
        RECT 3383.390 3634.865 3384.190 3634.945 ;
        RECT 3382.420 3634.615 3384.190 3634.865 ;
        RECT 3382.420 3634.575 3383.390 3634.615 ;
      LAYER li1 ;
        RECT 3384.410 3634.445 3384.580 3635.115 ;
        RECT 3382.030 3634.235 3383.050 3634.405 ;
        RECT 3382.030 3633.650 3382.200 3634.235 ;
      LAYER li1 ;
        RECT 3383.220 3634.115 3383.390 3634.405 ;
      LAYER li1 ;
        RECT 3383.560 3634.275 3384.580 3634.445 ;
      LAYER li1 ;
        RECT 3382.420 3633.945 3383.220 3634.065 ;
        RECT 3383.390 3633.945 3384.190 3634.025 ;
        RECT 3384.780 3634.015 3384.950 3636.465 ;
      LAYER li1 ;
        RECT 3385.120 3636.125 3385.290 3636.710 ;
      LAYER li1 ;
        RECT 3385.940 3636.625 3386.110 3636.705 ;
        RECT 3385.460 3636.415 3386.110 3636.625 ;
        RECT 3385.460 3636.295 3385.940 3636.415 ;
      LAYER li1 ;
        RECT 3385.120 3635.955 3385.770 3636.125 ;
      LAYER li1 ;
        RECT 3385.940 3635.955 3386.110 3636.245 ;
      LAYER li1 ;
        RECT 3385.120 3635.285 3385.290 3635.955 ;
      LAYER li1 ;
        RECT 3385.460 3635.495 3386.110 3635.785 ;
        RECT 3385.460 3635.455 3385.940 3635.495 ;
      LAYER li1 ;
        RECT 3385.120 3635.115 3385.770 3635.285 ;
        RECT 3385.120 3634.445 3385.290 3635.115 ;
      LAYER li1 ;
        RECT 3385.940 3635.035 3386.110 3635.325 ;
        RECT 3385.460 3634.865 3385.940 3634.945 ;
        RECT 3385.460 3634.615 3386.110 3634.865 ;
        RECT 3385.940 3634.575 3386.110 3634.615 ;
      LAYER li1 ;
        RECT 3385.120 3634.275 3385.770 3634.445 ;
      LAYER li1 ;
        RECT 3385.940 3634.115 3386.110 3634.405 ;
        RECT 3382.420 3633.855 3384.190 3633.945 ;
        RECT 3382.420 3633.735 3383.390 3633.855 ;
        RECT 3383.220 3633.655 3383.390 3633.735 ;
        RECT 3384.410 3633.840 3385.290 3634.015 ;
        RECT 3384.410 3633.685 3384.580 3633.840 ;
      LAYER li1 ;
        RECT 3381.320 3633.565 3382.200 3633.650 ;
      LAYER li1 ;
        RECT 3380.500 3633.225 3380.670 3633.485 ;
      LAYER li1 ;
        RECT 3380.840 3633.395 3383.050 3633.565 ;
      LAYER li1 ;
        RECT 3383.220 3633.225 3383.390 3633.485 ;
        RECT 3383.560 3633.355 3384.580 3633.685 ;
        RECT 3380.500 3633.195 3381.470 3633.225 ;
        RECT 3380.670 3633.025 3381.470 3633.195 ;
        RECT 3380.500 3632.895 3381.470 3633.025 ;
        RECT 3382.070 3633.195 3383.390 3633.225 ;
        RECT 3382.070 3633.025 3383.220 3633.195 ;
        RECT 3383.390 3633.025 3384.190 3633.185 ;
        RECT 3382.070 3633.015 3384.190 3633.025 ;
        RECT 3382.070 3632.895 3383.390 3633.015 ;
        RECT 3380.500 3632.735 3380.670 3632.895 ;
        RECT 3383.220 3632.735 3383.390 3632.895 ;
        RECT 3384.410 3632.845 3384.580 3633.355 ;
        RECT 3377.780 3632.335 3377.950 3632.420 ;
        RECT 3380.500 3632.335 3380.670 3632.565 ;
        RECT 3383.220 3632.335 3383.390 3632.565 ;
        RECT 3383.560 3632.515 3384.580 3632.845 ;
      LAYER li1 ;
        RECT 3384.750 3632.560 3384.950 3633.660 ;
      LAYER li1 ;
        RECT 3385.120 3633.605 3385.290 3633.840 ;
        RECT 3385.460 3633.945 3385.940 3634.105 ;
        RECT 3385.460 3633.775 3386.110 3633.945 ;
        RECT 3385.940 3633.655 3386.110 3633.775 ;
        RECT 3385.120 3633.435 3385.765 3633.605 ;
        RECT 3385.120 3632.765 3385.290 3633.435 ;
        RECT 3385.940 3633.265 3386.110 3633.485 ;
        RECT 3385.460 3633.195 3386.110 3633.265 ;
        RECT 3385.460 3633.025 3385.940 3633.195 ;
        RECT 3385.460 3632.935 3386.110 3633.025 ;
        RECT 3385.120 3632.595 3385.770 3632.765 ;
        RECT 3385.940 3632.735 3386.110 3632.935 ;
        RECT 3385.940 3632.335 3386.110 3632.565 ;
        RECT 3377.780 3632.275 3379.115 3632.335 ;
        RECT 3377.950 3632.105 3379.115 3632.275 ;
        RECT 3377.780 3632.045 3379.115 3632.105 ;
        RECT 3379.775 3632.275 3381.395 3632.335 ;
        RECT 3379.775 3632.105 3380.500 3632.275 ;
        RECT 3380.670 3632.105 3381.395 3632.275 ;
        RECT 3379.775 3632.045 3381.395 3632.105 ;
        RECT 3377.780 3631.960 3377.950 3632.045 ;
      LAYER li1 ;
        RECT 3379.955 3630.290 3380.500 3631.875 ;
      LAYER li1 ;
        RECT 3380.500 3631.815 3380.670 3632.045 ;
        RECT 3380.500 3631.445 3380.670 3631.645 ;
        RECT 3380.840 3631.615 3381.490 3631.785 ;
        RECT 3380.500 3631.355 3381.150 3631.445 ;
        RECT 3380.670 3631.185 3381.150 3631.355 ;
        RECT 3380.500 3631.115 3381.150 3631.185 ;
        RECT 3380.500 3630.895 3380.670 3631.115 ;
        RECT 3381.320 3630.945 3381.490 3631.615 ;
        RECT 3380.845 3630.775 3381.490 3630.945 ;
        RECT 3380.500 3630.605 3380.670 3630.725 ;
        RECT 3380.500 3630.435 3381.150 3630.605 ;
      LAYER li1 ;
        RECT 3379.125 3629.950 3380.500 3630.290 ;
      LAYER li1 ;
        RECT 3380.670 3630.275 3381.150 3630.435 ;
        RECT 3381.320 3630.540 3381.490 3630.775 ;
      LAYER li1 ;
        RECT 3381.660 3630.720 3381.860 3632.310 ;
      LAYER li1 ;
        RECT 3382.055 3632.275 3384.555 3632.335 ;
        RECT 3382.055 3632.105 3383.220 3632.275 ;
        RECT 3383.390 3632.105 3384.555 3632.275 ;
        RECT 3382.055 3632.045 3384.555 3632.105 ;
        RECT 3385.215 3632.275 3386.110 3632.335 ;
        RECT 3385.215 3632.105 3385.940 3632.275 ;
        RECT 3385.215 3632.045 3386.110 3632.105 ;
        RECT 3382.030 3631.535 3383.050 3631.865 ;
        RECT 3383.220 3631.815 3383.390 3632.045 ;
        RECT 3385.940 3631.815 3386.110 3632.045 ;
        RECT 3382.030 3631.025 3382.200 3631.535 ;
        RECT 3383.220 3631.485 3383.390 3631.645 ;
        RECT 3385.940 3631.485 3386.110 3631.645 ;
        RECT 3383.220 3631.365 3384.540 3631.485 ;
        RECT 3382.420 3631.355 3384.540 3631.365 ;
        RECT 3382.420 3631.195 3383.220 3631.355 ;
        RECT 3383.390 3631.185 3384.540 3631.355 ;
        RECT 3383.220 3631.155 3384.540 3631.185 ;
        RECT 3385.140 3631.355 3386.110 3631.485 ;
        RECT 3385.140 3631.185 3385.940 3631.355 ;
        RECT 3385.140 3631.155 3386.110 3631.185 ;
        RECT 3382.030 3630.695 3383.050 3631.025 ;
        RECT 3383.220 3630.895 3383.390 3631.155 ;
      LAYER li1 ;
        RECT 3383.560 3630.815 3385.770 3630.985 ;
      LAYER li1 ;
        RECT 3385.940 3630.895 3386.110 3631.155 ;
      LAYER li1 ;
        RECT 3384.410 3630.730 3385.290 3630.815 ;
      LAYER li1 ;
        RECT 3382.030 3630.540 3382.200 3630.695 ;
        RECT 3381.320 3630.365 3382.200 3630.540 ;
        RECT 3383.220 3630.645 3383.390 3630.725 ;
        RECT 3383.220 3630.525 3384.190 3630.645 ;
        RECT 3382.420 3630.435 3384.190 3630.525 ;
        RECT 3380.500 3629.975 3380.670 3630.265 ;
      LAYER li1 ;
        RECT 3379.955 3626.530 3380.500 3629.950 ;
        RECT 3380.840 3629.935 3381.490 3630.105 ;
      LAYER li1 ;
        RECT 3380.500 3629.765 3380.670 3629.805 ;
        RECT 3380.500 3629.515 3381.150 3629.765 ;
        RECT 3380.670 3629.435 3381.150 3629.515 ;
        RECT 3380.500 3629.055 3380.670 3629.345 ;
      LAYER li1 ;
        RECT 3381.320 3629.265 3381.490 3629.935 ;
        RECT 3380.840 3629.095 3381.490 3629.265 ;
      LAYER li1 ;
        RECT 3380.670 3628.885 3381.150 3628.925 ;
        RECT 3380.500 3628.595 3381.150 3628.885 ;
      LAYER li1 ;
        RECT 3381.320 3628.425 3381.490 3629.095 ;
      LAYER li1 ;
        RECT 3380.500 3628.135 3380.670 3628.425 ;
      LAYER li1 ;
        RECT 3380.840 3628.255 3381.490 3628.425 ;
      LAYER li1 ;
        RECT 3380.670 3627.965 3381.150 3628.085 ;
        RECT 3380.500 3627.755 3381.150 3627.965 ;
        RECT 3380.500 3627.675 3380.670 3627.755 ;
      LAYER li1 ;
        RECT 3381.320 3627.670 3381.490 3628.255 ;
      LAYER li1 ;
        RECT 3381.660 3627.915 3381.830 3630.365 ;
        RECT 3382.420 3630.355 3383.220 3630.435 ;
        RECT 3383.390 3630.315 3384.190 3630.435 ;
      LAYER li1 ;
        RECT 3382.030 3629.935 3383.050 3630.105 ;
      LAYER li1 ;
        RECT 3383.220 3629.975 3383.390 3630.265 ;
      LAYER li1 ;
        RECT 3384.410 3630.145 3384.580 3630.730 ;
        RECT 3383.560 3629.975 3384.580 3630.145 ;
        RECT 3382.030 3629.265 3382.200 3629.935 ;
      LAYER li1 ;
        RECT 3383.220 3629.765 3384.190 3629.805 ;
        RECT 3382.420 3629.515 3384.190 3629.765 ;
        RECT 3382.420 3629.435 3383.220 3629.515 ;
        RECT 3383.390 3629.475 3384.190 3629.515 ;
      LAYER li1 ;
        RECT 3382.030 3629.095 3383.050 3629.265 ;
        RECT 3382.030 3628.425 3382.200 3629.095 ;
      LAYER li1 ;
        RECT 3383.220 3629.055 3383.390 3629.345 ;
      LAYER li1 ;
        RECT 3384.410 3629.305 3384.580 3629.975 ;
        RECT 3383.560 3629.135 3384.580 3629.305 ;
      LAYER li1 ;
        RECT 3382.420 3628.885 3383.220 3628.925 ;
        RECT 3383.390 3628.885 3384.190 3628.965 ;
        RECT 3382.420 3628.635 3384.190 3628.885 ;
        RECT 3382.420 3628.595 3383.390 3628.635 ;
      LAYER li1 ;
        RECT 3384.410 3628.465 3384.580 3629.135 ;
        RECT 3382.030 3628.255 3383.050 3628.425 ;
        RECT 3382.030 3627.670 3382.200 3628.255 ;
      LAYER li1 ;
        RECT 3383.220 3628.135 3383.390 3628.425 ;
      LAYER li1 ;
        RECT 3383.560 3628.295 3384.580 3628.465 ;
      LAYER li1 ;
        RECT 3382.420 3627.965 3383.220 3628.085 ;
        RECT 3383.390 3627.965 3384.190 3628.045 ;
        RECT 3384.780 3628.035 3384.950 3630.485 ;
      LAYER li1 ;
        RECT 3385.120 3630.145 3385.290 3630.730 ;
      LAYER li1 ;
        RECT 3385.940 3630.645 3386.110 3630.725 ;
        RECT 3385.460 3630.435 3386.110 3630.645 ;
        RECT 3385.460 3630.315 3385.940 3630.435 ;
      LAYER li1 ;
        RECT 3385.120 3629.975 3385.770 3630.145 ;
      LAYER li1 ;
        RECT 3385.940 3629.975 3386.110 3630.265 ;
      LAYER li1 ;
        RECT 3385.120 3629.305 3385.290 3629.975 ;
      LAYER li1 ;
        RECT 3385.460 3629.515 3386.110 3629.805 ;
        RECT 3385.460 3629.475 3385.940 3629.515 ;
      LAYER li1 ;
        RECT 3385.120 3629.135 3385.770 3629.305 ;
        RECT 3385.120 3628.465 3385.290 3629.135 ;
      LAYER li1 ;
        RECT 3385.940 3629.055 3386.110 3629.345 ;
        RECT 3385.460 3628.885 3385.940 3628.965 ;
        RECT 3385.460 3628.635 3386.110 3628.885 ;
        RECT 3385.940 3628.595 3386.110 3628.635 ;
      LAYER li1 ;
        RECT 3385.120 3628.295 3385.770 3628.465 ;
      LAYER li1 ;
        RECT 3385.940 3628.135 3386.110 3628.425 ;
        RECT 3382.420 3627.875 3384.190 3627.965 ;
        RECT 3382.420 3627.755 3383.390 3627.875 ;
        RECT 3383.220 3627.675 3383.390 3627.755 ;
        RECT 3384.410 3627.860 3385.290 3628.035 ;
        RECT 3384.410 3627.705 3384.580 3627.860 ;
      LAYER li1 ;
        RECT 3381.320 3627.585 3382.200 3627.670 ;
      LAYER li1 ;
        RECT 3380.500 3627.245 3380.670 3627.505 ;
      LAYER li1 ;
        RECT 3380.840 3627.415 3383.050 3627.585 ;
      LAYER li1 ;
        RECT 3383.220 3627.245 3383.390 3627.505 ;
        RECT 3383.560 3627.375 3384.580 3627.705 ;
        RECT 3380.500 3627.215 3381.470 3627.245 ;
        RECT 3380.670 3627.045 3381.470 3627.215 ;
        RECT 3380.500 3626.915 3381.470 3627.045 ;
        RECT 3382.070 3627.215 3383.390 3627.245 ;
        RECT 3382.070 3627.045 3383.220 3627.215 ;
        RECT 3383.390 3627.045 3384.190 3627.205 ;
        RECT 3382.070 3627.035 3384.190 3627.045 ;
        RECT 3382.070 3626.915 3383.390 3627.035 ;
        RECT 3380.500 3626.755 3380.670 3626.915 ;
        RECT 3383.220 3626.755 3383.390 3626.915 ;
        RECT 3384.410 3626.865 3384.580 3627.375 ;
        RECT 3377.780 3626.355 3377.950 3626.440 ;
        RECT 3380.500 3626.355 3380.670 3626.585 ;
        RECT 3383.220 3626.355 3383.390 3626.585 ;
        RECT 3383.560 3626.535 3384.580 3626.865 ;
      LAYER li1 ;
        RECT 3384.750 3626.580 3384.950 3627.680 ;
      LAYER li1 ;
        RECT 3385.120 3627.625 3385.290 3627.860 ;
        RECT 3385.460 3627.965 3385.940 3628.125 ;
        RECT 3385.460 3627.795 3386.110 3627.965 ;
        RECT 3385.940 3627.675 3386.110 3627.795 ;
        RECT 3385.120 3627.455 3385.765 3627.625 ;
        RECT 3385.120 3626.785 3385.290 3627.455 ;
        RECT 3385.940 3627.285 3386.110 3627.505 ;
        RECT 3385.460 3627.215 3386.110 3627.285 ;
        RECT 3385.460 3627.045 3385.940 3627.215 ;
        RECT 3385.460 3626.955 3386.110 3627.045 ;
        RECT 3385.120 3626.615 3385.770 3626.785 ;
        RECT 3385.940 3626.755 3386.110 3626.955 ;
        RECT 3385.940 3626.355 3386.110 3626.585 ;
        RECT 3377.780 3626.295 3379.115 3626.355 ;
        RECT 3377.950 3626.125 3379.115 3626.295 ;
        RECT 3377.780 3626.065 3379.115 3626.125 ;
        RECT 3379.775 3626.295 3381.395 3626.355 ;
        RECT 3379.775 3626.125 3380.500 3626.295 ;
        RECT 3380.670 3626.125 3381.395 3626.295 ;
        RECT 3379.775 3626.065 3381.395 3626.125 ;
        RECT 3377.780 3625.980 3377.950 3626.065 ;
      LAYER li1 ;
        RECT 3379.955 3624.310 3380.500 3625.895 ;
      LAYER li1 ;
        RECT 3380.500 3625.835 3380.670 3626.065 ;
        RECT 3380.500 3625.465 3380.670 3625.665 ;
        RECT 3380.840 3625.635 3381.490 3625.805 ;
        RECT 3380.500 3625.375 3381.150 3625.465 ;
        RECT 3380.670 3625.205 3381.150 3625.375 ;
        RECT 3380.500 3625.135 3381.150 3625.205 ;
        RECT 3380.500 3624.915 3380.670 3625.135 ;
        RECT 3381.320 3624.965 3381.490 3625.635 ;
        RECT 3380.845 3624.795 3381.490 3624.965 ;
        RECT 3380.500 3624.625 3380.670 3624.745 ;
        RECT 3380.500 3624.455 3381.150 3624.625 ;
      LAYER li1 ;
        RECT 3379.125 3623.970 3380.500 3624.310 ;
      LAYER li1 ;
        RECT 3380.670 3624.295 3381.150 3624.455 ;
        RECT 3381.320 3624.560 3381.490 3624.795 ;
      LAYER li1 ;
        RECT 3381.660 3624.740 3381.860 3626.330 ;
      LAYER li1 ;
        RECT 3382.055 3626.295 3384.555 3626.355 ;
        RECT 3382.055 3626.125 3383.220 3626.295 ;
        RECT 3383.390 3626.125 3384.555 3626.295 ;
        RECT 3382.055 3626.065 3384.555 3626.125 ;
        RECT 3385.215 3626.295 3386.110 3626.355 ;
        RECT 3385.215 3626.125 3385.940 3626.295 ;
        RECT 3385.215 3626.065 3386.110 3626.125 ;
        RECT 3382.030 3625.555 3383.050 3625.885 ;
        RECT 3383.220 3625.835 3383.390 3626.065 ;
        RECT 3385.940 3625.835 3386.110 3626.065 ;
        RECT 3382.030 3625.045 3382.200 3625.555 ;
        RECT 3383.220 3625.505 3383.390 3625.665 ;
        RECT 3385.940 3625.505 3386.110 3625.665 ;
        RECT 3383.220 3625.385 3384.540 3625.505 ;
        RECT 3382.420 3625.375 3384.540 3625.385 ;
        RECT 3382.420 3625.215 3383.220 3625.375 ;
        RECT 3383.390 3625.205 3384.540 3625.375 ;
        RECT 3383.220 3625.175 3384.540 3625.205 ;
        RECT 3385.140 3625.375 3386.110 3625.505 ;
        RECT 3385.140 3625.205 3385.940 3625.375 ;
        RECT 3385.140 3625.175 3386.110 3625.205 ;
        RECT 3382.030 3624.715 3383.050 3625.045 ;
        RECT 3383.220 3624.915 3383.390 3625.175 ;
      LAYER li1 ;
        RECT 3383.560 3624.835 3385.770 3625.005 ;
      LAYER li1 ;
        RECT 3385.940 3624.915 3386.110 3625.175 ;
      LAYER li1 ;
        RECT 3384.410 3624.750 3385.290 3624.835 ;
      LAYER li1 ;
        RECT 3382.030 3624.560 3382.200 3624.715 ;
        RECT 3381.320 3624.385 3382.200 3624.560 ;
        RECT 3383.220 3624.665 3383.390 3624.745 ;
        RECT 3383.220 3624.545 3384.190 3624.665 ;
        RECT 3382.420 3624.455 3384.190 3624.545 ;
        RECT 3380.500 3623.995 3380.670 3624.285 ;
      LAYER li1 ;
        RECT 3379.955 3620.550 3380.500 3623.970 ;
        RECT 3380.840 3623.955 3381.490 3624.125 ;
      LAYER li1 ;
        RECT 3380.500 3623.785 3380.670 3623.825 ;
        RECT 3380.500 3623.535 3381.150 3623.785 ;
        RECT 3380.670 3623.455 3381.150 3623.535 ;
        RECT 3380.500 3623.075 3380.670 3623.365 ;
      LAYER li1 ;
        RECT 3381.320 3623.285 3381.490 3623.955 ;
        RECT 3380.840 3623.115 3381.490 3623.285 ;
      LAYER li1 ;
        RECT 3380.670 3622.905 3381.150 3622.945 ;
        RECT 3380.500 3622.615 3381.150 3622.905 ;
      LAYER li1 ;
        RECT 3381.320 3622.445 3381.490 3623.115 ;
      LAYER li1 ;
        RECT 3380.500 3622.155 3380.670 3622.445 ;
      LAYER li1 ;
        RECT 3380.840 3622.275 3381.490 3622.445 ;
      LAYER li1 ;
        RECT 3380.670 3621.985 3381.150 3622.105 ;
        RECT 3380.500 3621.775 3381.150 3621.985 ;
        RECT 3380.500 3621.695 3380.670 3621.775 ;
      LAYER li1 ;
        RECT 3381.320 3621.690 3381.490 3622.275 ;
      LAYER li1 ;
        RECT 3381.660 3621.935 3381.830 3624.385 ;
        RECT 3382.420 3624.375 3383.220 3624.455 ;
        RECT 3383.390 3624.335 3384.190 3624.455 ;
      LAYER li1 ;
        RECT 3382.030 3623.955 3383.050 3624.125 ;
      LAYER li1 ;
        RECT 3383.220 3623.995 3383.390 3624.285 ;
      LAYER li1 ;
        RECT 3384.410 3624.165 3384.580 3624.750 ;
        RECT 3383.560 3623.995 3384.580 3624.165 ;
        RECT 3382.030 3623.285 3382.200 3623.955 ;
      LAYER li1 ;
        RECT 3383.220 3623.785 3384.190 3623.825 ;
        RECT 3382.420 3623.535 3384.190 3623.785 ;
        RECT 3382.420 3623.455 3383.220 3623.535 ;
        RECT 3383.390 3623.495 3384.190 3623.535 ;
      LAYER li1 ;
        RECT 3382.030 3623.115 3383.050 3623.285 ;
        RECT 3382.030 3622.445 3382.200 3623.115 ;
      LAYER li1 ;
        RECT 3383.220 3623.075 3383.390 3623.365 ;
      LAYER li1 ;
        RECT 3384.410 3623.325 3384.580 3623.995 ;
        RECT 3383.560 3623.155 3384.580 3623.325 ;
      LAYER li1 ;
        RECT 3382.420 3622.905 3383.220 3622.945 ;
        RECT 3383.390 3622.905 3384.190 3622.985 ;
        RECT 3382.420 3622.655 3384.190 3622.905 ;
        RECT 3382.420 3622.615 3383.390 3622.655 ;
      LAYER li1 ;
        RECT 3384.410 3622.485 3384.580 3623.155 ;
        RECT 3382.030 3622.275 3383.050 3622.445 ;
        RECT 3382.030 3621.690 3382.200 3622.275 ;
      LAYER li1 ;
        RECT 3383.220 3622.155 3383.390 3622.445 ;
      LAYER li1 ;
        RECT 3383.560 3622.315 3384.580 3622.485 ;
      LAYER li1 ;
        RECT 3382.420 3621.985 3383.220 3622.105 ;
        RECT 3383.390 3621.985 3384.190 3622.065 ;
        RECT 3384.780 3622.055 3384.950 3624.505 ;
      LAYER li1 ;
        RECT 3385.120 3624.165 3385.290 3624.750 ;
      LAYER li1 ;
        RECT 3385.940 3624.665 3386.110 3624.745 ;
        RECT 3385.460 3624.455 3386.110 3624.665 ;
        RECT 3385.460 3624.335 3385.940 3624.455 ;
      LAYER li1 ;
        RECT 3385.120 3623.995 3385.770 3624.165 ;
      LAYER li1 ;
        RECT 3385.940 3623.995 3386.110 3624.285 ;
      LAYER li1 ;
        RECT 3385.120 3623.325 3385.290 3623.995 ;
      LAYER li1 ;
        RECT 3385.460 3623.535 3386.110 3623.825 ;
        RECT 3385.460 3623.495 3385.940 3623.535 ;
      LAYER li1 ;
        RECT 3385.120 3623.155 3385.770 3623.325 ;
        RECT 3385.120 3622.485 3385.290 3623.155 ;
      LAYER li1 ;
        RECT 3385.940 3623.075 3386.110 3623.365 ;
        RECT 3385.460 3622.905 3385.940 3622.985 ;
        RECT 3385.460 3622.655 3386.110 3622.905 ;
        RECT 3385.940 3622.615 3386.110 3622.655 ;
      LAYER li1 ;
        RECT 3385.120 3622.315 3385.770 3622.485 ;
      LAYER li1 ;
        RECT 3385.940 3622.155 3386.110 3622.445 ;
        RECT 3382.420 3621.895 3384.190 3621.985 ;
        RECT 3382.420 3621.775 3383.390 3621.895 ;
        RECT 3383.220 3621.695 3383.390 3621.775 ;
        RECT 3384.410 3621.880 3385.290 3622.055 ;
        RECT 3384.410 3621.725 3384.580 3621.880 ;
      LAYER li1 ;
        RECT 3381.320 3621.605 3382.200 3621.690 ;
      LAYER li1 ;
        RECT 3380.500 3621.265 3380.670 3621.525 ;
      LAYER li1 ;
        RECT 3380.840 3621.435 3383.050 3621.605 ;
      LAYER li1 ;
        RECT 3383.220 3621.265 3383.390 3621.525 ;
        RECT 3383.560 3621.395 3384.580 3621.725 ;
        RECT 3380.500 3621.235 3381.470 3621.265 ;
        RECT 3380.670 3621.065 3381.470 3621.235 ;
        RECT 3380.500 3620.935 3381.470 3621.065 ;
        RECT 3382.070 3621.235 3383.390 3621.265 ;
        RECT 3382.070 3621.065 3383.220 3621.235 ;
        RECT 3383.390 3621.065 3384.190 3621.225 ;
        RECT 3382.070 3621.055 3384.190 3621.065 ;
        RECT 3382.070 3620.935 3383.390 3621.055 ;
        RECT 3380.500 3620.775 3380.670 3620.935 ;
        RECT 3383.220 3620.775 3383.390 3620.935 ;
        RECT 3384.410 3620.885 3384.580 3621.395 ;
        RECT 3377.780 3620.375 3377.950 3620.460 ;
        RECT 3380.500 3620.375 3380.670 3620.605 ;
        RECT 3383.220 3620.375 3383.390 3620.605 ;
        RECT 3383.560 3620.555 3384.580 3620.885 ;
      LAYER li1 ;
        RECT 3384.750 3620.600 3384.950 3621.700 ;
      LAYER li1 ;
        RECT 3385.120 3621.645 3385.290 3621.880 ;
        RECT 3385.460 3621.985 3385.940 3622.145 ;
        RECT 3385.460 3621.815 3386.110 3621.985 ;
        RECT 3385.940 3621.695 3386.110 3621.815 ;
        RECT 3385.120 3621.475 3385.765 3621.645 ;
        RECT 3385.120 3620.805 3385.290 3621.475 ;
        RECT 3385.940 3621.305 3386.110 3621.525 ;
        RECT 3385.460 3621.235 3386.110 3621.305 ;
        RECT 3385.460 3621.065 3385.940 3621.235 ;
        RECT 3385.460 3620.975 3386.110 3621.065 ;
        RECT 3385.120 3620.635 3385.770 3620.805 ;
        RECT 3385.940 3620.775 3386.110 3620.975 ;
        RECT 3385.940 3620.375 3386.110 3620.605 ;
        RECT 3377.780 3620.315 3379.115 3620.375 ;
        RECT 3377.950 3620.145 3379.115 3620.315 ;
        RECT 3377.780 3620.085 3379.115 3620.145 ;
        RECT 3379.775 3620.315 3381.395 3620.375 ;
        RECT 3379.775 3620.145 3380.500 3620.315 ;
        RECT 3380.670 3620.145 3381.395 3620.315 ;
        RECT 3379.775 3620.085 3381.395 3620.145 ;
        RECT 3377.780 3620.000 3377.950 3620.085 ;
      LAYER li1 ;
        RECT 3379.955 3618.330 3380.500 3619.915 ;
      LAYER li1 ;
        RECT 3380.500 3619.855 3380.670 3620.085 ;
        RECT 3380.500 3619.485 3380.670 3619.685 ;
        RECT 3380.840 3619.655 3381.490 3619.825 ;
        RECT 3380.500 3619.395 3381.150 3619.485 ;
        RECT 3380.670 3619.225 3381.150 3619.395 ;
        RECT 3380.500 3619.155 3381.150 3619.225 ;
        RECT 3380.500 3618.935 3380.670 3619.155 ;
        RECT 3381.320 3618.985 3381.490 3619.655 ;
        RECT 3380.845 3618.815 3381.490 3618.985 ;
        RECT 3380.500 3618.645 3380.670 3618.765 ;
        RECT 3380.500 3618.475 3381.150 3618.645 ;
      LAYER li1 ;
        RECT 3379.125 3617.990 3380.500 3618.330 ;
      LAYER li1 ;
        RECT 3380.670 3618.315 3381.150 3618.475 ;
        RECT 3381.320 3618.580 3381.490 3618.815 ;
      LAYER li1 ;
        RECT 3381.660 3618.760 3381.860 3620.350 ;
      LAYER li1 ;
        RECT 3382.055 3620.315 3384.555 3620.375 ;
        RECT 3382.055 3620.145 3383.220 3620.315 ;
        RECT 3383.390 3620.145 3384.555 3620.315 ;
        RECT 3382.055 3620.085 3384.555 3620.145 ;
        RECT 3385.215 3620.315 3386.110 3620.375 ;
        RECT 3385.215 3620.145 3385.940 3620.315 ;
        RECT 3385.215 3620.085 3386.110 3620.145 ;
        RECT 3382.030 3619.575 3383.050 3619.905 ;
        RECT 3383.220 3619.855 3383.390 3620.085 ;
        RECT 3385.940 3619.855 3386.110 3620.085 ;
        RECT 3382.030 3619.065 3382.200 3619.575 ;
        RECT 3383.220 3619.525 3383.390 3619.685 ;
        RECT 3385.940 3619.525 3386.110 3619.685 ;
        RECT 3383.220 3619.405 3384.540 3619.525 ;
        RECT 3382.420 3619.395 3384.540 3619.405 ;
        RECT 3382.420 3619.235 3383.220 3619.395 ;
        RECT 3383.390 3619.225 3384.540 3619.395 ;
        RECT 3383.220 3619.195 3384.540 3619.225 ;
        RECT 3385.140 3619.395 3386.110 3619.525 ;
        RECT 3385.140 3619.225 3385.940 3619.395 ;
        RECT 3385.140 3619.195 3386.110 3619.225 ;
        RECT 3382.030 3618.735 3383.050 3619.065 ;
        RECT 3383.220 3618.935 3383.390 3619.195 ;
      LAYER li1 ;
        RECT 3383.560 3618.855 3385.770 3619.025 ;
      LAYER li1 ;
        RECT 3385.940 3618.935 3386.110 3619.195 ;
      LAYER li1 ;
        RECT 3384.410 3618.770 3385.290 3618.855 ;
      LAYER li1 ;
        RECT 3382.030 3618.580 3382.200 3618.735 ;
        RECT 3381.320 3618.405 3382.200 3618.580 ;
        RECT 3383.220 3618.685 3383.390 3618.765 ;
        RECT 3383.220 3618.565 3384.190 3618.685 ;
        RECT 3382.420 3618.475 3384.190 3618.565 ;
        RECT 3380.500 3618.015 3380.670 3618.305 ;
      LAYER li1 ;
        RECT 3379.955 3614.570 3380.500 3617.990 ;
        RECT 3380.840 3617.975 3381.490 3618.145 ;
      LAYER li1 ;
        RECT 3380.500 3617.805 3380.670 3617.845 ;
        RECT 3380.500 3617.555 3381.150 3617.805 ;
        RECT 3380.670 3617.475 3381.150 3617.555 ;
        RECT 3380.500 3617.095 3380.670 3617.385 ;
      LAYER li1 ;
        RECT 3381.320 3617.305 3381.490 3617.975 ;
        RECT 3380.840 3617.135 3381.490 3617.305 ;
      LAYER li1 ;
        RECT 3380.670 3616.925 3381.150 3616.965 ;
        RECT 3380.500 3616.635 3381.150 3616.925 ;
      LAYER li1 ;
        RECT 3381.320 3616.465 3381.490 3617.135 ;
      LAYER li1 ;
        RECT 3380.500 3616.175 3380.670 3616.465 ;
      LAYER li1 ;
        RECT 3380.840 3616.295 3381.490 3616.465 ;
      LAYER li1 ;
        RECT 3380.670 3616.005 3381.150 3616.125 ;
        RECT 3380.500 3615.795 3381.150 3616.005 ;
        RECT 3380.500 3615.715 3380.670 3615.795 ;
      LAYER li1 ;
        RECT 3381.320 3615.710 3381.490 3616.295 ;
      LAYER li1 ;
        RECT 3381.660 3615.955 3381.830 3618.405 ;
        RECT 3382.420 3618.395 3383.220 3618.475 ;
        RECT 3383.390 3618.355 3384.190 3618.475 ;
      LAYER li1 ;
        RECT 3382.030 3617.975 3383.050 3618.145 ;
      LAYER li1 ;
        RECT 3383.220 3618.015 3383.390 3618.305 ;
      LAYER li1 ;
        RECT 3384.410 3618.185 3384.580 3618.770 ;
        RECT 3383.560 3618.015 3384.580 3618.185 ;
        RECT 3382.030 3617.305 3382.200 3617.975 ;
      LAYER li1 ;
        RECT 3383.220 3617.805 3384.190 3617.845 ;
        RECT 3382.420 3617.555 3384.190 3617.805 ;
        RECT 3382.420 3617.475 3383.220 3617.555 ;
        RECT 3383.390 3617.515 3384.190 3617.555 ;
      LAYER li1 ;
        RECT 3382.030 3617.135 3383.050 3617.305 ;
        RECT 3382.030 3616.465 3382.200 3617.135 ;
      LAYER li1 ;
        RECT 3383.220 3617.095 3383.390 3617.385 ;
      LAYER li1 ;
        RECT 3384.410 3617.345 3384.580 3618.015 ;
        RECT 3383.560 3617.175 3384.580 3617.345 ;
      LAYER li1 ;
        RECT 3382.420 3616.925 3383.220 3616.965 ;
        RECT 3383.390 3616.925 3384.190 3617.005 ;
        RECT 3382.420 3616.675 3384.190 3616.925 ;
        RECT 3382.420 3616.635 3383.390 3616.675 ;
      LAYER li1 ;
        RECT 3384.410 3616.505 3384.580 3617.175 ;
        RECT 3382.030 3616.295 3383.050 3616.465 ;
        RECT 3382.030 3615.710 3382.200 3616.295 ;
      LAYER li1 ;
        RECT 3383.220 3616.175 3383.390 3616.465 ;
      LAYER li1 ;
        RECT 3383.560 3616.335 3384.580 3616.505 ;
      LAYER li1 ;
        RECT 3382.420 3616.005 3383.220 3616.125 ;
        RECT 3383.390 3616.005 3384.190 3616.085 ;
        RECT 3384.780 3616.075 3384.950 3618.525 ;
      LAYER li1 ;
        RECT 3385.120 3618.185 3385.290 3618.770 ;
      LAYER li1 ;
        RECT 3385.940 3618.685 3386.110 3618.765 ;
        RECT 3385.460 3618.475 3386.110 3618.685 ;
        RECT 3385.460 3618.355 3385.940 3618.475 ;
      LAYER li1 ;
        RECT 3385.120 3618.015 3385.770 3618.185 ;
      LAYER li1 ;
        RECT 3385.940 3618.015 3386.110 3618.305 ;
      LAYER li1 ;
        RECT 3385.120 3617.345 3385.290 3618.015 ;
      LAYER li1 ;
        RECT 3385.460 3617.555 3386.110 3617.845 ;
        RECT 3385.460 3617.515 3385.940 3617.555 ;
      LAYER li1 ;
        RECT 3385.120 3617.175 3385.770 3617.345 ;
        RECT 3385.120 3616.505 3385.290 3617.175 ;
      LAYER li1 ;
        RECT 3385.940 3617.095 3386.110 3617.385 ;
        RECT 3385.460 3616.925 3385.940 3617.005 ;
        RECT 3385.460 3616.675 3386.110 3616.925 ;
        RECT 3385.940 3616.635 3386.110 3616.675 ;
      LAYER li1 ;
        RECT 3385.120 3616.335 3385.770 3616.505 ;
      LAYER li1 ;
        RECT 3385.940 3616.175 3386.110 3616.465 ;
        RECT 3382.420 3615.915 3384.190 3616.005 ;
        RECT 3382.420 3615.795 3383.390 3615.915 ;
        RECT 3383.220 3615.715 3383.390 3615.795 ;
        RECT 3384.410 3615.900 3385.290 3616.075 ;
        RECT 3384.410 3615.745 3384.580 3615.900 ;
      LAYER li1 ;
        RECT 3381.320 3615.625 3382.200 3615.710 ;
      LAYER li1 ;
        RECT 3380.500 3615.285 3380.670 3615.545 ;
      LAYER li1 ;
        RECT 3380.840 3615.455 3383.050 3615.625 ;
      LAYER li1 ;
        RECT 3383.220 3615.285 3383.390 3615.545 ;
        RECT 3383.560 3615.415 3384.580 3615.745 ;
        RECT 3380.500 3615.255 3381.470 3615.285 ;
        RECT 3380.670 3615.085 3381.470 3615.255 ;
        RECT 3380.500 3614.955 3381.470 3615.085 ;
        RECT 3382.070 3615.255 3383.390 3615.285 ;
        RECT 3382.070 3615.085 3383.220 3615.255 ;
        RECT 3383.390 3615.085 3384.190 3615.245 ;
        RECT 3382.070 3615.075 3384.190 3615.085 ;
        RECT 3382.070 3614.955 3383.390 3615.075 ;
        RECT 3380.500 3614.795 3380.670 3614.955 ;
        RECT 3383.220 3614.795 3383.390 3614.955 ;
        RECT 3384.410 3614.905 3384.580 3615.415 ;
        RECT 3377.780 3614.395 3377.950 3614.480 ;
        RECT 3380.500 3614.395 3380.670 3614.625 ;
        RECT 3383.220 3614.395 3383.390 3614.625 ;
        RECT 3383.560 3614.575 3384.580 3614.905 ;
      LAYER li1 ;
        RECT 3384.750 3614.620 3384.950 3615.720 ;
      LAYER li1 ;
        RECT 3385.120 3615.665 3385.290 3615.900 ;
        RECT 3385.460 3616.005 3385.940 3616.165 ;
        RECT 3385.460 3615.835 3386.110 3616.005 ;
        RECT 3385.940 3615.715 3386.110 3615.835 ;
        RECT 3385.120 3615.495 3385.765 3615.665 ;
        RECT 3385.120 3614.825 3385.290 3615.495 ;
        RECT 3385.940 3615.325 3386.110 3615.545 ;
        RECT 3385.460 3615.255 3386.110 3615.325 ;
        RECT 3385.460 3615.085 3385.940 3615.255 ;
        RECT 3385.460 3614.995 3386.110 3615.085 ;
        RECT 3385.120 3614.655 3385.770 3614.825 ;
        RECT 3385.940 3614.795 3386.110 3614.995 ;
        RECT 3385.940 3614.395 3386.110 3614.625 ;
        RECT 3377.780 3614.335 3379.115 3614.395 ;
        RECT 3377.950 3614.165 3379.115 3614.335 ;
        RECT 3377.780 3614.105 3379.115 3614.165 ;
        RECT 3379.775 3614.335 3381.395 3614.395 ;
        RECT 3379.775 3614.165 3380.500 3614.335 ;
        RECT 3380.670 3614.165 3381.395 3614.335 ;
        RECT 3379.775 3614.105 3381.395 3614.165 ;
        RECT 3382.055 3614.335 3384.555 3614.395 ;
        RECT 3382.055 3614.165 3383.220 3614.335 ;
        RECT 3383.390 3614.165 3384.555 3614.335 ;
        RECT 3382.055 3614.105 3384.555 3614.165 ;
        RECT 3385.215 3614.335 3386.110 3614.395 ;
        RECT 3385.215 3614.165 3385.940 3614.335 ;
        RECT 3385.215 3614.105 3386.110 3614.165 ;
        RECT 3377.780 3614.020 3377.950 3614.105 ;
      LAYER li1 ;
        RECT 3379.955 3612.350 3380.500 3613.935 ;
      LAYER li1 ;
        RECT 3380.500 3613.875 3380.670 3614.105 ;
        RECT 3380.500 3613.505 3380.670 3613.705 ;
        RECT 3380.840 3613.675 3381.490 3613.845 ;
        RECT 3380.500 3613.415 3381.150 3613.505 ;
        RECT 3380.670 3613.245 3381.150 3613.415 ;
        RECT 3380.500 3613.175 3381.150 3613.245 ;
        RECT 3380.500 3612.955 3380.670 3613.175 ;
        RECT 3381.320 3613.005 3381.490 3613.675 ;
        RECT 3380.845 3612.835 3381.490 3613.005 ;
        RECT 3380.500 3612.665 3380.670 3612.785 ;
        RECT 3380.500 3612.495 3381.150 3612.665 ;
      LAYER li1 ;
        RECT 3379.125 3612.010 3380.500 3612.350 ;
      LAYER li1 ;
        RECT 3380.670 3612.335 3381.150 3612.495 ;
        RECT 3381.320 3612.600 3381.490 3612.835 ;
        RECT 3382.030 3613.595 3383.050 3613.925 ;
        RECT 3383.220 3613.875 3383.390 3614.105 ;
        RECT 3385.940 3613.875 3386.110 3614.105 ;
        RECT 3382.030 3613.085 3382.200 3613.595 ;
        RECT 3383.220 3613.545 3383.390 3613.705 ;
        RECT 3385.940 3613.545 3386.110 3613.705 ;
        RECT 3383.220 3613.425 3384.540 3613.545 ;
        RECT 3382.420 3613.415 3384.540 3613.425 ;
        RECT 3382.420 3613.255 3383.220 3613.415 ;
        RECT 3383.390 3613.245 3384.540 3613.415 ;
        RECT 3383.220 3613.215 3384.540 3613.245 ;
        RECT 3385.140 3613.415 3386.110 3613.545 ;
        RECT 3385.140 3613.245 3385.940 3613.415 ;
        RECT 3385.140 3613.215 3386.110 3613.245 ;
        RECT 3382.030 3612.755 3383.050 3613.085 ;
        RECT 3383.220 3612.955 3383.390 3613.215 ;
        RECT 3385.940 3612.955 3386.110 3613.215 ;
        RECT 3382.030 3612.600 3382.200 3612.755 ;
        RECT 3381.320 3612.425 3382.200 3612.600 ;
        RECT 3383.220 3612.705 3383.390 3612.785 ;
        RECT 3385.940 3612.705 3386.110 3612.785 ;
        RECT 3383.220 3612.585 3384.190 3612.705 ;
        RECT 3382.420 3612.495 3384.190 3612.585 ;
        RECT 3380.500 3612.035 3380.670 3612.325 ;
      LAYER li1 ;
        RECT 3379.955 3608.590 3380.500 3612.010 ;
        RECT 3380.840 3611.995 3381.490 3612.165 ;
      LAYER li1 ;
        RECT 3380.500 3611.825 3380.670 3611.865 ;
        RECT 3380.500 3611.575 3381.150 3611.825 ;
        RECT 3380.670 3611.495 3381.150 3611.575 ;
        RECT 3380.500 3611.115 3380.670 3611.405 ;
      LAYER li1 ;
        RECT 3381.320 3611.325 3381.490 3611.995 ;
        RECT 3380.840 3611.155 3381.490 3611.325 ;
      LAYER li1 ;
        RECT 3380.670 3610.945 3381.150 3610.985 ;
        RECT 3380.500 3610.655 3381.150 3610.945 ;
      LAYER li1 ;
        RECT 3381.320 3610.485 3381.490 3611.155 ;
      LAYER li1 ;
        RECT 3380.500 3610.195 3380.670 3610.485 ;
      LAYER li1 ;
        RECT 3380.840 3610.315 3381.490 3610.485 ;
      LAYER li1 ;
        RECT 3380.670 3610.025 3381.150 3610.145 ;
        RECT 3380.500 3609.815 3381.150 3610.025 ;
        RECT 3380.500 3609.735 3380.670 3609.815 ;
      LAYER li1 ;
        RECT 3381.320 3609.730 3381.490 3610.315 ;
      LAYER li1 ;
        RECT 3381.660 3609.975 3381.830 3612.425 ;
        RECT 3382.420 3612.415 3383.220 3612.495 ;
        RECT 3383.390 3612.375 3384.190 3612.495 ;
      LAYER li1 ;
        RECT 3382.030 3611.995 3383.050 3612.165 ;
      LAYER li1 ;
        RECT 3383.220 3612.035 3383.390 3612.325 ;
      LAYER li1 ;
        RECT 3382.030 3611.325 3382.200 3611.995 ;
      LAYER li1 ;
        RECT 3383.220 3611.825 3384.190 3611.865 ;
        RECT 3382.420 3611.575 3384.190 3611.825 ;
        RECT 3382.420 3611.495 3383.220 3611.575 ;
        RECT 3383.390 3611.535 3384.190 3611.575 ;
      LAYER li1 ;
        RECT 3382.030 3611.155 3383.050 3611.325 ;
        RECT 3382.030 3610.485 3382.200 3611.155 ;
      LAYER li1 ;
        RECT 3383.220 3611.115 3383.390 3611.405 ;
        RECT 3382.420 3610.945 3383.220 3610.985 ;
        RECT 3383.390 3610.945 3384.190 3611.025 ;
        RECT 3382.420 3610.695 3384.190 3610.945 ;
        RECT 3382.420 3610.655 3383.390 3610.695 ;
      LAYER li1 ;
        RECT 3382.030 3610.315 3383.050 3610.485 ;
        RECT 3382.030 3609.730 3382.200 3610.315 ;
      LAYER li1 ;
        RECT 3383.220 3610.195 3383.390 3610.485 ;
        RECT 3382.420 3610.025 3383.220 3610.145 ;
        RECT 3383.390 3610.025 3384.190 3610.105 ;
        RECT 3384.780 3610.095 3384.950 3612.545 ;
        RECT 3385.460 3612.495 3386.110 3612.705 ;
        RECT 3385.460 3612.375 3385.940 3612.495 ;
        RECT 3385.940 3612.035 3386.110 3612.325 ;
        RECT 3385.460 3611.575 3386.110 3611.865 ;
        RECT 3385.460 3611.535 3385.940 3611.575 ;
        RECT 3385.940 3611.115 3386.110 3611.405 ;
        RECT 3385.460 3610.945 3385.940 3611.025 ;
        RECT 3385.460 3610.695 3386.110 3610.945 ;
        RECT 3385.940 3610.655 3386.110 3610.695 ;
        RECT 3385.940 3610.195 3386.110 3610.485 ;
        RECT 3382.420 3609.935 3384.190 3610.025 ;
        RECT 3382.420 3609.815 3383.390 3609.935 ;
        RECT 3383.220 3609.735 3383.390 3609.815 ;
        RECT 3384.410 3609.920 3385.290 3610.095 ;
        RECT 3384.410 3609.765 3384.580 3609.920 ;
      LAYER li1 ;
        RECT 3381.320 3609.645 3382.200 3609.730 ;
      LAYER li1 ;
        RECT 3380.500 3609.305 3380.670 3609.565 ;
      LAYER li1 ;
        RECT 3380.840 3609.475 3383.050 3609.645 ;
      LAYER li1 ;
        RECT 3383.220 3609.305 3383.390 3609.565 ;
        RECT 3383.560 3609.435 3384.580 3609.765 ;
        RECT 3380.500 3609.275 3381.470 3609.305 ;
        RECT 3380.670 3609.105 3381.470 3609.275 ;
        RECT 3380.500 3608.975 3381.470 3609.105 ;
        RECT 3382.070 3609.275 3383.390 3609.305 ;
        RECT 3382.070 3609.105 3383.220 3609.275 ;
        RECT 3383.390 3609.105 3384.190 3609.265 ;
        RECT 3382.070 3609.095 3384.190 3609.105 ;
        RECT 3382.070 3608.975 3383.390 3609.095 ;
        RECT 3380.500 3608.815 3380.670 3608.975 ;
        RECT 3383.220 3608.815 3383.390 3608.975 ;
        RECT 3384.410 3608.925 3384.580 3609.435 ;
        RECT 3377.780 3608.415 3377.950 3608.500 ;
        RECT 3380.500 3608.415 3380.670 3608.645 ;
        RECT 3383.220 3608.415 3383.390 3608.645 ;
        RECT 3383.560 3608.595 3384.580 3608.925 ;
      LAYER li1 ;
        RECT 3384.750 3608.640 3384.950 3609.740 ;
      LAYER li1 ;
        RECT 3385.120 3609.685 3385.290 3609.920 ;
        RECT 3385.460 3610.025 3385.940 3610.185 ;
        RECT 3385.460 3609.855 3386.110 3610.025 ;
        RECT 3385.940 3609.735 3386.110 3609.855 ;
        RECT 3385.120 3609.515 3385.765 3609.685 ;
        RECT 3385.120 3608.845 3385.290 3609.515 ;
        RECT 3385.940 3609.345 3386.110 3609.565 ;
        RECT 3385.460 3609.275 3386.110 3609.345 ;
        RECT 3385.460 3609.105 3385.940 3609.275 ;
        RECT 3385.460 3609.015 3386.110 3609.105 ;
        RECT 3385.120 3608.675 3385.770 3608.845 ;
        RECT 3385.940 3608.815 3386.110 3609.015 ;
        RECT 3385.940 3608.415 3386.110 3608.645 ;
        RECT 3377.780 3608.355 3379.115 3608.415 ;
        RECT 3377.950 3608.185 3379.115 3608.355 ;
        RECT 3377.780 3608.125 3379.115 3608.185 ;
        RECT 3379.775 3608.355 3381.395 3608.415 ;
        RECT 3379.775 3608.185 3380.500 3608.355 ;
        RECT 3380.670 3608.185 3381.395 3608.355 ;
        RECT 3379.775 3608.125 3381.395 3608.185 ;
        RECT 3382.055 3608.355 3384.555 3608.415 ;
        RECT 3382.055 3608.185 3383.220 3608.355 ;
        RECT 3383.390 3608.185 3384.555 3608.355 ;
        RECT 3382.055 3608.125 3384.555 3608.185 ;
        RECT 3385.215 3608.355 3386.110 3608.415 ;
        RECT 3385.215 3608.185 3385.940 3608.355 ;
        RECT 3385.215 3608.125 3386.110 3608.185 ;
        RECT 3377.780 3608.040 3377.950 3608.125 ;
      LAYER li1 ;
        RECT 3379.955 3606.370 3380.500 3607.955 ;
      LAYER li1 ;
        RECT 3380.500 3607.895 3380.670 3608.125 ;
        RECT 3380.500 3607.525 3380.670 3607.725 ;
        RECT 3380.840 3607.695 3381.490 3607.865 ;
        RECT 3380.500 3607.435 3381.150 3607.525 ;
        RECT 3380.670 3607.265 3381.150 3607.435 ;
        RECT 3380.500 3607.195 3381.150 3607.265 ;
        RECT 3380.500 3606.975 3380.670 3607.195 ;
        RECT 3381.320 3607.025 3381.490 3607.695 ;
        RECT 3380.845 3606.855 3381.490 3607.025 ;
        RECT 3380.500 3606.685 3380.670 3606.805 ;
        RECT 3380.500 3606.515 3381.150 3606.685 ;
      LAYER li1 ;
        RECT 3379.125 3606.030 3380.500 3606.370 ;
      LAYER li1 ;
        RECT 3380.670 3606.355 3381.150 3606.515 ;
        RECT 3381.320 3606.620 3381.490 3606.855 ;
        RECT 3382.030 3607.615 3383.050 3607.945 ;
        RECT 3383.220 3607.895 3383.390 3608.125 ;
        RECT 3385.940 3607.895 3386.110 3608.125 ;
        RECT 3382.030 3607.105 3382.200 3607.615 ;
        RECT 3383.220 3607.565 3383.390 3607.725 ;
        RECT 3385.940 3607.565 3386.110 3607.725 ;
        RECT 3383.220 3607.445 3384.540 3607.565 ;
        RECT 3382.420 3607.435 3384.540 3607.445 ;
        RECT 3382.420 3607.275 3383.220 3607.435 ;
        RECT 3383.390 3607.265 3384.540 3607.435 ;
        RECT 3383.220 3607.235 3384.540 3607.265 ;
        RECT 3385.140 3607.435 3386.110 3607.565 ;
        RECT 3385.140 3607.265 3385.940 3607.435 ;
        RECT 3385.140 3607.235 3386.110 3607.265 ;
        RECT 3382.030 3606.775 3383.050 3607.105 ;
        RECT 3383.220 3606.975 3383.390 3607.235 ;
        RECT 3385.940 3606.975 3386.110 3607.235 ;
        RECT 3382.030 3606.620 3382.200 3606.775 ;
        RECT 3381.320 3606.445 3382.200 3606.620 ;
        RECT 3383.220 3606.725 3383.390 3606.805 ;
        RECT 3385.940 3606.725 3386.110 3606.805 ;
        RECT 3383.220 3606.605 3384.190 3606.725 ;
        RECT 3382.420 3606.515 3384.190 3606.605 ;
        RECT 3380.500 3606.055 3380.670 3606.345 ;
      LAYER li1 ;
        RECT 3379.955 3602.610 3380.500 3606.030 ;
        RECT 3380.840 3606.015 3381.490 3606.185 ;
      LAYER li1 ;
        RECT 3380.500 3605.845 3380.670 3605.885 ;
        RECT 3380.500 3605.595 3381.150 3605.845 ;
        RECT 3380.670 3605.515 3381.150 3605.595 ;
        RECT 3380.500 3605.135 3380.670 3605.425 ;
      LAYER li1 ;
        RECT 3381.320 3605.345 3381.490 3606.015 ;
        RECT 3380.840 3605.175 3381.490 3605.345 ;
      LAYER li1 ;
        RECT 3380.670 3604.965 3381.150 3605.005 ;
        RECT 3380.500 3604.675 3381.150 3604.965 ;
      LAYER li1 ;
        RECT 3381.320 3604.505 3381.490 3605.175 ;
      LAYER li1 ;
        RECT 3380.500 3604.215 3380.670 3604.505 ;
      LAYER li1 ;
        RECT 3380.840 3604.335 3381.490 3604.505 ;
      LAYER li1 ;
        RECT 3380.670 3604.045 3381.150 3604.165 ;
        RECT 3380.500 3603.835 3381.150 3604.045 ;
        RECT 3380.500 3603.755 3380.670 3603.835 ;
      LAYER li1 ;
        RECT 3381.320 3603.750 3381.490 3604.335 ;
      LAYER li1 ;
        RECT 3381.660 3603.995 3381.830 3606.445 ;
        RECT 3382.420 3606.435 3383.220 3606.515 ;
        RECT 3383.390 3606.395 3384.190 3606.515 ;
      LAYER li1 ;
        RECT 3382.030 3606.015 3383.050 3606.185 ;
      LAYER li1 ;
        RECT 3383.220 3606.055 3383.390 3606.345 ;
      LAYER li1 ;
        RECT 3382.030 3605.345 3382.200 3606.015 ;
      LAYER li1 ;
        RECT 3383.220 3605.845 3384.190 3605.885 ;
        RECT 3382.420 3605.595 3384.190 3605.845 ;
        RECT 3382.420 3605.515 3383.220 3605.595 ;
        RECT 3383.390 3605.555 3384.190 3605.595 ;
      LAYER li1 ;
        RECT 3382.030 3605.175 3383.050 3605.345 ;
        RECT 3382.030 3604.505 3382.200 3605.175 ;
      LAYER li1 ;
        RECT 3383.220 3605.135 3383.390 3605.425 ;
        RECT 3382.420 3604.965 3383.220 3605.005 ;
        RECT 3383.390 3604.965 3384.190 3605.045 ;
        RECT 3382.420 3604.715 3384.190 3604.965 ;
        RECT 3382.420 3604.675 3383.390 3604.715 ;
      LAYER li1 ;
        RECT 3382.030 3604.335 3383.050 3604.505 ;
        RECT 3382.030 3603.750 3382.200 3604.335 ;
      LAYER li1 ;
        RECT 3383.220 3604.215 3383.390 3604.505 ;
        RECT 3382.420 3604.045 3383.220 3604.165 ;
        RECT 3383.390 3604.045 3384.190 3604.125 ;
        RECT 3384.780 3604.115 3384.950 3606.565 ;
        RECT 3385.460 3606.515 3386.110 3606.725 ;
        RECT 3385.460 3606.395 3385.940 3606.515 ;
        RECT 3385.940 3606.055 3386.110 3606.345 ;
        RECT 3385.460 3605.595 3386.110 3605.885 ;
        RECT 3385.460 3605.555 3385.940 3605.595 ;
        RECT 3385.940 3605.135 3386.110 3605.425 ;
        RECT 3385.460 3604.965 3385.940 3605.045 ;
        RECT 3385.460 3604.715 3386.110 3604.965 ;
        RECT 3385.940 3604.675 3386.110 3604.715 ;
        RECT 3385.940 3604.215 3386.110 3604.505 ;
        RECT 3382.420 3603.955 3384.190 3604.045 ;
        RECT 3382.420 3603.835 3383.390 3603.955 ;
        RECT 3383.220 3603.755 3383.390 3603.835 ;
        RECT 3384.410 3603.940 3385.290 3604.115 ;
        RECT 3384.410 3603.785 3384.580 3603.940 ;
      LAYER li1 ;
        RECT 3381.320 3603.665 3382.200 3603.750 ;
      LAYER li1 ;
        RECT 3380.500 3603.325 3380.670 3603.585 ;
      LAYER li1 ;
        RECT 3380.840 3603.495 3383.050 3603.665 ;
      LAYER li1 ;
        RECT 3383.220 3603.325 3383.390 3603.585 ;
        RECT 3383.560 3603.455 3384.580 3603.785 ;
        RECT 3380.500 3603.295 3381.470 3603.325 ;
        RECT 3380.670 3603.125 3381.470 3603.295 ;
        RECT 3380.500 3602.995 3381.470 3603.125 ;
        RECT 3382.070 3603.295 3383.390 3603.325 ;
        RECT 3382.070 3603.125 3383.220 3603.295 ;
        RECT 3383.390 3603.125 3384.190 3603.285 ;
        RECT 3382.070 3603.115 3384.190 3603.125 ;
        RECT 3382.070 3602.995 3383.390 3603.115 ;
        RECT 3380.500 3602.835 3380.670 3602.995 ;
        RECT 3383.220 3602.835 3383.390 3602.995 ;
        RECT 3384.410 3602.945 3384.580 3603.455 ;
        RECT 3377.780 3602.435 3377.950 3602.520 ;
        RECT 3380.500 3602.435 3380.670 3602.665 ;
        RECT 3383.220 3602.435 3383.390 3602.665 ;
        RECT 3383.560 3602.615 3384.580 3602.945 ;
      LAYER li1 ;
        RECT 3384.750 3602.660 3384.950 3603.760 ;
      LAYER li1 ;
        RECT 3385.120 3603.705 3385.290 3603.940 ;
        RECT 3385.460 3604.045 3385.940 3604.205 ;
        RECT 3385.460 3603.875 3386.110 3604.045 ;
        RECT 3385.940 3603.755 3386.110 3603.875 ;
        RECT 3385.120 3603.535 3385.765 3603.705 ;
        RECT 3385.120 3602.865 3385.290 3603.535 ;
        RECT 3385.940 3603.365 3386.110 3603.585 ;
        RECT 3385.460 3603.295 3386.110 3603.365 ;
        RECT 3385.460 3603.125 3385.940 3603.295 ;
        RECT 3385.460 3603.035 3386.110 3603.125 ;
        RECT 3385.120 3602.695 3385.770 3602.865 ;
        RECT 3385.940 3602.835 3386.110 3603.035 ;
        RECT 3385.940 3602.435 3386.110 3602.665 ;
        RECT 3377.780 3602.375 3379.115 3602.435 ;
        RECT 3377.950 3602.205 3379.115 3602.375 ;
        RECT 3377.780 3602.145 3379.115 3602.205 ;
        RECT 3379.775 3602.375 3381.395 3602.435 ;
        RECT 3379.775 3602.205 3380.500 3602.375 ;
        RECT 3380.670 3602.205 3381.395 3602.375 ;
        RECT 3379.775 3602.145 3381.395 3602.205 ;
        RECT 3382.055 3602.375 3384.555 3602.435 ;
        RECT 3382.055 3602.205 3383.220 3602.375 ;
        RECT 3383.390 3602.205 3384.555 3602.375 ;
        RECT 3382.055 3602.145 3384.555 3602.205 ;
        RECT 3385.215 3602.375 3386.110 3602.435 ;
        RECT 3385.215 3602.205 3385.940 3602.375 ;
        RECT 3385.215 3602.145 3386.110 3602.205 ;
        RECT 3377.780 3602.060 3377.950 3602.145 ;
        RECT 3380.500 3602.060 3380.670 3602.145 ;
        RECT 3383.220 3602.060 3383.390 3602.145 ;
        RECT 3385.940 3602.060 3386.110 3602.145 ;
        RECT 201.885 3050.885 202.055 3050.970 ;
        RECT 204.605 3050.885 204.775 3050.970 ;
        RECT 207.325 3050.885 207.495 3050.970 ;
        RECT 210.045 3050.885 210.215 3050.970 ;
        RECT 201.885 3050.825 202.780 3050.885 ;
        RECT 202.055 3050.655 202.780 3050.825 ;
        RECT 201.885 3050.595 202.780 3050.655 ;
        RECT 203.440 3050.825 205.940 3050.885 ;
        RECT 203.440 3050.655 204.605 3050.825 ;
        RECT 204.775 3050.655 205.940 3050.825 ;
        RECT 203.440 3050.595 205.940 3050.655 ;
        RECT 201.885 3050.365 202.055 3050.595 ;
        RECT 204.605 3050.365 204.775 3050.595 ;
        RECT 201.885 3050.035 202.055 3050.195 ;
        RECT 204.605 3050.035 204.775 3050.195 ;
        RECT 204.945 3050.085 205.965 3050.415 ;
        RECT 201.885 3049.905 202.855 3050.035 ;
        RECT 202.055 3049.735 202.855 3049.905 ;
        RECT 201.885 3049.705 202.855 3049.735 ;
        RECT 203.455 3049.915 204.775 3050.035 ;
        RECT 203.455 3049.905 205.575 3049.915 ;
        RECT 203.455 3049.735 204.605 3049.905 ;
        RECT 204.775 3049.745 205.575 3049.905 ;
        RECT 203.455 3049.705 204.775 3049.735 ;
        RECT 201.885 3049.445 202.055 3049.705 ;
      LAYER li1 ;
        RECT 202.225 3049.365 204.435 3049.535 ;
      LAYER li1 ;
        RECT 204.605 3049.445 204.775 3049.705 ;
        RECT 205.795 3049.575 205.965 3050.085 ;
      LAYER li1 ;
        RECT 202.705 3049.280 203.585 3049.365 ;
      LAYER li1 ;
        RECT 201.885 3049.195 202.055 3049.275 ;
        RECT 201.885 3048.985 202.535 3049.195 ;
        RECT 202.055 3048.865 202.535 3048.985 ;
        RECT 201.885 3048.525 202.055 3048.815 ;
      LAYER li1 ;
        RECT 202.705 3048.695 202.875 3049.280 ;
        RECT 202.225 3048.525 202.875 3048.695 ;
      LAYER li1 ;
        RECT 201.885 3048.065 202.535 3048.355 ;
        RECT 202.055 3048.025 202.535 3048.065 ;
        RECT 201.885 3047.605 202.055 3047.895 ;
      LAYER li1 ;
        RECT 202.705 3047.855 202.875 3048.525 ;
        RECT 202.225 3047.685 202.875 3047.855 ;
      LAYER li1 ;
        RECT 202.055 3047.435 202.535 3047.515 ;
        RECT 201.885 3047.185 202.535 3047.435 ;
        RECT 201.885 3047.145 202.055 3047.185 ;
      LAYER li1 ;
        RECT 202.705 3047.015 202.875 3047.685 ;
      LAYER li1 ;
        RECT 201.885 3046.685 202.055 3046.975 ;
      LAYER li1 ;
        RECT 202.225 3046.845 202.875 3047.015 ;
      LAYER li1 ;
        RECT 202.055 3046.515 202.535 3046.675 ;
        RECT 203.045 3046.585 203.215 3049.035 ;
      LAYER li1 ;
        RECT 203.415 3048.695 203.585 3049.280 ;
      LAYER li1 ;
        RECT 204.605 3049.195 204.775 3049.275 ;
        RECT 204.945 3049.245 205.965 3049.575 ;
      LAYER li1 ;
        RECT 206.135 3049.270 206.335 3050.860 ;
      LAYER li1 ;
        RECT 206.600 3050.825 208.220 3050.885 ;
        RECT 206.600 3050.655 207.325 3050.825 ;
        RECT 207.495 3050.655 208.220 3050.825 ;
        RECT 206.600 3050.595 208.220 3050.655 ;
        RECT 208.880 3050.825 210.215 3050.885 ;
        RECT 208.880 3050.655 210.045 3050.825 ;
        RECT 208.880 3050.595 210.215 3050.655 ;
        RECT 207.325 3050.365 207.495 3050.595 ;
        RECT 210.045 3050.510 210.215 3050.595 ;
        RECT 206.505 3050.165 207.155 3050.335 ;
        RECT 206.505 3049.495 206.675 3050.165 ;
        RECT 207.325 3049.995 207.495 3050.195 ;
        RECT 206.845 3049.905 207.495 3049.995 ;
        RECT 206.845 3049.735 207.325 3049.905 ;
        RECT 206.845 3049.665 207.495 3049.735 ;
        RECT 206.505 3049.325 207.150 3049.495 ;
        RECT 207.325 3049.445 207.495 3049.665 ;
        RECT 203.805 3049.075 204.775 3049.195 ;
        RECT 205.795 3049.090 205.965 3049.245 ;
        RECT 206.505 3049.090 206.675 3049.325 ;
        RECT 207.325 3049.155 207.495 3049.275 ;
        RECT 203.805 3048.985 205.575 3049.075 ;
        RECT 203.805 3048.865 204.605 3048.985 ;
        RECT 204.775 3048.905 205.575 3048.985 ;
        RECT 205.795 3048.915 206.675 3049.090 ;
        RECT 206.845 3048.985 207.495 3049.155 ;
      LAYER li1 ;
        RECT 203.415 3048.525 204.435 3048.695 ;
      LAYER li1 ;
        RECT 204.605 3048.525 204.775 3048.815 ;
      LAYER li1 ;
        RECT 203.415 3047.855 203.585 3048.525 ;
        RECT 204.945 3048.485 205.965 3048.655 ;
      LAYER li1 ;
        RECT 203.805 3048.315 204.775 3048.355 ;
        RECT 203.805 3048.065 205.575 3048.315 ;
        RECT 203.805 3048.025 204.605 3048.065 ;
        RECT 204.775 3047.985 205.575 3048.065 ;
      LAYER li1 ;
        RECT 203.415 3047.685 204.435 3047.855 ;
        RECT 203.415 3047.015 203.585 3047.685 ;
      LAYER li1 ;
        RECT 204.605 3047.605 204.775 3047.895 ;
      LAYER li1 ;
        RECT 205.795 3047.815 205.965 3048.485 ;
        RECT 204.945 3047.645 205.965 3047.815 ;
      LAYER li1 ;
        RECT 203.805 3047.435 204.605 3047.515 ;
        RECT 204.775 3047.435 205.575 3047.475 ;
        RECT 203.805 3047.185 205.575 3047.435 ;
        RECT 204.605 3047.145 205.575 3047.185 ;
      LAYER li1 ;
        RECT 203.415 3046.845 204.435 3047.015 ;
        RECT 205.795 3046.975 205.965 3047.645 ;
      LAYER li1 ;
        RECT 204.605 3046.685 204.775 3046.975 ;
      LAYER li1 ;
        RECT 204.945 3046.805 205.965 3046.975 ;
      LAYER li1 ;
        RECT 201.885 3046.345 202.535 3046.515 ;
        RECT 202.705 3046.410 203.585 3046.585 ;
        RECT 203.805 3046.515 204.605 3046.595 ;
        RECT 204.775 3046.515 205.575 3046.635 ;
        RECT 203.805 3046.425 205.575 3046.515 ;
        RECT 201.885 3046.225 202.055 3046.345 ;
        RECT 202.705 3046.175 202.875 3046.410 ;
        RECT 203.415 3046.255 203.585 3046.410 ;
        RECT 204.605 3046.305 205.575 3046.425 ;
        RECT 201.885 3045.835 202.055 3046.055 ;
        RECT 202.230 3046.005 202.875 3046.175 ;
        RECT 201.885 3045.765 202.535 3045.835 ;
        RECT 202.055 3045.595 202.535 3045.765 ;
        RECT 201.885 3045.505 202.535 3045.595 ;
        RECT 201.885 3045.305 202.055 3045.505 ;
        RECT 202.705 3045.335 202.875 3046.005 ;
        RECT 202.225 3045.165 202.875 3045.335 ;
        RECT 201.885 3044.905 202.055 3045.135 ;
      LAYER li1 ;
        RECT 203.045 3045.130 203.245 3046.230 ;
      LAYER li1 ;
        RECT 203.415 3045.925 204.435 3046.255 ;
        RECT 204.605 3046.225 204.775 3046.305 ;
      LAYER li1 ;
        RECT 205.795 3046.220 205.965 3046.805 ;
      LAYER li1 ;
        RECT 206.165 3046.465 206.335 3048.915 ;
        RECT 206.845 3048.825 207.325 3048.985 ;
      LAYER li1 ;
        RECT 207.495 3048.840 208.040 3050.425 ;
        RECT 206.505 3048.485 207.155 3048.655 ;
      LAYER li1 ;
        RECT 207.325 3048.525 207.495 3048.815 ;
      LAYER li1 ;
        RECT 207.495 3048.500 208.870 3048.840 ;
        RECT 206.505 3047.815 206.675 3048.485 ;
      LAYER li1 ;
        RECT 207.325 3048.315 207.495 3048.355 ;
        RECT 206.845 3048.065 207.495 3048.315 ;
        RECT 206.845 3047.985 207.325 3048.065 ;
      LAYER li1 ;
        RECT 206.505 3047.645 207.155 3047.815 ;
        RECT 206.505 3046.975 206.675 3047.645 ;
      LAYER li1 ;
        RECT 207.325 3047.605 207.495 3047.895 ;
        RECT 206.845 3047.435 207.325 3047.475 ;
        RECT 206.845 3047.145 207.495 3047.435 ;
      LAYER li1 ;
        RECT 206.505 3046.805 207.155 3046.975 ;
        RECT 206.505 3046.220 206.675 3046.805 ;
      LAYER li1 ;
        RECT 207.325 3046.685 207.495 3046.975 ;
        RECT 206.845 3046.515 207.325 3046.635 ;
        RECT 206.845 3046.305 207.495 3046.515 ;
        RECT 207.325 3046.225 207.495 3046.305 ;
      LAYER li1 ;
        RECT 205.795 3046.135 206.675 3046.220 ;
      LAYER li1 ;
        RECT 203.415 3045.415 203.585 3045.925 ;
        RECT 204.605 3045.795 204.775 3046.055 ;
      LAYER li1 ;
        RECT 204.945 3045.965 207.155 3046.135 ;
      LAYER li1 ;
        RECT 207.325 3045.795 207.495 3046.055 ;
        RECT 204.605 3045.765 205.925 3045.795 ;
        RECT 203.805 3045.595 204.605 3045.755 ;
        RECT 204.775 3045.595 205.925 3045.765 ;
        RECT 203.805 3045.585 205.925 3045.595 ;
        RECT 204.605 3045.465 205.925 3045.585 ;
        RECT 206.525 3045.765 207.495 3045.795 ;
        RECT 206.525 3045.595 207.325 3045.765 ;
        RECT 206.525 3045.465 207.495 3045.595 ;
        RECT 203.415 3045.085 204.435 3045.415 ;
        RECT 204.605 3045.305 204.775 3045.465 ;
        RECT 207.325 3045.305 207.495 3045.465 ;
        RECT 204.605 3044.905 204.775 3045.135 ;
        RECT 207.325 3044.905 207.495 3045.135 ;
      LAYER li1 ;
        RECT 207.495 3045.080 208.040 3048.500 ;
      LAYER li1 ;
        RECT 210.045 3044.905 210.215 3044.990 ;
        RECT 201.885 3044.845 202.780 3044.905 ;
        RECT 202.055 3044.675 202.780 3044.845 ;
        RECT 201.885 3044.615 202.780 3044.675 ;
        RECT 203.440 3044.845 205.940 3044.905 ;
        RECT 203.440 3044.675 204.605 3044.845 ;
        RECT 204.775 3044.675 205.940 3044.845 ;
        RECT 203.440 3044.615 205.940 3044.675 ;
        RECT 201.885 3044.385 202.055 3044.615 ;
        RECT 204.605 3044.385 204.775 3044.615 ;
        RECT 201.885 3044.055 202.055 3044.215 ;
        RECT 204.605 3044.055 204.775 3044.215 ;
        RECT 204.945 3044.105 205.965 3044.435 ;
        RECT 201.885 3043.925 202.855 3044.055 ;
        RECT 202.055 3043.755 202.855 3043.925 ;
        RECT 201.885 3043.725 202.855 3043.755 ;
        RECT 203.455 3043.935 204.775 3044.055 ;
        RECT 203.455 3043.925 205.575 3043.935 ;
        RECT 203.455 3043.755 204.605 3043.925 ;
        RECT 204.775 3043.765 205.575 3043.925 ;
        RECT 203.455 3043.725 204.775 3043.755 ;
        RECT 201.885 3043.465 202.055 3043.725 ;
      LAYER li1 ;
        RECT 202.225 3043.385 204.435 3043.555 ;
      LAYER li1 ;
        RECT 204.605 3043.465 204.775 3043.725 ;
        RECT 205.795 3043.595 205.965 3044.105 ;
      LAYER li1 ;
        RECT 202.705 3043.300 203.585 3043.385 ;
      LAYER li1 ;
        RECT 201.885 3043.215 202.055 3043.295 ;
        RECT 201.885 3043.005 202.535 3043.215 ;
        RECT 202.055 3042.885 202.535 3043.005 ;
        RECT 201.885 3042.545 202.055 3042.835 ;
      LAYER li1 ;
        RECT 202.705 3042.715 202.875 3043.300 ;
        RECT 202.225 3042.545 202.875 3042.715 ;
      LAYER li1 ;
        RECT 201.885 3042.085 202.535 3042.375 ;
        RECT 202.055 3042.045 202.535 3042.085 ;
        RECT 201.885 3041.625 202.055 3041.915 ;
      LAYER li1 ;
        RECT 202.705 3041.875 202.875 3042.545 ;
        RECT 202.225 3041.705 202.875 3041.875 ;
      LAYER li1 ;
        RECT 202.055 3041.455 202.535 3041.535 ;
        RECT 201.885 3041.205 202.535 3041.455 ;
        RECT 201.885 3041.165 202.055 3041.205 ;
      LAYER li1 ;
        RECT 202.705 3041.035 202.875 3041.705 ;
      LAYER li1 ;
        RECT 201.885 3040.705 202.055 3040.995 ;
      LAYER li1 ;
        RECT 202.225 3040.865 202.875 3041.035 ;
      LAYER li1 ;
        RECT 202.055 3040.535 202.535 3040.695 ;
        RECT 203.045 3040.605 203.215 3043.055 ;
      LAYER li1 ;
        RECT 203.415 3042.715 203.585 3043.300 ;
      LAYER li1 ;
        RECT 204.605 3043.215 204.775 3043.295 ;
        RECT 204.945 3043.265 205.965 3043.595 ;
      LAYER li1 ;
        RECT 206.135 3043.290 206.335 3044.880 ;
      LAYER li1 ;
        RECT 206.600 3044.845 208.220 3044.905 ;
        RECT 206.600 3044.675 207.325 3044.845 ;
        RECT 207.495 3044.675 208.220 3044.845 ;
        RECT 206.600 3044.615 208.220 3044.675 ;
        RECT 208.880 3044.845 210.215 3044.905 ;
        RECT 208.880 3044.675 210.045 3044.845 ;
        RECT 208.880 3044.615 210.215 3044.675 ;
        RECT 207.325 3044.385 207.495 3044.615 ;
        RECT 210.045 3044.530 210.215 3044.615 ;
        RECT 206.505 3044.185 207.155 3044.355 ;
        RECT 206.505 3043.515 206.675 3044.185 ;
        RECT 207.325 3044.015 207.495 3044.215 ;
        RECT 206.845 3043.925 207.495 3044.015 ;
        RECT 206.845 3043.755 207.325 3043.925 ;
        RECT 206.845 3043.685 207.495 3043.755 ;
        RECT 206.505 3043.345 207.150 3043.515 ;
        RECT 207.325 3043.465 207.495 3043.685 ;
        RECT 203.805 3043.095 204.775 3043.215 ;
        RECT 205.795 3043.110 205.965 3043.265 ;
        RECT 206.505 3043.110 206.675 3043.345 ;
        RECT 207.325 3043.175 207.495 3043.295 ;
        RECT 203.805 3043.005 205.575 3043.095 ;
        RECT 203.805 3042.885 204.605 3043.005 ;
        RECT 204.775 3042.925 205.575 3043.005 ;
        RECT 205.795 3042.935 206.675 3043.110 ;
        RECT 206.845 3043.005 207.495 3043.175 ;
      LAYER li1 ;
        RECT 203.415 3042.545 204.435 3042.715 ;
      LAYER li1 ;
        RECT 204.605 3042.545 204.775 3042.835 ;
      LAYER li1 ;
        RECT 203.415 3041.875 203.585 3042.545 ;
        RECT 204.945 3042.505 205.965 3042.675 ;
      LAYER li1 ;
        RECT 203.805 3042.335 204.775 3042.375 ;
        RECT 203.805 3042.085 205.575 3042.335 ;
        RECT 203.805 3042.045 204.605 3042.085 ;
        RECT 204.775 3042.005 205.575 3042.085 ;
      LAYER li1 ;
        RECT 203.415 3041.705 204.435 3041.875 ;
        RECT 203.415 3041.035 203.585 3041.705 ;
      LAYER li1 ;
        RECT 204.605 3041.625 204.775 3041.915 ;
      LAYER li1 ;
        RECT 205.795 3041.835 205.965 3042.505 ;
        RECT 204.945 3041.665 205.965 3041.835 ;
      LAYER li1 ;
        RECT 203.805 3041.455 204.605 3041.535 ;
        RECT 204.775 3041.455 205.575 3041.495 ;
        RECT 203.805 3041.205 205.575 3041.455 ;
        RECT 204.605 3041.165 205.575 3041.205 ;
      LAYER li1 ;
        RECT 203.415 3040.865 204.435 3041.035 ;
        RECT 205.795 3040.995 205.965 3041.665 ;
      LAYER li1 ;
        RECT 204.605 3040.705 204.775 3040.995 ;
      LAYER li1 ;
        RECT 204.945 3040.825 205.965 3040.995 ;
      LAYER li1 ;
        RECT 201.885 3040.365 202.535 3040.535 ;
        RECT 202.705 3040.430 203.585 3040.605 ;
        RECT 203.805 3040.535 204.605 3040.615 ;
        RECT 204.775 3040.535 205.575 3040.655 ;
        RECT 203.805 3040.445 205.575 3040.535 ;
        RECT 201.885 3040.245 202.055 3040.365 ;
        RECT 202.705 3040.195 202.875 3040.430 ;
        RECT 203.415 3040.275 203.585 3040.430 ;
        RECT 204.605 3040.325 205.575 3040.445 ;
        RECT 201.885 3039.855 202.055 3040.075 ;
        RECT 202.230 3040.025 202.875 3040.195 ;
        RECT 201.885 3039.785 202.535 3039.855 ;
        RECT 202.055 3039.615 202.535 3039.785 ;
        RECT 201.885 3039.525 202.535 3039.615 ;
        RECT 201.885 3039.325 202.055 3039.525 ;
        RECT 202.705 3039.355 202.875 3040.025 ;
        RECT 202.225 3039.185 202.875 3039.355 ;
        RECT 201.885 3038.925 202.055 3039.155 ;
      LAYER li1 ;
        RECT 203.045 3039.150 203.245 3040.250 ;
      LAYER li1 ;
        RECT 203.415 3039.945 204.435 3040.275 ;
        RECT 204.605 3040.245 204.775 3040.325 ;
      LAYER li1 ;
        RECT 205.795 3040.240 205.965 3040.825 ;
      LAYER li1 ;
        RECT 206.165 3040.485 206.335 3042.935 ;
        RECT 206.845 3042.845 207.325 3043.005 ;
      LAYER li1 ;
        RECT 207.495 3042.860 208.040 3044.445 ;
        RECT 206.505 3042.505 207.155 3042.675 ;
      LAYER li1 ;
        RECT 207.325 3042.545 207.495 3042.835 ;
      LAYER li1 ;
        RECT 207.495 3042.520 208.870 3042.860 ;
        RECT 206.505 3041.835 206.675 3042.505 ;
      LAYER li1 ;
        RECT 207.325 3042.335 207.495 3042.375 ;
        RECT 206.845 3042.085 207.495 3042.335 ;
        RECT 206.845 3042.005 207.325 3042.085 ;
      LAYER li1 ;
        RECT 206.505 3041.665 207.155 3041.835 ;
        RECT 206.505 3040.995 206.675 3041.665 ;
      LAYER li1 ;
        RECT 207.325 3041.625 207.495 3041.915 ;
        RECT 206.845 3041.455 207.325 3041.495 ;
        RECT 206.845 3041.165 207.495 3041.455 ;
      LAYER li1 ;
        RECT 206.505 3040.825 207.155 3040.995 ;
        RECT 206.505 3040.240 206.675 3040.825 ;
      LAYER li1 ;
        RECT 207.325 3040.705 207.495 3040.995 ;
        RECT 206.845 3040.535 207.325 3040.655 ;
        RECT 206.845 3040.325 207.495 3040.535 ;
        RECT 207.325 3040.245 207.495 3040.325 ;
      LAYER li1 ;
        RECT 205.795 3040.155 206.675 3040.240 ;
      LAYER li1 ;
        RECT 203.415 3039.435 203.585 3039.945 ;
        RECT 204.605 3039.815 204.775 3040.075 ;
      LAYER li1 ;
        RECT 204.945 3039.985 207.155 3040.155 ;
      LAYER li1 ;
        RECT 207.325 3039.815 207.495 3040.075 ;
        RECT 204.605 3039.785 205.925 3039.815 ;
        RECT 203.805 3039.615 204.605 3039.775 ;
        RECT 204.775 3039.615 205.925 3039.785 ;
        RECT 203.805 3039.605 205.925 3039.615 ;
        RECT 204.605 3039.485 205.925 3039.605 ;
        RECT 206.525 3039.785 207.495 3039.815 ;
        RECT 206.525 3039.615 207.325 3039.785 ;
        RECT 206.525 3039.485 207.495 3039.615 ;
        RECT 203.415 3039.105 204.435 3039.435 ;
        RECT 204.605 3039.325 204.775 3039.485 ;
        RECT 207.325 3039.325 207.495 3039.485 ;
        RECT 204.605 3038.925 204.775 3039.155 ;
        RECT 207.325 3038.925 207.495 3039.155 ;
      LAYER li1 ;
        RECT 207.495 3039.100 208.040 3042.520 ;
      LAYER li1 ;
        RECT 210.045 3038.925 210.215 3039.010 ;
        RECT 201.885 3038.865 202.780 3038.925 ;
        RECT 202.055 3038.695 202.780 3038.865 ;
        RECT 201.885 3038.635 202.780 3038.695 ;
        RECT 203.440 3038.865 205.940 3038.925 ;
        RECT 203.440 3038.695 204.605 3038.865 ;
        RECT 204.775 3038.695 205.940 3038.865 ;
        RECT 203.440 3038.635 205.940 3038.695 ;
        RECT 201.885 3038.405 202.055 3038.635 ;
        RECT 204.605 3038.405 204.775 3038.635 ;
        RECT 201.885 3038.075 202.055 3038.235 ;
        RECT 204.605 3038.075 204.775 3038.235 ;
        RECT 204.945 3038.125 205.965 3038.455 ;
        RECT 201.885 3037.945 202.855 3038.075 ;
        RECT 202.055 3037.775 202.855 3037.945 ;
        RECT 201.885 3037.745 202.855 3037.775 ;
        RECT 203.455 3037.955 204.775 3038.075 ;
        RECT 203.455 3037.945 205.575 3037.955 ;
        RECT 203.455 3037.775 204.605 3037.945 ;
        RECT 204.775 3037.785 205.575 3037.945 ;
        RECT 203.455 3037.745 204.775 3037.775 ;
        RECT 201.885 3037.485 202.055 3037.745 ;
      LAYER li1 ;
        RECT 202.225 3037.405 204.435 3037.575 ;
      LAYER li1 ;
        RECT 204.605 3037.485 204.775 3037.745 ;
        RECT 205.795 3037.615 205.965 3038.125 ;
      LAYER li1 ;
        RECT 202.705 3037.320 203.585 3037.405 ;
      LAYER li1 ;
        RECT 201.885 3037.235 202.055 3037.315 ;
        RECT 201.885 3037.025 202.535 3037.235 ;
        RECT 202.055 3036.905 202.535 3037.025 ;
        RECT 201.885 3036.565 202.055 3036.855 ;
      LAYER li1 ;
        RECT 202.705 3036.735 202.875 3037.320 ;
        RECT 202.225 3036.565 202.875 3036.735 ;
      LAYER li1 ;
        RECT 201.885 3036.105 202.535 3036.395 ;
        RECT 202.055 3036.065 202.535 3036.105 ;
        RECT 201.885 3035.645 202.055 3035.935 ;
      LAYER li1 ;
        RECT 202.705 3035.895 202.875 3036.565 ;
        RECT 202.225 3035.725 202.875 3035.895 ;
      LAYER li1 ;
        RECT 202.055 3035.475 202.535 3035.555 ;
        RECT 201.885 3035.225 202.535 3035.475 ;
        RECT 201.885 3035.185 202.055 3035.225 ;
      LAYER li1 ;
        RECT 202.705 3035.055 202.875 3035.725 ;
      LAYER li1 ;
        RECT 201.885 3034.725 202.055 3035.015 ;
      LAYER li1 ;
        RECT 202.225 3034.885 202.875 3035.055 ;
      LAYER li1 ;
        RECT 202.055 3034.555 202.535 3034.715 ;
        RECT 203.045 3034.625 203.215 3037.075 ;
      LAYER li1 ;
        RECT 203.415 3036.735 203.585 3037.320 ;
      LAYER li1 ;
        RECT 204.605 3037.235 204.775 3037.315 ;
        RECT 204.945 3037.285 205.965 3037.615 ;
      LAYER li1 ;
        RECT 206.135 3037.310 206.335 3038.900 ;
      LAYER li1 ;
        RECT 206.600 3038.865 208.220 3038.925 ;
        RECT 206.600 3038.695 207.325 3038.865 ;
        RECT 207.495 3038.695 208.220 3038.865 ;
        RECT 206.600 3038.635 208.220 3038.695 ;
        RECT 208.880 3038.865 210.215 3038.925 ;
        RECT 208.880 3038.695 210.045 3038.865 ;
        RECT 208.880 3038.635 210.215 3038.695 ;
        RECT 207.325 3038.405 207.495 3038.635 ;
        RECT 210.045 3038.550 210.215 3038.635 ;
        RECT 206.505 3038.205 207.155 3038.375 ;
        RECT 206.505 3037.535 206.675 3038.205 ;
        RECT 207.325 3038.035 207.495 3038.235 ;
        RECT 206.845 3037.945 207.495 3038.035 ;
        RECT 206.845 3037.775 207.325 3037.945 ;
        RECT 206.845 3037.705 207.495 3037.775 ;
        RECT 206.505 3037.365 207.150 3037.535 ;
        RECT 207.325 3037.485 207.495 3037.705 ;
        RECT 203.805 3037.115 204.775 3037.235 ;
        RECT 205.795 3037.130 205.965 3037.285 ;
        RECT 206.505 3037.130 206.675 3037.365 ;
        RECT 207.325 3037.195 207.495 3037.315 ;
        RECT 203.805 3037.025 205.575 3037.115 ;
        RECT 203.805 3036.905 204.605 3037.025 ;
        RECT 204.775 3036.945 205.575 3037.025 ;
        RECT 205.795 3036.955 206.675 3037.130 ;
        RECT 206.845 3037.025 207.495 3037.195 ;
      LAYER li1 ;
        RECT 203.415 3036.565 204.435 3036.735 ;
      LAYER li1 ;
        RECT 204.605 3036.565 204.775 3036.855 ;
      LAYER li1 ;
        RECT 203.415 3035.895 203.585 3036.565 ;
        RECT 204.945 3036.525 205.965 3036.695 ;
      LAYER li1 ;
        RECT 203.805 3036.355 204.775 3036.395 ;
        RECT 203.805 3036.105 205.575 3036.355 ;
        RECT 203.805 3036.065 204.605 3036.105 ;
        RECT 204.775 3036.025 205.575 3036.105 ;
      LAYER li1 ;
        RECT 203.415 3035.725 204.435 3035.895 ;
        RECT 203.415 3035.055 203.585 3035.725 ;
      LAYER li1 ;
        RECT 204.605 3035.645 204.775 3035.935 ;
      LAYER li1 ;
        RECT 205.795 3035.855 205.965 3036.525 ;
        RECT 204.945 3035.685 205.965 3035.855 ;
      LAYER li1 ;
        RECT 203.805 3035.475 204.605 3035.555 ;
        RECT 204.775 3035.475 205.575 3035.515 ;
        RECT 203.805 3035.225 205.575 3035.475 ;
        RECT 204.605 3035.185 205.575 3035.225 ;
      LAYER li1 ;
        RECT 203.415 3034.885 204.435 3035.055 ;
        RECT 205.795 3035.015 205.965 3035.685 ;
      LAYER li1 ;
        RECT 204.605 3034.725 204.775 3035.015 ;
      LAYER li1 ;
        RECT 204.945 3034.845 205.965 3035.015 ;
      LAYER li1 ;
        RECT 201.885 3034.385 202.535 3034.555 ;
        RECT 202.705 3034.450 203.585 3034.625 ;
        RECT 203.805 3034.555 204.605 3034.635 ;
        RECT 204.775 3034.555 205.575 3034.675 ;
        RECT 203.805 3034.465 205.575 3034.555 ;
        RECT 201.885 3034.265 202.055 3034.385 ;
        RECT 202.705 3034.215 202.875 3034.450 ;
        RECT 203.415 3034.295 203.585 3034.450 ;
        RECT 204.605 3034.345 205.575 3034.465 ;
        RECT 201.885 3033.875 202.055 3034.095 ;
        RECT 202.230 3034.045 202.875 3034.215 ;
        RECT 201.885 3033.805 202.535 3033.875 ;
        RECT 202.055 3033.635 202.535 3033.805 ;
        RECT 201.885 3033.545 202.535 3033.635 ;
        RECT 201.885 3033.345 202.055 3033.545 ;
        RECT 202.705 3033.375 202.875 3034.045 ;
        RECT 202.225 3033.205 202.875 3033.375 ;
        RECT 201.885 3032.945 202.055 3033.175 ;
      LAYER li1 ;
        RECT 203.045 3033.170 203.245 3034.270 ;
      LAYER li1 ;
        RECT 203.415 3033.965 204.435 3034.295 ;
        RECT 204.605 3034.265 204.775 3034.345 ;
      LAYER li1 ;
        RECT 205.795 3034.260 205.965 3034.845 ;
      LAYER li1 ;
        RECT 206.165 3034.505 206.335 3036.955 ;
        RECT 206.845 3036.865 207.325 3037.025 ;
      LAYER li1 ;
        RECT 207.495 3036.880 208.040 3038.465 ;
        RECT 206.505 3036.525 207.155 3036.695 ;
      LAYER li1 ;
        RECT 207.325 3036.565 207.495 3036.855 ;
      LAYER li1 ;
        RECT 207.495 3036.540 208.870 3036.880 ;
        RECT 206.505 3035.855 206.675 3036.525 ;
      LAYER li1 ;
        RECT 207.325 3036.355 207.495 3036.395 ;
        RECT 206.845 3036.105 207.495 3036.355 ;
        RECT 206.845 3036.025 207.325 3036.105 ;
      LAYER li1 ;
        RECT 206.505 3035.685 207.155 3035.855 ;
        RECT 206.505 3035.015 206.675 3035.685 ;
      LAYER li1 ;
        RECT 207.325 3035.645 207.495 3035.935 ;
        RECT 206.845 3035.475 207.325 3035.515 ;
        RECT 206.845 3035.185 207.495 3035.475 ;
      LAYER li1 ;
        RECT 206.505 3034.845 207.155 3035.015 ;
        RECT 206.505 3034.260 206.675 3034.845 ;
      LAYER li1 ;
        RECT 207.325 3034.725 207.495 3035.015 ;
        RECT 206.845 3034.555 207.325 3034.675 ;
        RECT 206.845 3034.345 207.495 3034.555 ;
        RECT 207.325 3034.265 207.495 3034.345 ;
      LAYER li1 ;
        RECT 205.795 3034.175 206.675 3034.260 ;
      LAYER li1 ;
        RECT 203.415 3033.455 203.585 3033.965 ;
        RECT 204.605 3033.835 204.775 3034.095 ;
      LAYER li1 ;
        RECT 204.945 3034.005 207.155 3034.175 ;
      LAYER li1 ;
        RECT 207.325 3033.835 207.495 3034.095 ;
        RECT 204.605 3033.805 205.925 3033.835 ;
        RECT 203.805 3033.635 204.605 3033.795 ;
        RECT 204.775 3033.635 205.925 3033.805 ;
        RECT 203.805 3033.625 205.925 3033.635 ;
        RECT 204.605 3033.505 205.925 3033.625 ;
        RECT 206.525 3033.805 207.495 3033.835 ;
        RECT 206.525 3033.635 207.325 3033.805 ;
        RECT 206.525 3033.505 207.495 3033.635 ;
        RECT 203.415 3033.125 204.435 3033.455 ;
        RECT 204.605 3033.345 204.775 3033.505 ;
        RECT 207.325 3033.345 207.495 3033.505 ;
        RECT 204.605 3032.945 204.775 3033.175 ;
        RECT 207.325 3032.945 207.495 3033.175 ;
      LAYER li1 ;
        RECT 207.495 3033.120 208.040 3036.540 ;
      LAYER li1 ;
        RECT 210.045 3032.945 210.215 3033.030 ;
        RECT 201.885 3032.885 202.780 3032.945 ;
        RECT 202.055 3032.715 202.780 3032.885 ;
        RECT 201.885 3032.655 202.780 3032.715 ;
        RECT 203.440 3032.885 205.940 3032.945 ;
        RECT 203.440 3032.715 204.605 3032.885 ;
        RECT 204.775 3032.715 205.940 3032.885 ;
        RECT 203.440 3032.655 205.940 3032.715 ;
        RECT 201.885 3032.425 202.055 3032.655 ;
        RECT 204.605 3032.425 204.775 3032.655 ;
        RECT 201.885 3032.095 202.055 3032.255 ;
        RECT 204.605 3032.095 204.775 3032.255 ;
        RECT 204.945 3032.145 205.965 3032.475 ;
        RECT 201.885 3031.965 202.855 3032.095 ;
        RECT 202.055 3031.795 202.855 3031.965 ;
        RECT 201.885 3031.765 202.855 3031.795 ;
        RECT 203.455 3031.975 204.775 3032.095 ;
        RECT 203.455 3031.965 205.575 3031.975 ;
        RECT 203.455 3031.795 204.605 3031.965 ;
        RECT 204.775 3031.805 205.575 3031.965 ;
        RECT 203.455 3031.765 204.775 3031.795 ;
        RECT 201.885 3031.505 202.055 3031.765 ;
      LAYER li1 ;
        RECT 202.225 3031.425 204.435 3031.595 ;
      LAYER li1 ;
        RECT 204.605 3031.505 204.775 3031.765 ;
        RECT 205.795 3031.635 205.965 3032.145 ;
      LAYER li1 ;
        RECT 202.705 3031.340 203.585 3031.425 ;
      LAYER li1 ;
        RECT 201.885 3031.255 202.055 3031.335 ;
        RECT 201.885 3031.045 202.535 3031.255 ;
        RECT 202.055 3030.925 202.535 3031.045 ;
        RECT 201.885 3030.585 202.055 3030.875 ;
      LAYER li1 ;
        RECT 202.705 3030.755 202.875 3031.340 ;
        RECT 202.225 3030.585 202.875 3030.755 ;
      LAYER li1 ;
        RECT 201.885 3030.125 202.535 3030.415 ;
        RECT 202.055 3030.085 202.535 3030.125 ;
        RECT 201.885 3029.665 202.055 3029.955 ;
      LAYER li1 ;
        RECT 202.705 3029.915 202.875 3030.585 ;
        RECT 202.225 3029.745 202.875 3029.915 ;
      LAYER li1 ;
        RECT 202.055 3029.495 202.535 3029.575 ;
        RECT 201.885 3029.245 202.535 3029.495 ;
        RECT 201.885 3029.205 202.055 3029.245 ;
      LAYER li1 ;
        RECT 202.705 3029.075 202.875 3029.745 ;
      LAYER li1 ;
        RECT 201.885 3028.745 202.055 3029.035 ;
      LAYER li1 ;
        RECT 202.225 3028.905 202.875 3029.075 ;
      LAYER li1 ;
        RECT 202.055 3028.575 202.535 3028.735 ;
        RECT 203.045 3028.645 203.215 3031.095 ;
      LAYER li1 ;
        RECT 203.415 3030.755 203.585 3031.340 ;
      LAYER li1 ;
        RECT 204.605 3031.255 204.775 3031.335 ;
        RECT 204.945 3031.305 205.965 3031.635 ;
      LAYER li1 ;
        RECT 206.135 3031.330 206.335 3032.920 ;
      LAYER li1 ;
        RECT 206.600 3032.885 208.220 3032.945 ;
        RECT 206.600 3032.715 207.325 3032.885 ;
        RECT 207.495 3032.715 208.220 3032.885 ;
        RECT 206.600 3032.655 208.220 3032.715 ;
        RECT 208.880 3032.885 210.215 3032.945 ;
        RECT 208.880 3032.715 210.045 3032.885 ;
        RECT 208.880 3032.655 210.215 3032.715 ;
        RECT 207.325 3032.425 207.495 3032.655 ;
        RECT 210.045 3032.570 210.215 3032.655 ;
        RECT 206.505 3032.225 207.155 3032.395 ;
        RECT 206.505 3031.555 206.675 3032.225 ;
        RECT 207.325 3032.055 207.495 3032.255 ;
        RECT 206.845 3031.965 207.495 3032.055 ;
        RECT 206.845 3031.795 207.325 3031.965 ;
        RECT 206.845 3031.725 207.495 3031.795 ;
        RECT 206.505 3031.385 207.150 3031.555 ;
        RECT 207.325 3031.505 207.495 3031.725 ;
        RECT 203.805 3031.135 204.775 3031.255 ;
        RECT 205.795 3031.150 205.965 3031.305 ;
        RECT 206.505 3031.150 206.675 3031.385 ;
        RECT 207.325 3031.215 207.495 3031.335 ;
        RECT 203.805 3031.045 205.575 3031.135 ;
        RECT 203.805 3030.925 204.605 3031.045 ;
        RECT 204.775 3030.965 205.575 3031.045 ;
        RECT 205.795 3030.975 206.675 3031.150 ;
        RECT 206.845 3031.045 207.495 3031.215 ;
      LAYER li1 ;
        RECT 203.415 3030.585 204.435 3030.755 ;
      LAYER li1 ;
        RECT 204.605 3030.585 204.775 3030.875 ;
      LAYER li1 ;
        RECT 203.415 3029.915 203.585 3030.585 ;
        RECT 204.945 3030.545 205.965 3030.715 ;
      LAYER li1 ;
        RECT 203.805 3030.375 204.775 3030.415 ;
        RECT 203.805 3030.125 205.575 3030.375 ;
        RECT 203.805 3030.085 204.605 3030.125 ;
        RECT 204.775 3030.045 205.575 3030.125 ;
      LAYER li1 ;
        RECT 203.415 3029.745 204.435 3029.915 ;
        RECT 203.415 3029.075 203.585 3029.745 ;
      LAYER li1 ;
        RECT 204.605 3029.665 204.775 3029.955 ;
      LAYER li1 ;
        RECT 205.795 3029.875 205.965 3030.545 ;
        RECT 204.945 3029.705 205.965 3029.875 ;
      LAYER li1 ;
        RECT 203.805 3029.495 204.605 3029.575 ;
        RECT 204.775 3029.495 205.575 3029.535 ;
        RECT 203.805 3029.245 205.575 3029.495 ;
        RECT 204.605 3029.205 205.575 3029.245 ;
      LAYER li1 ;
        RECT 203.415 3028.905 204.435 3029.075 ;
        RECT 205.795 3029.035 205.965 3029.705 ;
      LAYER li1 ;
        RECT 204.605 3028.745 204.775 3029.035 ;
      LAYER li1 ;
        RECT 204.945 3028.865 205.965 3029.035 ;
      LAYER li1 ;
        RECT 201.885 3028.405 202.535 3028.575 ;
        RECT 202.705 3028.470 203.585 3028.645 ;
        RECT 203.805 3028.575 204.605 3028.655 ;
        RECT 204.775 3028.575 205.575 3028.695 ;
        RECT 203.805 3028.485 205.575 3028.575 ;
        RECT 201.885 3028.285 202.055 3028.405 ;
        RECT 202.705 3028.235 202.875 3028.470 ;
        RECT 203.415 3028.315 203.585 3028.470 ;
        RECT 204.605 3028.365 205.575 3028.485 ;
        RECT 201.885 3027.895 202.055 3028.115 ;
        RECT 202.230 3028.065 202.875 3028.235 ;
        RECT 201.885 3027.825 202.535 3027.895 ;
        RECT 202.055 3027.655 202.535 3027.825 ;
        RECT 201.885 3027.565 202.535 3027.655 ;
        RECT 201.885 3027.365 202.055 3027.565 ;
        RECT 202.705 3027.395 202.875 3028.065 ;
        RECT 202.225 3027.225 202.875 3027.395 ;
        RECT 201.885 3026.965 202.055 3027.195 ;
      LAYER li1 ;
        RECT 203.045 3027.190 203.245 3028.290 ;
      LAYER li1 ;
        RECT 203.415 3027.985 204.435 3028.315 ;
        RECT 204.605 3028.285 204.775 3028.365 ;
      LAYER li1 ;
        RECT 205.795 3028.280 205.965 3028.865 ;
      LAYER li1 ;
        RECT 206.165 3028.525 206.335 3030.975 ;
        RECT 206.845 3030.885 207.325 3031.045 ;
      LAYER li1 ;
        RECT 207.495 3030.900 208.040 3032.485 ;
        RECT 206.505 3030.545 207.155 3030.715 ;
      LAYER li1 ;
        RECT 207.325 3030.585 207.495 3030.875 ;
      LAYER li1 ;
        RECT 207.495 3030.560 208.870 3030.900 ;
        RECT 206.505 3029.875 206.675 3030.545 ;
      LAYER li1 ;
        RECT 207.325 3030.375 207.495 3030.415 ;
        RECT 206.845 3030.125 207.495 3030.375 ;
        RECT 206.845 3030.045 207.325 3030.125 ;
      LAYER li1 ;
        RECT 206.505 3029.705 207.155 3029.875 ;
        RECT 206.505 3029.035 206.675 3029.705 ;
      LAYER li1 ;
        RECT 207.325 3029.665 207.495 3029.955 ;
        RECT 206.845 3029.495 207.325 3029.535 ;
        RECT 206.845 3029.205 207.495 3029.495 ;
      LAYER li1 ;
        RECT 206.505 3028.865 207.155 3029.035 ;
        RECT 206.505 3028.280 206.675 3028.865 ;
      LAYER li1 ;
        RECT 207.325 3028.745 207.495 3029.035 ;
        RECT 206.845 3028.575 207.325 3028.695 ;
        RECT 206.845 3028.365 207.495 3028.575 ;
        RECT 207.325 3028.285 207.495 3028.365 ;
      LAYER li1 ;
        RECT 205.795 3028.195 206.675 3028.280 ;
      LAYER li1 ;
        RECT 203.415 3027.475 203.585 3027.985 ;
        RECT 204.605 3027.855 204.775 3028.115 ;
      LAYER li1 ;
        RECT 204.945 3028.025 207.155 3028.195 ;
      LAYER li1 ;
        RECT 207.325 3027.855 207.495 3028.115 ;
        RECT 204.605 3027.825 205.925 3027.855 ;
        RECT 203.805 3027.655 204.605 3027.815 ;
        RECT 204.775 3027.655 205.925 3027.825 ;
        RECT 203.805 3027.645 205.925 3027.655 ;
        RECT 204.605 3027.525 205.925 3027.645 ;
        RECT 206.525 3027.825 207.495 3027.855 ;
        RECT 206.525 3027.655 207.325 3027.825 ;
        RECT 206.525 3027.525 207.495 3027.655 ;
        RECT 203.415 3027.145 204.435 3027.475 ;
        RECT 204.605 3027.365 204.775 3027.525 ;
        RECT 207.325 3027.365 207.495 3027.525 ;
        RECT 204.605 3026.965 204.775 3027.195 ;
        RECT 207.325 3026.965 207.495 3027.195 ;
      LAYER li1 ;
        RECT 207.495 3027.140 208.040 3030.560 ;
      LAYER li1 ;
        RECT 210.045 3026.965 210.215 3027.050 ;
        RECT 201.885 3026.905 202.780 3026.965 ;
        RECT 202.055 3026.735 202.780 3026.905 ;
        RECT 201.885 3026.675 202.780 3026.735 ;
        RECT 203.440 3026.905 205.940 3026.965 ;
        RECT 203.440 3026.735 204.605 3026.905 ;
        RECT 204.775 3026.735 205.940 3026.905 ;
        RECT 203.440 3026.675 205.940 3026.735 ;
        RECT 201.885 3026.445 202.055 3026.675 ;
        RECT 204.605 3026.445 204.775 3026.675 ;
        RECT 201.885 3026.115 202.055 3026.275 ;
        RECT 204.605 3026.115 204.775 3026.275 ;
        RECT 204.945 3026.165 205.965 3026.495 ;
        RECT 201.885 3025.985 202.855 3026.115 ;
        RECT 202.055 3025.815 202.855 3025.985 ;
        RECT 201.885 3025.785 202.855 3025.815 ;
        RECT 203.455 3025.995 204.775 3026.115 ;
        RECT 203.455 3025.985 205.575 3025.995 ;
        RECT 203.455 3025.815 204.605 3025.985 ;
        RECT 204.775 3025.825 205.575 3025.985 ;
        RECT 203.455 3025.785 204.775 3025.815 ;
        RECT 201.885 3025.525 202.055 3025.785 ;
      LAYER li1 ;
        RECT 202.225 3025.445 204.435 3025.615 ;
      LAYER li1 ;
        RECT 204.605 3025.525 204.775 3025.785 ;
        RECT 205.795 3025.655 205.965 3026.165 ;
      LAYER li1 ;
        RECT 202.705 3025.360 203.585 3025.445 ;
      LAYER li1 ;
        RECT 201.885 3025.275 202.055 3025.355 ;
        RECT 201.885 3025.065 202.535 3025.275 ;
        RECT 202.055 3024.945 202.535 3025.065 ;
        RECT 201.885 3024.605 202.055 3024.895 ;
      LAYER li1 ;
        RECT 202.705 3024.775 202.875 3025.360 ;
        RECT 202.225 3024.605 202.875 3024.775 ;
      LAYER li1 ;
        RECT 201.885 3024.145 202.535 3024.435 ;
        RECT 202.055 3024.105 202.535 3024.145 ;
        RECT 201.885 3023.685 202.055 3023.975 ;
      LAYER li1 ;
        RECT 202.705 3023.935 202.875 3024.605 ;
        RECT 202.225 3023.765 202.875 3023.935 ;
      LAYER li1 ;
        RECT 202.055 3023.515 202.535 3023.595 ;
        RECT 201.885 3023.265 202.535 3023.515 ;
        RECT 201.885 3023.225 202.055 3023.265 ;
      LAYER li1 ;
        RECT 202.705 3023.095 202.875 3023.765 ;
      LAYER li1 ;
        RECT 201.885 3022.765 202.055 3023.055 ;
      LAYER li1 ;
        RECT 202.225 3022.925 202.875 3023.095 ;
      LAYER li1 ;
        RECT 202.055 3022.595 202.535 3022.755 ;
        RECT 203.045 3022.665 203.215 3025.115 ;
      LAYER li1 ;
        RECT 203.415 3024.775 203.585 3025.360 ;
      LAYER li1 ;
        RECT 204.605 3025.275 204.775 3025.355 ;
        RECT 204.945 3025.325 205.965 3025.655 ;
      LAYER li1 ;
        RECT 206.135 3025.350 206.335 3026.940 ;
      LAYER li1 ;
        RECT 206.600 3026.905 208.220 3026.965 ;
        RECT 206.600 3026.735 207.325 3026.905 ;
        RECT 207.495 3026.735 208.220 3026.905 ;
        RECT 206.600 3026.675 208.220 3026.735 ;
        RECT 208.880 3026.905 210.215 3026.965 ;
        RECT 208.880 3026.735 210.045 3026.905 ;
        RECT 208.880 3026.675 210.215 3026.735 ;
        RECT 207.325 3026.445 207.495 3026.675 ;
        RECT 210.045 3026.590 210.215 3026.675 ;
        RECT 206.505 3026.245 207.155 3026.415 ;
        RECT 206.505 3025.575 206.675 3026.245 ;
        RECT 207.325 3026.075 207.495 3026.275 ;
        RECT 206.845 3025.985 207.495 3026.075 ;
        RECT 206.845 3025.815 207.325 3025.985 ;
        RECT 206.845 3025.745 207.495 3025.815 ;
        RECT 206.505 3025.405 207.150 3025.575 ;
        RECT 207.325 3025.525 207.495 3025.745 ;
        RECT 203.805 3025.155 204.775 3025.275 ;
        RECT 205.795 3025.170 205.965 3025.325 ;
        RECT 206.505 3025.170 206.675 3025.405 ;
        RECT 207.325 3025.235 207.495 3025.355 ;
        RECT 203.805 3025.065 205.575 3025.155 ;
        RECT 203.805 3024.945 204.605 3025.065 ;
        RECT 204.775 3024.985 205.575 3025.065 ;
        RECT 205.795 3024.995 206.675 3025.170 ;
        RECT 206.845 3025.065 207.495 3025.235 ;
      LAYER li1 ;
        RECT 203.415 3024.605 204.435 3024.775 ;
      LAYER li1 ;
        RECT 204.605 3024.605 204.775 3024.895 ;
      LAYER li1 ;
        RECT 203.415 3023.935 203.585 3024.605 ;
        RECT 204.945 3024.565 205.965 3024.735 ;
      LAYER li1 ;
        RECT 203.805 3024.395 204.775 3024.435 ;
        RECT 203.805 3024.145 205.575 3024.395 ;
        RECT 203.805 3024.105 204.605 3024.145 ;
        RECT 204.775 3024.065 205.575 3024.145 ;
      LAYER li1 ;
        RECT 203.415 3023.765 204.435 3023.935 ;
        RECT 203.415 3023.095 203.585 3023.765 ;
      LAYER li1 ;
        RECT 204.605 3023.685 204.775 3023.975 ;
      LAYER li1 ;
        RECT 205.795 3023.895 205.965 3024.565 ;
        RECT 204.945 3023.725 205.965 3023.895 ;
      LAYER li1 ;
        RECT 203.805 3023.515 204.605 3023.595 ;
        RECT 204.775 3023.515 205.575 3023.555 ;
        RECT 203.805 3023.265 205.575 3023.515 ;
        RECT 204.605 3023.225 205.575 3023.265 ;
      LAYER li1 ;
        RECT 203.415 3022.925 204.435 3023.095 ;
        RECT 205.795 3023.055 205.965 3023.725 ;
      LAYER li1 ;
        RECT 204.605 3022.765 204.775 3023.055 ;
      LAYER li1 ;
        RECT 204.945 3022.885 205.965 3023.055 ;
      LAYER li1 ;
        RECT 201.885 3022.425 202.535 3022.595 ;
        RECT 202.705 3022.490 203.585 3022.665 ;
        RECT 203.805 3022.595 204.605 3022.675 ;
        RECT 204.775 3022.595 205.575 3022.715 ;
        RECT 203.805 3022.505 205.575 3022.595 ;
        RECT 201.885 3022.305 202.055 3022.425 ;
        RECT 202.705 3022.255 202.875 3022.490 ;
        RECT 203.415 3022.335 203.585 3022.490 ;
        RECT 204.605 3022.385 205.575 3022.505 ;
        RECT 201.885 3021.915 202.055 3022.135 ;
        RECT 202.230 3022.085 202.875 3022.255 ;
        RECT 201.885 3021.845 202.535 3021.915 ;
        RECT 202.055 3021.675 202.535 3021.845 ;
        RECT 201.885 3021.585 202.535 3021.675 ;
        RECT 201.885 3021.385 202.055 3021.585 ;
        RECT 202.705 3021.415 202.875 3022.085 ;
        RECT 202.225 3021.245 202.875 3021.415 ;
        RECT 201.885 3020.985 202.055 3021.215 ;
      LAYER li1 ;
        RECT 203.045 3021.210 203.245 3022.310 ;
      LAYER li1 ;
        RECT 203.415 3022.005 204.435 3022.335 ;
        RECT 204.605 3022.305 204.775 3022.385 ;
      LAYER li1 ;
        RECT 205.795 3022.300 205.965 3022.885 ;
      LAYER li1 ;
        RECT 206.165 3022.545 206.335 3024.995 ;
        RECT 206.845 3024.905 207.325 3025.065 ;
      LAYER li1 ;
        RECT 207.495 3024.920 208.040 3026.505 ;
        RECT 206.505 3024.565 207.155 3024.735 ;
      LAYER li1 ;
        RECT 207.325 3024.605 207.495 3024.895 ;
      LAYER li1 ;
        RECT 207.495 3024.580 208.870 3024.920 ;
        RECT 206.505 3023.895 206.675 3024.565 ;
      LAYER li1 ;
        RECT 207.325 3024.395 207.495 3024.435 ;
        RECT 206.845 3024.145 207.495 3024.395 ;
        RECT 206.845 3024.065 207.325 3024.145 ;
      LAYER li1 ;
        RECT 206.505 3023.725 207.155 3023.895 ;
        RECT 206.505 3023.055 206.675 3023.725 ;
      LAYER li1 ;
        RECT 207.325 3023.685 207.495 3023.975 ;
        RECT 206.845 3023.515 207.325 3023.555 ;
        RECT 206.845 3023.225 207.495 3023.515 ;
      LAYER li1 ;
        RECT 206.505 3022.885 207.155 3023.055 ;
        RECT 206.505 3022.300 206.675 3022.885 ;
      LAYER li1 ;
        RECT 207.325 3022.765 207.495 3023.055 ;
        RECT 206.845 3022.595 207.325 3022.715 ;
        RECT 206.845 3022.385 207.495 3022.595 ;
        RECT 207.325 3022.305 207.495 3022.385 ;
      LAYER li1 ;
        RECT 205.795 3022.215 206.675 3022.300 ;
      LAYER li1 ;
        RECT 203.415 3021.495 203.585 3022.005 ;
        RECT 204.605 3021.875 204.775 3022.135 ;
      LAYER li1 ;
        RECT 204.945 3022.045 207.155 3022.215 ;
      LAYER li1 ;
        RECT 207.325 3021.875 207.495 3022.135 ;
        RECT 204.605 3021.845 205.925 3021.875 ;
        RECT 203.805 3021.675 204.605 3021.835 ;
        RECT 204.775 3021.675 205.925 3021.845 ;
        RECT 203.805 3021.665 205.925 3021.675 ;
        RECT 204.605 3021.545 205.925 3021.665 ;
        RECT 206.525 3021.845 207.495 3021.875 ;
        RECT 206.525 3021.675 207.325 3021.845 ;
        RECT 206.525 3021.545 207.495 3021.675 ;
        RECT 203.415 3021.165 204.435 3021.495 ;
        RECT 204.605 3021.385 204.775 3021.545 ;
        RECT 207.325 3021.385 207.495 3021.545 ;
        RECT 204.605 3020.985 204.775 3021.215 ;
        RECT 207.325 3020.985 207.495 3021.215 ;
      LAYER li1 ;
        RECT 207.495 3021.160 208.040 3024.580 ;
      LAYER li1 ;
        RECT 210.045 3020.985 210.215 3021.070 ;
        RECT 201.885 3020.925 202.780 3020.985 ;
        RECT 202.055 3020.755 202.780 3020.925 ;
        RECT 201.885 3020.695 202.780 3020.755 ;
        RECT 203.440 3020.925 205.940 3020.985 ;
        RECT 203.440 3020.755 204.605 3020.925 ;
        RECT 204.775 3020.755 205.940 3020.925 ;
        RECT 203.440 3020.695 205.940 3020.755 ;
        RECT 206.600 3020.925 208.220 3020.985 ;
        RECT 206.600 3020.755 207.325 3020.925 ;
        RECT 207.495 3020.755 208.220 3020.925 ;
        RECT 206.600 3020.695 208.220 3020.755 ;
        RECT 208.880 3020.925 210.215 3020.985 ;
        RECT 208.880 3020.755 210.045 3020.925 ;
        RECT 208.880 3020.695 210.215 3020.755 ;
        RECT 201.885 3020.465 202.055 3020.695 ;
        RECT 204.605 3020.465 204.775 3020.695 ;
        RECT 201.885 3020.135 202.055 3020.295 ;
        RECT 204.605 3020.135 204.775 3020.295 ;
        RECT 204.945 3020.185 205.965 3020.515 ;
        RECT 207.325 3020.465 207.495 3020.695 ;
        RECT 210.045 3020.610 210.215 3020.695 ;
        RECT 201.885 3020.005 202.855 3020.135 ;
        RECT 202.055 3019.835 202.855 3020.005 ;
        RECT 201.885 3019.805 202.855 3019.835 ;
        RECT 203.455 3020.015 204.775 3020.135 ;
        RECT 203.455 3020.005 205.575 3020.015 ;
        RECT 203.455 3019.835 204.605 3020.005 ;
        RECT 204.775 3019.845 205.575 3020.005 ;
        RECT 203.455 3019.805 204.775 3019.835 ;
        RECT 201.885 3019.545 202.055 3019.805 ;
        RECT 204.605 3019.545 204.775 3019.805 ;
        RECT 205.795 3019.675 205.965 3020.185 ;
        RECT 201.885 3019.295 202.055 3019.375 ;
        RECT 204.605 3019.295 204.775 3019.375 ;
        RECT 204.945 3019.345 205.965 3019.675 ;
        RECT 201.885 3019.085 202.535 3019.295 ;
        RECT 203.805 3019.175 204.775 3019.295 ;
        RECT 205.795 3019.190 205.965 3019.345 ;
        RECT 206.505 3020.265 207.155 3020.435 ;
        RECT 206.505 3019.595 206.675 3020.265 ;
        RECT 207.325 3020.095 207.495 3020.295 ;
        RECT 206.845 3020.005 207.495 3020.095 ;
        RECT 206.845 3019.835 207.325 3020.005 ;
        RECT 206.845 3019.765 207.495 3019.835 ;
        RECT 206.505 3019.425 207.150 3019.595 ;
        RECT 207.325 3019.545 207.495 3019.765 ;
        RECT 206.505 3019.190 206.675 3019.425 ;
        RECT 207.325 3019.255 207.495 3019.375 ;
        RECT 202.055 3018.965 202.535 3019.085 ;
        RECT 201.885 3018.625 202.055 3018.915 ;
        RECT 201.885 3018.165 202.535 3018.455 ;
        RECT 202.055 3018.125 202.535 3018.165 ;
        RECT 201.885 3017.705 202.055 3017.995 ;
        RECT 202.055 3017.535 202.535 3017.615 ;
        RECT 201.885 3017.285 202.535 3017.535 ;
        RECT 201.885 3017.245 202.055 3017.285 ;
        RECT 201.885 3016.785 202.055 3017.075 ;
        RECT 202.055 3016.615 202.535 3016.775 ;
        RECT 203.045 3016.685 203.215 3019.135 ;
        RECT 203.805 3019.085 205.575 3019.175 ;
        RECT 203.805 3018.965 204.605 3019.085 ;
        RECT 204.775 3019.005 205.575 3019.085 ;
        RECT 205.795 3019.015 206.675 3019.190 ;
        RECT 206.845 3019.085 207.495 3019.255 ;
        RECT 204.605 3018.625 204.775 3018.915 ;
      LAYER li1 ;
        RECT 204.945 3018.585 205.965 3018.755 ;
      LAYER li1 ;
        RECT 203.805 3018.415 204.775 3018.455 ;
        RECT 203.805 3018.165 205.575 3018.415 ;
        RECT 203.805 3018.125 204.605 3018.165 ;
        RECT 204.775 3018.085 205.575 3018.165 ;
        RECT 204.605 3017.705 204.775 3017.995 ;
      LAYER li1 ;
        RECT 205.795 3017.915 205.965 3018.585 ;
        RECT 204.945 3017.745 205.965 3017.915 ;
      LAYER li1 ;
        RECT 203.805 3017.535 204.605 3017.615 ;
        RECT 204.775 3017.535 205.575 3017.575 ;
        RECT 203.805 3017.285 205.575 3017.535 ;
        RECT 204.605 3017.245 205.575 3017.285 ;
      LAYER li1 ;
        RECT 205.795 3017.075 205.965 3017.745 ;
      LAYER li1 ;
        RECT 204.605 3016.785 204.775 3017.075 ;
      LAYER li1 ;
        RECT 204.945 3016.905 205.965 3017.075 ;
      LAYER li1 ;
        RECT 201.885 3016.445 202.535 3016.615 ;
        RECT 202.705 3016.510 203.585 3016.685 ;
        RECT 203.805 3016.615 204.605 3016.695 ;
        RECT 204.775 3016.615 205.575 3016.735 ;
        RECT 203.805 3016.525 205.575 3016.615 ;
        RECT 201.885 3016.325 202.055 3016.445 ;
        RECT 202.705 3016.275 202.875 3016.510 ;
        RECT 203.415 3016.355 203.585 3016.510 ;
        RECT 204.605 3016.405 205.575 3016.525 ;
        RECT 201.885 3015.935 202.055 3016.155 ;
        RECT 202.230 3016.105 202.875 3016.275 ;
        RECT 201.885 3015.865 202.535 3015.935 ;
        RECT 202.055 3015.695 202.535 3015.865 ;
        RECT 201.885 3015.605 202.535 3015.695 ;
        RECT 201.885 3015.405 202.055 3015.605 ;
        RECT 202.705 3015.435 202.875 3016.105 ;
        RECT 202.225 3015.265 202.875 3015.435 ;
        RECT 201.885 3015.005 202.055 3015.235 ;
      LAYER li1 ;
        RECT 203.045 3015.230 203.245 3016.330 ;
      LAYER li1 ;
        RECT 203.415 3016.025 204.435 3016.355 ;
        RECT 204.605 3016.325 204.775 3016.405 ;
      LAYER li1 ;
        RECT 205.795 3016.320 205.965 3016.905 ;
      LAYER li1 ;
        RECT 206.165 3016.565 206.335 3019.015 ;
        RECT 206.845 3018.925 207.325 3019.085 ;
      LAYER li1 ;
        RECT 207.495 3018.940 208.040 3020.525 ;
        RECT 206.505 3018.585 207.155 3018.755 ;
      LAYER li1 ;
        RECT 207.325 3018.625 207.495 3018.915 ;
      LAYER li1 ;
        RECT 207.495 3018.600 208.870 3018.940 ;
        RECT 206.505 3017.915 206.675 3018.585 ;
      LAYER li1 ;
        RECT 207.325 3018.415 207.495 3018.455 ;
        RECT 206.845 3018.165 207.495 3018.415 ;
        RECT 206.845 3018.085 207.325 3018.165 ;
      LAYER li1 ;
        RECT 206.505 3017.745 207.155 3017.915 ;
        RECT 206.505 3017.075 206.675 3017.745 ;
      LAYER li1 ;
        RECT 207.325 3017.705 207.495 3017.995 ;
        RECT 206.845 3017.535 207.325 3017.575 ;
        RECT 206.845 3017.245 207.495 3017.535 ;
      LAYER li1 ;
        RECT 206.505 3016.905 207.155 3017.075 ;
        RECT 206.505 3016.320 206.675 3016.905 ;
      LAYER li1 ;
        RECT 207.325 3016.785 207.495 3017.075 ;
        RECT 206.845 3016.615 207.325 3016.735 ;
        RECT 206.845 3016.405 207.495 3016.615 ;
        RECT 207.325 3016.325 207.495 3016.405 ;
      LAYER li1 ;
        RECT 205.795 3016.235 206.675 3016.320 ;
      LAYER li1 ;
        RECT 203.415 3015.515 203.585 3016.025 ;
        RECT 204.605 3015.895 204.775 3016.155 ;
      LAYER li1 ;
        RECT 204.945 3016.065 207.155 3016.235 ;
      LAYER li1 ;
        RECT 207.325 3015.895 207.495 3016.155 ;
        RECT 204.605 3015.865 205.925 3015.895 ;
        RECT 203.805 3015.695 204.605 3015.855 ;
        RECT 204.775 3015.695 205.925 3015.865 ;
        RECT 203.805 3015.685 205.925 3015.695 ;
        RECT 204.605 3015.565 205.925 3015.685 ;
        RECT 206.525 3015.865 207.495 3015.895 ;
        RECT 206.525 3015.695 207.325 3015.865 ;
        RECT 206.525 3015.565 207.495 3015.695 ;
        RECT 203.415 3015.185 204.435 3015.515 ;
        RECT 204.605 3015.405 204.775 3015.565 ;
        RECT 207.325 3015.405 207.495 3015.565 ;
        RECT 204.605 3015.005 204.775 3015.235 ;
        RECT 207.325 3015.005 207.495 3015.235 ;
      LAYER li1 ;
        RECT 207.495 3015.180 208.040 3018.600 ;
      LAYER li1 ;
        RECT 210.045 3015.005 210.215 3015.090 ;
        RECT 201.885 3014.945 202.780 3015.005 ;
        RECT 202.055 3014.775 202.780 3014.945 ;
        RECT 201.885 3014.715 202.780 3014.775 ;
        RECT 203.440 3014.945 205.940 3015.005 ;
        RECT 203.440 3014.775 204.605 3014.945 ;
        RECT 204.775 3014.775 205.940 3014.945 ;
        RECT 203.440 3014.715 205.940 3014.775 ;
        RECT 206.600 3014.945 208.220 3015.005 ;
        RECT 206.600 3014.775 207.325 3014.945 ;
        RECT 207.495 3014.775 208.220 3014.945 ;
        RECT 206.600 3014.715 208.220 3014.775 ;
        RECT 208.880 3014.945 210.215 3015.005 ;
        RECT 208.880 3014.775 210.045 3014.945 ;
        RECT 208.880 3014.715 210.215 3014.775 ;
        RECT 201.885 3014.485 202.055 3014.715 ;
        RECT 204.605 3014.485 204.775 3014.715 ;
        RECT 201.885 3014.155 202.055 3014.315 ;
        RECT 204.605 3014.155 204.775 3014.315 ;
        RECT 204.945 3014.205 205.965 3014.535 ;
        RECT 207.325 3014.485 207.495 3014.715 ;
        RECT 210.045 3014.630 210.215 3014.715 ;
        RECT 201.885 3014.025 202.855 3014.155 ;
        RECT 202.055 3013.855 202.855 3014.025 ;
        RECT 201.885 3013.825 202.855 3013.855 ;
        RECT 203.455 3014.035 204.775 3014.155 ;
        RECT 203.455 3014.025 205.575 3014.035 ;
        RECT 203.455 3013.855 204.605 3014.025 ;
        RECT 204.775 3013.865 205.575 3014.025 ;
        RECT 203.455 3013.825 204.775 3013.855 ;
        RECT 201.885 3013.565 202.055 3013.825 ;
        RECT 204.605 3013.565 204.775 3013.825 ;
        RECT 205.795 3013.695 205.965 3014.205 ;
        RECT 201.885 3013.315 202.055 3013.395 ;
        RECT 204.605 3013.315 204.775 3013.395 ;
        RECT 204.945 3013.365 205.965 3013.695 ;
        RECT 201.885 3013.105 202.535 3013.315 ;
        RECT 203.805 3013.195 204.775 3013.315 ;
        RECT 205.795 3013.210 205.965 3013.365 ;
        RECT 206.505 3014.285 207.155 3014.455 ;
        RECT 206.505 3013.615 206.675 3014.285 ;
        RECT 207.325 3014.115 207.495 3014.315 ;
        RECT 206.845 3014.025 207.495 3014.115 ;
        RECT 206.845 3013.855 207.325 3014.025 ;
        RECT 206.845 3013.785 207.495 3013.855 ;
        RECT 206.505 3013.445 207.150 3013.615 ;
        RECT 207.325 3013.565 207.495 3013.785 ;
        RECT 206.505 3013.210 206.675 3013.445 ;
        RECT 207.325 3013.275 207.495 3013.395 ;
        RECT 202.055 3012.985 202.535 3013.105 ;
        RECT 201.885 3012.645 202.055 3012.935 ;
        RECT 201.885 3012.185 202.535 3012.475 ;
        RECT 202.055 3012.145 202.535 3012.185 ;
        RECT 201.885 3011.725 202.055 3012.015 ;
        RECT 202.055 3011.555 202.535 3011.635 ;
        RECT 201.885 3011.305 202.535 3011.555 ;
        RECT 201.885 3011.265 202.055 3011.305 ;
        RECT 201.885 3010.805 202.055 3011.095 ;
        RECT 202.055 3010.635 202.535 3010.795 ;
        RECT 203.045 3010.705 203.215 3013.155 ;
        RECT 203.805 3013.105 205.575 3013.195 ;
        RECT 203.805 3012.985 204.605 3013.105 ;
        RECT 204.775 3013.025 205.575 3013.105 ;
        RECT 205.795 3013.035 206.675 3013.210 ;
        RECT 206.845 3013.105 207.495 3013.275 ;
        RECT 204.605 3012.645 204.775 3012.935 ;
      LAYER li1 ;
        RECT 204.945 3012.605 205.965 3012.775 ;
      LAYER li1 ;
        RECT 203.805 3012.435 204.775 3012.475 ;
        RECT 203.805 3012.185 205.575 3012.435 ;
        RECT 203.805 3012.145 204.605 3012.185 ;
        RECT 204.775 3012.105 205.575 3012.185 ;
        RECT 204.605 3011.725 204.775 3012.015 ;
      LAYER li1 ;
        RECT 205.795 3011.935 205.965 3012.605 ;
        RECT 204.945 3011.765 205.965 3011.935 ;
      LAYER li1 ;
        RECT 203.805 3011.555 204.605 3011.635 ;
        RECT 204.775 3011.555 205.575 3011.595 ;
        RECT 203.805 3011.305 205.575 3011.555 ;
        RECT 204.605 3011.265 205.575 3011.305 ;
      LAYER li1 ;
        RECT 205.795 3011.095 205.965 3011.765 ;
      LAYER li1 ;
        RECT 204.605 3010.805 204.775 3011.095 ;
      LAYER li1 ;
        RECT 204.945 3010.925 205.965 3011.095 ;
      LAYER li1 ;
        RECT 201.885 3010.465 202.535 3010.635 ;
        RECT 202.705 3010.530 203.585 3010.705 ;
        RECT 203.805 3010.635 204.605 3010.715 ;
        RECT 204.775 3010.635 205.575 3010.755 ;
        RECT 203.805 3010.545 205.575 3010.635 ;
        RECT 201.885 3010.345 202.055 3010.465 ;
        RECT 202.705 3010.295 202.875 3010.530 ;
        RECT 203.415 3010.375 203.585 3010.530 ;
        RECT 204.605 3010.425 205.575 3010.545 ;
        RECT 201.885 3009.955 202.055 3010.175 ;
        RECT 202.230 3010.125 202.875 3010.295 ;
        RECT 201.885 3009.885 202.535 3009.955 ;
        RECT 202.055 3009.715 202.535 3009.885 ;
        RECT 201.885 3009.625 202.535 3009.715 ;
        RECT 201.885 3009.425 202.055 3009.625 ;
        RECT 202.705 3009.455 202.875 3010.125 ;
        RECT 202.225 3009.285 202.875 3009.455 ;
        RECT 201.885 3009.025 202.055 3009.255 ;
      LAYER li1 ;
        RECT 203.045 3009.250 203.245 3010.350 ;
      LAYER li1 ;
        RECT 203.415 3010.045 204.435 3010.375 ;
        RECT 204.605 3010.345 204.775 3010.425 ;
      LAYER li1 ;
        RECT 205.795 3010.340 205.965 3010.925 ;
      LAYER li1 ;
        RECT 206.165 3010.585 206.335 3013.035 ;
        RECT 206.845 3012.945 207.325 3013.105 ;
      LAYER li1 ;
        RECT 207.495 3012.960 208.040 3014.545 ;
        RECT 206.505 3012.605 207.155 3012.775 ;
      LAYER li1 ;
        RECT 207.325 3012.645 207.495 3012.935 ;
      LAYER li1 ;
        RECT 207.495 3012.620 208.870 3012.960 ;
        RECT 206.505 3011.935 206.675 3012.605 ;
      LAYER li1 ;
        RECT 207.325 3012.435 207.495 3012.475 ;
        RECT 206.845 3012.185 207.495 3012.435 ;
        RECT 206.845 3012.105 207.325 3012.185 ;
      LAYER li1 ;
        RECT 206.505 3011.765 207.155 3011.935 ;
        RECT 206.505 3011.095 206.675 3011.765 ;
      LAYER li1 ;
        RECT 207.325 3011.725 207.495 3012.015 ;
        RECT 206.845 3011.555 207.325 3011.595 ;
        RECT 206.845 3011.265 207.495 3011.555 ;
      LAYER li1 ;
        RECT 206.505 3010.925 207.155 3011.095 ;
        RECT 206.505 3010.340 206.675 3010.925 ;
      LAYER li1 ;
        RECT 207.325 3010.805 207.495 3011.095 ;
        RECT 206.845 3010.635 207.325 3010.755 ;
        RECT 206.845 3010.425 207.495 3010.635 ;
        RECT 207.325 3010.345 207.495 3010.425 ;
      LAYER li1 ;
        RECT 205.795 3010.255 206.675 3010.340 ;
      LAYER li1 ;
        RECT 203.415 3009.535 203.585 3010.045 ;
        RECT 204.605 3009.915 204.775 3010.175 ;
      LAYER li1 ;
        RECT 204.945 3010.085 207.155 3010.255 ;
      LAYER li1 ;
        RECT 207.325 3009.915 207.495 3010.175 ;
        RECT 204.605 3009.885 205.925 3009.915 ;
        RECT 203.805 3009.715 204.605 3009.875 ;
        RECT 204.775 3009.715 205.925 3009.885 ;
        RECT 203.805 3009.705 205.925 3009.715 ;
        RECT 204.605 3009.585 205.925 3009.705 ;
        RECT 206.525 3009.885 207.495 3009.915 ;
        RECT 206.525 3009.715 207.325 3009.885 ;
        RECT 206.525 3009.585 207.495 3009.715 ;
        RECT 203.415 3009.205 204.435 3009.535 ;
        RECT 204.605 3009.425 204.775 3009.585 ;
        RECT 207.325 3009.425 207.495 3009.585 ;
        RECT 204.605 3009.025 204.775 3009.255 ;
        RECT 207.325 3009.025 207.495 3009.255 ;
      LAYER li1 ;
        RECT 207.495 3009.200 208.040 3012.620 ;
      LAYER li1 ;
        RECT 210.045 3009.025 210.215 3009.110 ;
        RECT 201.885 3008.965 202.780 3009.025 ;
        RECT 202.055 3008.795 202.780 3008.965 ;
        RECT 201.885 3008.735 202.780 3008.795 ;
        RECT 203.440 3008.965 205.940 3009.025 ;
        RECT 203.440 3008.795 204.605 3008.965 ;
        RECT 204.775 3008.795 205.940 3008.965 ;
        RECT 203.440 3008.735 205.940 3008.795 ;
        RECT 206.600 3008.965 208.220 3009.025 ;
        RECT 206.600 3008.795 207.325 3008.965 ;
        RECT 207.495 3008.795 208.220 3008.965 ;
        RECT 206.600 3008.735 208.220 3008.795 ;
        RECT 208.880 3008.965 210.215 3009.025 ;
        RECT 208.880 3008.795 210.045 3008.965 ;
        RECT 208.880 3008.735 210.215 3008.795 ;
        RECT 201.885 3008.505 202.055 3008.735 ;
        RECT 204.605 3008.505 204.775 3008.735 ;
        RECT 201.885 3008.175 202.055 3008.335 ;
        RECT 204.605 3008.175 204.775 3008.335 ;
        RECT 204.945 3008.225 205.965 3008.555 ;
        RECT 207.325 3008.505 207.495 3008.735 ;
        RECT 210.045 3008.650 210.215 3008.735 ;
        RECT 201.885 3008.045 202.855 3008.175 ;
        RECT 202.055 3007.875 202.855 3008.045 ;
        RECT 201.885 3007.845 202.855 3007.875 ;
        RECT 203.455 3008.055 204.775 3008.175 ;
        RECT 203.455 3008.045 205.575 3008.055 ;
        RECT 203.455 3007.875 204.605 3008.045 ;
        RECT 204.775 3007.885 205.575 3008.045 ;
        RECT 203.455 3007.845 204.775 3007.875 ;
        RECT 201.885 3007.585 202.055 3007.845 ;
        RECT 204.605 3007.585 204.775 3007.845 ;
        RECT 205.795 3007.715 205.965 3008.225 ;
        RECT 201.885 3007.335 202.055 3007.415 ;
        RECT 204.605 3007.335 204.775 3007.415 ;
        RECT 204.945 3007.385 205.965 3007.715 ;
        RECT 201.885 3007.125 202.535 3007.335 ;
        RECT 203.805 3007.215 204.775 3007.335 ;
        RECT 205.795 3007.230 205.965 3007.385 ;
        RECT 206.505 3008.305 207.155 3008.475 ;
        RECT 206.505 3007.635 206.675 3008.305 ;
        RECT 207.325 3008.135 207.495 3008.335 ;
        RECT 206.845 3008.045 207.495 3008.135 ;
        RECT 206.845 3007.875 207.325 3008.045 ;
        RECT 206.845 3007.805 207.495 3007.875 ;
        RECT 206.505 3007.465 207.150 3007.635 ;
        RECT 207.325 3007.585 207.495 3007.805 ;
        RECT 206.505 3007.230 206.675 3007.465 ;
        RECT 207.325 3007.295 207.495 3007.415 ;
        RECT 202.055 3007.005 202.535 3007.125 ;
        RECT 201.885 3006.665 202.055 3006.955 ;
        RECT 201.885 3006.205 202.535 3006.495 ;
        RECT 202.055 3006.165 202.535 3006.205 ;
        RECT 201.885 3005.745 202.055 3006.035 ;
        RECT 202.055 3005.575 202.535 3005.655 ;
        RECT 201.885 3005.325 202.535 3005.575 ;
        RECT 201.885 3005.285 202.055 3005.325 ;
        RECT 201.885 3004.825 202.055 3005.115 ;
        RECT 202.055 3004.655 202.535 3004.815 ;
        RECT 203.045 3004.725 203.215 3007.175 ;
        RECT 203.805 3007.125 205.575 3007.215 ;
        RECT 203.805 3007.005 204.605 3007.125 ;
        RECT 204.775 3007.045 205.575 3007.125 ;
        RECT 205.795 3007.055 206.675 3007.230 ;
        RECT 206.845 3007.125 207.495 3007.295 ;
        RECT 204.605 3006.665 204.775 3006.955 ;
      LAYER li1 ;
        RECT 204.945 3006.625 205.965 3006.795 ;
      LAYER li1 ;
        RECT 203.805 3006.455 204.775 3006.495 ;
        RECT 203.805 3006.205 205.575 3006.455 ;
        RECT 203.805 3006.165 204.605 3006.205 ;
        RECT 204.775 3006.125 205.575 3006.205 ;
        RECT 204.605 3005.745 204.775 3006.035 ;
      LAYER li1 ;
        RECT 205.795 3005.955 205.965 3006.625 ;
        RECT 204.945 3005.785 205.965 3005.955 ;
      LAYER li1 ;
        RECT 203.805 3005.575 204.605 3005.655 ;
        RECT 204.775 3005.575 205.575 3005.615 ;
        RECT 203.805 3005.325 205.575 3005.575 ;
        RECT 204.605 3005.285 205.575 3005.325 ;
      LAYER li1 ;
        RECT 205.795 3005.115 205.965 3005.785 ;
      LAYER li1 ;
        RECT 204.605 3004.825 204.775 3005.115 ;
      LAYER li1 ;
        RECT 204.945 3004.945 205.965 3005.115 ;
      LAYER li1 ;
        RECT 201.885 3004.485 202.535 3004.655 ;
        RECT 202.705 3004.550 203.585 3004.725 ;
        RECT 203.805 3004.655 204.605 3004.735 ;
        RECT 204.775 3004.655 205.575 3004.775 ;
        RECT 203.805 3004.565 205.575 3004.655 ;
        RECT 201.885 3004.365 202.055 3004.485 ;
        RECT 202.705 3004.315 202.875 3004.550 ;
        RECT 203.415 3004.395 203.585 3004.550 ;
        RECT 204.605 3004.445 205.575 3004.565 ;
        RECT 201.885 3003.975 202.055 3004.195 ;
        RECT 202.230 3004.145 202.875 3004.315 ;
        RECT 201.885 3003.905 202.535 3003.975 ;
        RECT 202.055 3003.735 202.535 3003.905 ;
        RECT 201.885 3003.645 202.535 3003.735 ;
        RECT 201.885 3003.445 202.055 3003.645 ;
        RECT 202.705 3003.475 202.875 3004.145 ;
        RECT 202.225 3003.305 202.875 3003.475 ;
        RECT 201.885 3003.045 202.055 3003.275 ;
      LAYER li1 ;
        RECT 203.045 3003.270 203.245 3004.370 ;
      LAYER li1 ;
        RECT 203.415 3004.065 204.435 3004.395 ;
        RECT 204.605 3004.365 204.775 3004.445 ;
      LAYER li1 ;
        RECT 205.795 3004.360 205.965 3004.945 ;
      LAYER li1 ;
        RECT 206.165 3004.605 206.335 3007.055 ;
        RECT 206.845 3006.965 207.325 3007.125 ;
      LAYER li1 ;
        RECT 207.495 3006.980 208.040 3008.565 ;
        RECT 206.505 3006.625 207.155 3006.795 ;
      LAYER li1 ;
        RECT 207.325 3006.665 207.495 3006.955 ;
      LAYER li1 ;
        RECT 207.495 3006.640 208.870 3006.980 ;
        RECT 206.505 3005.955 206.675 3006.625 ;
      LAYER li1 ;
        RECT 207.325 3006.455 207.495 3006.495 ;
        RECT 206.845 3006.205 207.495 3006.455 ;
        RECT 206.845 3006.125 207.325 3006.205 ;
      LAYER li1 ;
        RECT 206.505 3005.785 207.155 3005.955 ;
        RECT 206.505 3005.115 206.675 3005.785 ;
      LAYER li1 ;
        RECT 207.325 3005.745 207.495 3006.035 ;
        RECT 206.845 3005.575 207.325 3005.615 ;
        RECT 206.845 3005.285 207.495 3005.575 ;
      LAYER li1 ;
        RECT 206.505 3004.945 207.155 3005.115 ;
        RECT 206.505 3004.360 206.675 3004.945 ;
      LAYER li1 ;
        RECT 207.325 3004.825 207.495 3005.115 ;
        RECT 206.845 3004.655 207.325 3004.775 ;
        RECT 206.845 3004.445 207.495 3004.655 ;
        RECT 207.325 3004.365 207.495 3004.445 ;
      LAYER li1 ;
        RECT 205.795 3004.275 206.675 3004.360 ;
      LAYER li1 ;
        RECT 203.415 3003.555 203.585 3004.065 ;
        RECT 204.605 3003.935 204.775 3004.195 ;
      LAYER li1 ;
        RECT 204.945 3004.105 207.155 3004.275 ;
      LAYER li1 ;
        RECT 207.325 3003.935 207.495 3004.195 ;
        RECT 204.605 3003.905 205.925 3003.935 ;
        RECT 203.805 3003.735 204.605 3003.895 ;
        RECT 204.775 3003.735 205.925 3003.905 ;
        RECT 203.805 3003.725 205.925 3003.735 ;
        RECT 204.605 3003.605 205.925 3003.725 ;
        RECT 206.525 3003.905 207.495 3003.935 ;
        RECT 206.525 3003.735 207.325 3003.905 ;
        RECT 206.525 3003.605 207.495 3003.735 ;
        RECT 203.415 3003.225 204.435 3003.555 ;
        RECT 204.605 3003.445 204.775 3003.605 ;
        RECT 207.325 3003.445 207.495 3003.605 ;
        RECT 204.605 3003.045 204.775 3003.275 ;
        RECT 207.325 3003.045 207.495 3003.275 ;
      LAYER li1 ;
        RECT 207.495 3003.220 208.040 3006.640 ;
      LAYER li1 ;
        RECT 210.045 3003.045 210.215 3003.130 ;
        RECT 201.885 3002.985 202.780 3003.045 ;
        RECT 202.055 3002.815 202.780 3002.985 ;
        RECT 201.885 3002.755 202.780 3002.815 ;
        RECT 203.440 3002.985 205.940 3003.045 ;
        RECT 203.440 3002.815 204.605 3002.985 ;
        RECT 204.775 3002.815 205.940 3002.985 ;
        RECT 203.440 3002.755 205.940 3002.815 ;
        RECT 206.600 3002.985 208.220 3003.045 ;
        RECT 206.600 3002.815 207.325 3002.985 ;
        RECT 207.495 3002.815 208.220 3002.985 ;
        RECT 206.600 3002.755 208.220 3002.815 ;
        RECT 208.880 3002.985 210.215 3003.045 ;
        RECT 208.880 3002.815 210.045 3002.985 ;
        RECT 208.880 3002.755 210.215 3002.815 ;
        RECT 201.885 3002.525 202.055 3002.755 ;
        RECT 204.605 3002.525 204.775 3002.755 ;
        RECT 201.885 3002.195 202.055 3002.355 ;
        RECT 204.605 3002.195 204.775 3002.355 ;
        RECT 204.945 3002.245 205.965 3002.575 ;
        RECT 207.325 3002.525 207.495 3002.755 ;
        RECT 210.045 3002.670 210.215 3002.755 ;
        RECT 201.885 3002.065 202.855 3002.195 ;
        RECT 202.055 3001.895 202.855 3002.065 ;
        RECT 201.885 3001.865 202.855 3001.895 ;
        RECT 203.455 3002.075 204.775 3002.195 ;
        RECT 203.455 3002.065 205.575 3002.075 ;
        RECT 203.455 3001.895 204.605 3002.065 ;
        RECT 204.775 3001.905 205.575 3002.065 ;
        RECT 203.455 3001.865 204.775 3001.895 ;
        RECT 201.885 3001.605 202.055 3001.865 ;
        RECT 204.605 3001.605 204.775 3001.865 ;
        RECT 205.795 3001.735 205.965 3002.245 ;
        RECT 201.885 3001.355 202.055 3001.435 ;
        RECT 204.605 3001.355 204.775 3001.435 ;
        RECT 204.945 3001.405 205.965 3001.735 ;
        RECT 201.885 3001.145 202.535 3001.355 ;
        RECT 203.805 3001.235 204.775 3001.355 ;
        RECT 205.795 3001.250 205.965 3001.405 ;
        RECT 206.505 3002.325 207.155 3002.495 ;
        RECT 206.505 3001.655 206.675 3002.325 ;
        RECT 207.325 3002.155 207.495 3002.355 ;
        RECT 206.845 3002.065 207.495 3002.155 ;
        RECT 206.845 3001.895 207.325 3002.065 ;
        RECT 206.845 3001.825 207.495 3001.895 ;
        RECT 206.505 3001.485 207.150 3001.655 ;
        RECT 207.325 3001.605 207.495 3001.825 ;
        RECT 206.505 3001.250 206.675 3001.485 ;
        RECT 207.325 3001.315 207.495 3001.435 ;
        RECT 202.055 3001.025 202.535 3001.145 ;
        RECT 201.885 3000.685 202.055 3000.975 ;
        RECT 201.885 3000.225 202.535 3000.515 ;
        RECT 202.055 3000.185 202.535 3000.225 ;
        RECT 201.885 2999.765 202.055 3000.055 ;
        RECT 202.055 2999.595 202.535 2999.675 ;
        RECT 201.885 2999.345 202.535 2999.595 ;
        RECT 201.885 2999.305 202.055 2999.345 ;
        RECT 201.885 2998.845 202.055 2999.135 ;
        RECT 202.055 2998.675 202.535 2998.835 ;
        RECT 203.045 2998.745 203.215 3001.195 ;
        RECT 203.805 3001.145 205.575 3001.235 ;
        RECT 203.805 3001.025 204.605 3001.145 ;
        RECT 204.775 3001.065 205.575 3001.145 ;
        RECT 205.795 3001.075 206.675 3001.250 ;
        RECT 206.845 3001.145 207.495 3001.315 ;
        RECT 204.605 3000.685 204.775 3000.975 ;
      LAYER li1 ;
        RECT 204.945 3000.645 205.965 3000.815 ;
      LAYER li1 ;
        RECT 203.805 3000.475 204.775 3000.515 ;
        RECT 203.805 3000.225 205.575 3000.475 ;
        RECT 203.805 3000.185 204.605 3000.225 ;
        RECT 204.775 3000.145 205.575 3000.225 ;
        RECT 204.605 2999.765 204.775 3000.055 ;
      LAYER li1 ;
        RECT 205.795 2999.975 205.965 3000.645 ;
        RECT 204.945 2999.805 205.965 2999.975 ;
      LAYER li1 ;
        RECT 203.805 2999.595 204.605 2999.675 ;
        RECT 204.775 2999.595 205.575 2999.635 ;
        RECT 203.805 2999.345 205.575 2999.595 ;
        RECT 204.605 2999.305 205.575 2999.345 ;
      LAYER li1 ;
        RECT 205.795 2999.135 205.965 2999.805 ;
      LAYER li1 ;
        RECT 204.605 2998.845 204.775 2999.135 ;
      LAYER li1 ;
        RECT 204.945 2998.965 205.965 2999.135 ;
      LAYER li1 ;
        RECT 201.885 2998.505 202.535 2998.675 ;
        RECT 202.705 2998.570 203.585 2998.745 ;
        RECT 203.805 2998.675 204.605 2998.755 ;
        RECT 204.775 2998.675 205.575 2998.795 ;
        RECT 203.805 2998.585 205.575 2998.675 ;
        RECT 201.885 2998.385 202.055 2998.505 ;
        RECT 202.705 2998.335 202.875 2998.570 ;
        RECT 203.415 2998.415 203.585 2998.570 ;
        RECT 204.605 2998.465 205.575 2998.585 ;
        RECT 201.885 2997.995 202.055 2998.215 ;
        RECT 202.230 2998.165 202.875 2998.335 ;
        RECT 201.885 2997.925 202.535 2997.995 ;
        RECT 202.055 2997.755 202.535 2997.925 ;
        RECT 201.885 2997.665 202.535 2997.755 ;
        RECT 201.885 2997.465 202.055 2997.665 ;
        RECT 202.705 2997.495 202.875 2998.165 ;
        RECT 202.225 2997.325 202.875 2997.495 ;
        RECT 201.885 2997.065 202.055 2997.295 ;
      LAYER li1 ;
        RECT 203.045 2997.290 203.245 2998.390 ;
      LAYER li1 ;
        RECT 203.415 2998.085 204.435 2998.415 ;
        RECT 204.605 2998.385 204.775 2998.465 ;
      LAYER li1 ;
        RECT 205.795 2998.380 205.965 2998.965 ;
      LAYER li1 ;
        RECT 206.165 2998.625 206.335 3001.075 ;
        RECT 206.845 3000.985 207.325 3001.145 ;
      LAYER li1 ;
        RECT 207.495 3001.000 208.040 3002.585 ;
        RECT 206.505 3000.645 207.155 3000.815 ;
      LAYER li1 ;
        RECT 207.325 3000.685 207.495 3000.975 ;
      LAYER li1 ;
        RECT 207.495 3000.660 208.870 3001.000 ;
        RECT 206.505 2999.975 206.675 3000.645 ;
      LAYER li1 ;
        RECT 207.325 3000.475 207.495 3000.515 ;
        RECT 206.845 3000.225 207.495 3000.475 ;
        RECT 206.845 3000.145 207.325 3000.225 ;
      LAYER li1 ;
        RECT 206.505 2999.805 207.155 2999.975 ;
        RECT 206.505 2999.135 206.675 2999.805 ;
      LAYER li1 ;
        RECT 207.325 2999.765 207.495 3000.055 ;
        RECT 206.845 2999.595 207.325 2999.635 ;
        RECT 206.845 2999.305 207.495 2999.595 ;
      LAYER li1 ;
        RECT 206.505 2998.965 207.155 2999.135 ;
        RECT 206.505 2998.380 206.675 2998.965 ;
      LAYER li1 ;
        RECT 207.325 2998.845 207.495 2999.135 ;
        RECT 206.845 2998.675 207.325 2998.795 ;
        RECT 206.845 2998.465 207.495 2998.675 ;
        RECT 207.325 2998.385 207.495 2998.465 ;
      LAYER li1 ;
        RECT 205.795 2998.295 206.675 2998.380 ;
      LAYER li1 ;
        RECT 203.415 2997.575 203.585 2998.085 ;
        RECT 204.605 2997.955 204.775 2998.215 ;
      LAYER li1 ;
        RECT 204.945 2998.125 207.155 2998.295 ;
      LAYER li1 ;
        RECT 207.325 2997.955 207.495 2998.215 ;
        RECT 204.605 2997.925 205.925 2997.955 ;
        RECT 203.805 2997.755 204.605 2997.915 ;
        RECT 204.775 2997.755 205.925 2997.925 ;
        RECT 203.805 2997.745 205.925 2997.755 ;
        RECT 204.605 2997.625 205.925 2997.745 ;
        RECT 206.525 2997.925 207.495 2997.955 ;
        RECT 206.525 2997.755 207.325 2997.925 ;
        RECT 206.525 2997.625 207.495 2997.755 ;
        RECT 203.415 2997.245 204.435 2997.575 ;
        RECT 204.605 2997.465 204.775 2997.625 ;
        RECT 207.325 2997.465 207.495 2997.625 ;
        RECT 204.605 2997.065 204.775 2997.295 ;
        RECT 207.325 2997.065 207.495 2997.295 ;
      LAYER li1 ;
        RECT 207.495 2997.240 208.040 3000.660 ;
      LAYER li1 ;
        RECT 210.045 2997.065 210.215 2997.150 ;
        RECT 201.885 2997.005 202.780 2997.065 ;
        RECT 202.055 2996.835 202.780 2997.005 ;
        RECT 201.885 2996.775 202.780 2996.835 ;
        RECT 203.440 2997.005 205.940 2997.065 ;
        RECT 203.440 2996.835 204.605 2997.005 ;
        RECT 204.775 2996.835 205.940 2997.005 ;
        RECT 203.440 2996.775 205.940 2996.835 ;
        RECT 206.600 2997.005 208.220 2997.065 ;
        RECT 206.600 2996.835 207.325 2997.005 ;
        RECT 207.495 2996.835 208.220 2997.005 ;
        RECT 206.600 2996.775 208.220 2996.835 ;
        RECT 208.880 2997.005 210.215 2997.065 ;
        RECT 208.880 2996.835 210.045 2997.005 ;
        RECT 208.880 2996.775 210.215 2996.835 ;
        RECT 201.885 2996.545 202.055 2996.775 ;
        RECT 204.605 2996.545 204.775 2996.775 ;
        RECT 201.885 2996.215 202.055 2996.375 ;
        RECT 204.605 2996.215 204.775 2996.375 ;
        RECT 204.945 2996.265 205.965 2996.595 ;
        RECT 207.325 2996.545 207.495 2996.775 ;
        RECT 210.045 2996.690 210.215 2996.775 ;
        RECT 201.885 2996.085 202.855 2996.215 ;
        RECT 202.055 2995.915 202.855 2996.085 ;
        RECT 201.885 2995.885 202.855 2995.915 ;
        RECT 203.455 2996.095 204.775 2996.215 ;
        RECT 203.455 2996.085 205.575 2996.095 ;
        RECT 203.455 2995.915 204.605 2996.085 ;
        RECT 204.775 2995.925 205.575 2996.085 ;
        RECT 203.455 2995.885 204.775 2995.915 ;
        RECT 201.885 2995.625 202.055 2995.885 ;
        RECT 204.605 2995.625 204.775 2995.885 ;
        RECT 205.795 2995.755 205.965 2996.265 ;
        RECT 201.885 2995.375 202.055 2995.455 ;
        RECT 204.605 2995.375 204.775 2995.455 ;
        RECT 204.945 2995.425 205.965 2995.755 ;
        RECT 201.885 2995.165 202.535 2995.375 ;
        RECT 203.805 2995.255 204.775 2995.375 ;
        RECT 205.795 2995.270 205.965 2995.425 ;
        RECT 206.505 2996.345 207.155 2996.515 ;
        RECT 206.505 2995.675 206.675 2996.345 ;
        RECT 207.325 2996.175 207.495 2996.375 ;
        RECT 206.845 2996.085 207.495 2996.175 ;
        RECT 206.845 2995.915 207.325 2996.085 ;
        RECT 206.845 2995.845 207.495 2995.915 ;
        RECT 206.505 2995.505 207.150 2995.675 ;
        RECT 207.325 2995.625 207.495 2995.845 ;
        RECT 206.505 2995.270 206.675 2995.505 ;
        RECT 207.325 2995.335 207.495 2995.455 ;
        RECT 202.055 2995.045 202.535 2995.165 ;
        RECT 201.885 2994.705 202.055 2994.995 ;
        RECT 201.885 2994.245 202.535 2994.535 ;
        RECT 202.055 2994.205 202.535 2994.245 ;
        RECT 201.885 2993.785 202.055 2994.075 ;
        RECT 202.055 2993.615 202.535 2993.695 ;
        RECT 201.885 2993.365 202.535 2993.615 ;
        RECT 201.885 2993.325 202.055 2993.365 ;
        RECT 201.885 2992.865 202.055 2993.155 ;
        RECT 202.055 2992.695 202.535 2992.855 ;
        RECT 203.045 2992.765 203.215 2995.215 ;
        RECT 203.805 2995.165 205.575 2995.255 ;
        RECT 203.805 2995.045 204.605 2995.165 ;
        RECT 204.775 2995.085 205.575 2995.165 ;
        RECT 205.795 2995.095 206.675 2995.270 ;
        RECT 206.845 2995.165 207.495 2995.335 ;
        RECT 204.605 2994.705 204.775 2994.995 ;
      LAYER li1 ;
        RECT 204.945 2994.665 205.965 2994.835 ;
      LAYER li1 ;
        RECT 203.805 2994.495 204.775 2994.535 ;
        RECT 203.805 2994.245 205.575 2994.495 ;
        RECT 203.805 2994.205 204.605 2994.245 ;
        RECT 204.775 2994.165 205.575 2994.245 ;
        RECT 204.605 2993.785 204.775 2994.075 ;
      LAYER li1 ;
        RECT 205.795 2993.995 205.965 2994.665 ;
        RECT 204.945 2993.825 205.965 2993.995 ;
      LAYER li1 ;
        RECT 203.805 2993.615 204.605 2993.695 ;
        RECT 204.775 2993.615 205.575 2993.655 ;
        RECT 203.805 2993.365 205.575 2993.615 ;
        RECT 204.605 2993.325 205.575 2993.365 ;
      LAYER li1 ;
        RECT 205.795 2993.155 205.965 2993.825 ;
      LAYER li1 ;
        RECT 204.605 2992.865 204.775 2993.155 ;
      LAYER li1 ;
        RECT 204.945 2992.985 205.965 2993.155 ;
      LAYER li1 ;
        RECT 201.885 2992.525 202.535 2992.695 ;
        RECT 202.705 2992.590 203.585 2992.765 ;
        RECT 203.805 2992.695 204.605 2992.775 ;
        RECT 204.775 2992.695 205.575 2992.815 ;
        RECT 203.805 2992.605 205.575 2992.695 ;
        RECT 201.885 2992.405 202.055 2992.525 ;
        RECT 202.705 2992.355 202.875 2992.590 ;
        RECT 203.415 2992.435 203.585 2992.590 ;
        RECT 204.605 2992.485 205.575 2992.605 ;
        RECT 201.885 2992.015 202.055 2992.235 ;
        RECT 202.230 2992.185 202.875 2992.355 ;
        RECT 201.885 2991.945 202.535 2992.015 ;
        RECT 202.055 2991.775 202.535 2991.945 ;
        RECT 201.885 2991.685 202.535 2991.775 ;
        RECT 201.885 2991.485 202.055 2991.685 ;
        RECT 202.705 2991.515 202.875 2992.185 ;
        RECT 202.225 2991.345 202.875 2991.515 ;
        RECT 201.885 2991.085 202.055 2991.315 ;
      LAYER li1 ;
        RECT 203.045 2991.310 203.245 2992.410 ;
      LAYER li1 ;
        RECT 203.415 2992.105 204.435 2992.435 ;
        RECT 204.605 2992.405 204.775 2992.485 ;
      LAYER li1 ;
        RECT 205.795 2992.400 205.965 2992.985 ;
      LAYER li1 ;
        RECT 206.165 2992.645 206.335 2995.095 ;
        RECT 206.845 2995.005 207.325 2995.165 ;
      LAYER li1 ;
        RECT 207.495 2995.020 208.040 2996.605 ;
        RECT 206.505 2994.665 207.155 2994.835 ;
      LAYER li1 ;
        RECT 207.325 2994.705 207.495 2994.995 ;
      LAYER li1 ;
        RECT 207.495 2994.680 208.870 2995.020 ;
        RECT 206.505 2993.995 206.675 2994.665 ;
      LAYER li1 ;
        RECT 207.325 2994.495 207.495 2994.535 ;
        RECT 206.845 2994.245 207.495 2994.495 ;
        RECT 206.845 2994.165 207.325 2994.245 ;
      LAYER li1 ;
        RECT 206.505 2993.825 207.155 2993.995 ;
        RECT 206.505 2993.155 206.675 2993.825 ;
      LAYER li1 ;
        RECT 207.325 2993.785 207.495 2994.075 ;
        RECT 206.845 2993.615 207.325 2993.655 ;
        RECT 206.845 2993.325 207.495 2993.615 ;
      LAYER li1 ;
        RECT 206.505 2992.985 207.155 2993.155 ;
        RECT 206.505 2992.400 206.675 2992.985 ;
      LAYER li1 ;
        RECT 207.325 2992.865 207.495 2993.155 ;
        RECT 206.845 2992.695 207.325 2992.815 ;
        RECT 206.845 2992.485 207.495 2992.695 ;
        RECT 207.325 2992.405 207.495 2992.485 ;
      LAYER li1 ;
        RECT 205.795 2992.315 206.675 2992.400 ;
      LAYER li1 ;
        RECT 203.415 2991.595 203.585 2992.105 ;
        RECT 204.605 2991.975 204.775 2992.235 ;
      LAYER li1 ;
        RECT 204.945 2992.145 207.155 2992.315 ;
      LAYER li1 ;
        RECT 207.325 2991.975 207.495 2992.235 ;
        RECT 204.605 2991.945 205.925 2991.975 ;
        RECT 203.805 2991.775 204.605 2991.935 ;
        RECT 204.775 2991.775 205.925 2991.945 ;
        RECT 203.805 2991.765 205.925 2991.775 ;
        RECT 204.605 2991.645 205.925 2991.765 ;
        RECT 206.525 2991.945 207.495 2991.975 ;
        RECT 206.525 2991.775 207.325 2991.945 ;
        RECT 206.525 2991.645 207.495 2991.775 ;
        RECT 203.415 2991.265 204.435 2991.595 ;
        RECT 204.605 2991.485 204.775 2991.645 ;
        RECT 207.325 2991.485 207.495 2991.645 ;
        RECT 204.605 2991.085 204.775 2991.315 ;
        RECT 207.325 2991.085 207.495 2991.315 ;
      LAYER li1 ;
        RECT 207.495 2991.260 208.040 2994.680 ;
      LAYER li1 ;
        RECT 210.045 2991.085 210.215 2991.170 ;
        RECT 201.885 2991.025 202.780 2991.085 ;
        RECT 202.055 2990.855 202.780 2991.025 ;
        RECT 201.885 2990.795 202.780 2990.855 ;
        RECT 203.440 2991.025 205.940 2991.085 ;
        RECT 203.440 2990.855 204.605 2991.025 ;
        RECT 204.775 2990.855 205.940 2991.025 ;
        RECT 203.440 2990.795 205.940 2990.855 ;
        RECT 206.600 2991.025 208.220 2991.085 ;
        RECT 206.600 2990.855 207.325 2991.025 ;
        RECT 207.495 2990.855 208.220 2991.025 ;
        RECT 206.600 2990.795 208.220 2990.855 ;
        RECT 208.880 2991.025 210.215 2991.085 ;
        RECT 208.880 2990.855 210.045 2991.025 ;
        RECT 208.880 2990.795 210.215 2990.855 ;
        RECT 201.885 2990.565 202.055 2990.795 ;
        RECT 204.605 2990.565 204.775 2990.795 ;
        RECT 207.325 2990.710 207.495 2990.795 ;
        RECT 210.045 2990.710 210.215 2990.795 ;
        RECT 201.885 2990.235 202.055 2990.395 ;
        RECT 204.605 2990.235 204.775 2990.395 ;
        RECT 204.945 2990.285 205.965 2990.615 ;
        RECT 201.885 2990.105 202.855 2990.235 ;
        RECT 202.055 2989.935 202.855 2990.105 ;
        RECT 201.885 2989.905 202.855 2989.935 ;
        RECT 203.455 2990.115 204.775 2990.235 ;
        RECT 203.455 2990.105 205.575 2990.115 ;
        RECT 203.455 2989.935 204.605 2990.105 ;
        RECT 204.775 2989.945 205.575 2990.105 ;
        RECT 203.455 2989.905 204.775 2989.935 ;
        RECT 201.885 2989.645 202.055 2989.905 ;
        RECT 204.605 2989.645 204.775 2989.905 ;
        RECT 205.795 2989.775 205.965 2990.285 ;
        RECT 201.885 2989.395 202.055 2989.475 ;
        RECT 204.605 2989.395 204.775 2989.475 ;
        RECT 204.945 2989.445 205.965 2989.775 ;
        RECT 201.885 2989.185 202.535 2989.395 ;
        RECT 203.805 2989.275 204.775 2989.395 ;
        RECT 205.795 2989.290 205.965 2989.445 ;
        RECT 206.505 2990.365 207.155 2990.535 ;
        RECT 206.505 2989.695 206.675 2990.365 ;
        RECT 206.845 2989.865 207.325 2990.195 ;
        RECT 206.505 2989.525 207.150 2989.695 ;
        RECT 206.505 2989.290 206.675 2989.525 ;
        RECT 202.055 2989.065 202.535 2989.185 ;
        RECT 201.885 2988.725 202.055 2989.015 ;
        RECT 201.885 2988.265 202.535 2988.555 ;
        RECT 202.055 2988.225 202.535 2988.265 ;
        RECT 201.885 2987.805 202.055 2988.095 ;
        RECT 202.055 2987.635 202.535 2987.715 ;
        RECT 201.885 2987.385 202.535 2987.635 ;
        RECT 201.885 2987.345 202.055 2987.385 ;
        RECT 201.885 2986.885 202.055 2987.175 ;
        RECT 202.055 2986.715 202.535 2986.875 ;
        RECT 203.045 2986.785 203.215 2989.235 ;
        RECT 203.805 2989.185 205.575 2989.275 ;
        RECT 203.805 2989.065 204.605 2989.185 ;
        RECT 204.775 2989.105 205.575 2989.185 ;
        RECT 205.795 2989.115 206.675 2989.290 ;
        RECT 204.605 2988.725 204.775 2989.015 ;
      LAYER li1 ;
        RECT 204.945 2988.685 205.965 2988.855 ;
      LAYER li1 ;
        RECT 203.805 2988.515 204.775 2988.555 ;
        RECT 203.805 2988.265 205.575 2988.515 ;
        RECT 203.805 2988.225 204.605 2988.265 ;
        RECT 204.775 2988.185 205.575 2988.265 ;
        RECT 204.605 2987.805 204.775 2988.095 ;
      LAYER li1 ;
        RECT 205.795 2988.015 205.965 2988.685 ;
        RECT 204.945 2987.845 205.965 2988.015 ;
      LAYER li1 ;
        RECT 203.805 2987.635 204.605 2987.715 ;
        RECT 204.775 2987.635 205.575 2987.675 ;
        RECT 203.805 2987.385 205.575 2987.635 ;
        RECT 204.605 2987.345 205.575 2987.385 ;
      LAYER li1 ;
        RECT 205.795 2987.175 205.965 2987.845 ;
      LAYER li1 ;
        RECT 204.605 2986.885 204.775 2987.175 ;
      LAYER li1 ;
        RECT 204.945 2987.005 205.965 2987.175 ;
      LAYER li1 ;
        RECT 201.885 2986.545 202.535 2986.715 ;
        RECT 202.705 2986.610 203.585 2986.785 ;
        RECT 203.805 2986.715 204.605 2986.795 ;
        RECT 204.775 2986.715 205.575 2986.835 ;
        RECT 203.805 2986.625 205.575 2986.715 ;
        RECT 201.885 2986.425 202.055 2986.545 ;
        RECT 202.705 2986.375 202.875 2986.610 ;
        RECT 203.415 2986.455 203.585 2986.610 ;
        RECT 204.605 2986.505 205.575 2986.625 ;
        RECT 201.885 2986.035 202.055 2986.255 ;
        RECT 202.230 2986.205 202.875 2986.375 ;
        RECT 201.885 2985.965 202.535 2986.035 ;
        RECT 202.055 2985.795 202.535 2985.965 ;
        RECT 201.885 2985.705 202.535 2985.795 ;
        RECT 201.885 2985.505 202.055 2985.705 ;
        RECT 202.705 2985.535 202.875 2986.205 ;
        RECT 202.225 2985.365 202.875 2985.535 ;
        RECT 201.885 2985.105 202.055 2985.335 ;
      LAYER li1 ;
        RECT 203.045 2985.330 203.245 2986.430 ;
      LAYER li1 ;
        RECT 203.415 2986.125 204.435 2986.455 ;
        RECT 204.605 2986.425 204.775 2986.505 ;
      LAYER li1 ;
        RECT 205.795 2986.420 205.965 2987.005 ;
      LAYER li1 ;
        RECT 206.165 2986.665 206.335 2989.115 ;
        RECT 206.845 2989.025 207.325 2989.355 ;
      LAYER li1 ;
        RECT 206.505 2988.685 207.155 2988.855 ;
        RECT 206.505 2988.015 206.675 2988.685 ;
      LAYER li1 ;
        RECT 206.845 2988.185 207.325 2988.515 ;
      LAYER li1 ;
        RECT 206.505 2987.845 207.155 2988.015 ;
        RECT 206.505 2987.175 206.675 2987.845 ;
      LAYER li1 ;
        RECT 206.845 2987.345 207.325 2987.675 ;
      LAYER li1 ;
        RECT 206.505 2987.005 207.155 2987.175 ;
        RECT 206.505 2986.420 206.675 2987.005 ;
      LAYER li1 ;
        RECT 206.845 2986.505 207.325 2986.835 ;
      LAYER li1 ;
        RECT 205.795 2986.335 206.675 2986.420 ;
      LAYER li1 ;
        RECT 203.415 2985.615 203.585 2986.125 ;
        RECT 204.605 2985.995 204.775 2986.255 ;
      LAYER li1 ;
        RECT 204.945 2986.165 207.155 2986.335 ;
      LAYER li1 ;
        RECT 204.605 2985.965 205.925 2985.995 ;
        RECT 203.805 2985.795 204.605 2985.955 ;
        RECT 204.775 2985.795 205.925 2985.965 ;
        RECT 203.805 2985.785 205.925 2985.795 ;
        RECT 204.605 2985.665 205.925 2985.785 ;
        RECT 206.525 2985.665 207.325 2985.995 ;
        RECT 203.415 2985.285 204.435 2985.615 ;
        RECT 204.605 2985.505 204.775 2985.665 ;
        RECT 204.605 2985.105 204.775 2985.335 ;
        RECT 207.325 2985.105 207.495 2985.190 ;
        RECT 210.045 2985.105 210.215 2985.190 ;
        RECT 201.885 2985.045 202.780 2985.105 ;
        RECT 202.055 2984.875 202.780 2985.045 ;
        RECT 201.885 2984.815 202.780 2984.875 ;
        RECT 203.440 2985.045 205.940 2985.105 ;
        RECT 203.440 2984.875 204.605 2985.045 ;
        RECT 204.775 2984.875 205.940 2985.045 ;
        RECT 203.440 2984.815 205.940 2984.875 ;
        RECT 206.600 2985.045 208.220 2985.105 ;
        RECT 206.600 2984.875 207.325 2985.045 ;
        RECT 207.495 2984.875 208.220 2985.045 ;
        RECT 206.600 2984.815 208.220 2984.875 ;
        RECT 208.880 2985.045 210.215 2985.105 ;
        RECT 208.880 2984.875 210.045 2985.045 ;
        RECT 208.880 2984.815 210.215 2984.875 ;
        RECT 201.885 2984.730 202.055 2984.815 ;
        RECT 204.605 2984.730 204.775 2984.815 ;
        RECT 207.325 2984.730 207.495 2984.815 ;
        RECT 210.045 2984.730 210.215 2984.815 ;
        RECT 3377.780 2268.195 3377.950 2268.280 ;
        RECT 3380.500 2268.195 3380.670 2268.280 ;
        RECT 3383.220 2268.195 3383.390 2268.280 ;
        RECT 3385.940 2268.195 3386.110 2268.280 ;
        RECT 3377.780 2268.135 3379.115 2268.195 ;
        RECT 3377.950 2267.965 3379.115 2268.135 ;
        RECT 3377.780 2267.905 3379.115 2267.965 ;
        RECT 3379.775 2268.135 3381.395 2268.195 ;
        RECT 3379.775 2267.965 3380.500 2268.135 ;
        RECT 3380.670 2267.965 3381.395 2268.135 ;
        RECT 3379.775 2267.905 3381.395 2267.965 ;
        RECT 3377.780 2267.820 3377.950 2267.905 ;
      LAYER li1 ;
        RECT 3379.955 2266.150 3380.500 2267.735 ;
      LAYER li1 ;
        RECT 3380.500 2267.675 3380.670 2267.905 ;
        RECT 3380.500 2267.305 3380.670 2267.505 ;
        RECT 3380.840 2267.475 3381.490 2267.645 ;
        RECT 3380.500 2267.215 3381.150 2267.305 ;
        RECT 3380.670 2267.045 3381.150 2267.215 ;
        RECT 3380.500 2266.975 3381.150 2267.045 ;
        RECT 3380.500 2266.755 3380.670 2266.975 ;
        RECT 3381.320 2266.805 3381.490 2267.475 ;
        RECT 3380.845 2266.635 3381.490 2266.805 ;
        RECT 3380.500 2266.465 3380.670 2266.585 ;
        RECT 3380.500 2266.295 3381.150 2266.465 ;
      LAYER li1 ;
        RECT 3379.125 2265.810 3380.500 2266.150 ;
      LAYER li1 ;
        RECT 3380.670 2266.135 3381.150 2266.295 ;
        RECT 3381.320 2266.400 3381.490 2266.635 ;
      LAYER li1 ;
        RECT 3381.660 2266.580 3381.860 2268.170 ;
      LAYER li1 ;
        RECT 3382.055 2268.135 3384.555 2268.195 ;
        RECT 3382.055 2267.965 3383.220 2268.135 ;
        RECT 3383.390 2267.965 3384.555 2268.135 ;
        RECT 3382.055 2267.905 3384.555 2267.965 ;
        RECT 3385.215 2268.135 3386.110 2268.195 ;
        RECT 3385.215 2267.965 3385.940 2268.135 ;
        RECT 3385.215 2267.905 3386.110 2267.965 ;
        RECT 3382.030 2267.395 3383.050 2267.725 ;
        RECT 3383.220 2267.675 3383.390 2267.905 ;
        RECT 3385.940 2267.675 3386.110 2267.905 ;
        RECT 3382.030 2266.885 3382.200 2267.395 ;
        RECT 3383.220 2267.345 3383.390 2267.505 ;
        RECT 3385.940 2267.345 3386.110 2267.505 ;
        RECT 3383.220 2267.225 3384.540 2267.345 ;
        RECT 3382.420 2267.215 3384.540 2267.225 ;
        RECT 3382.420 2267.055 3383.220 2267.215 ;
        RECT 3383.390 2267.045 3384.540 2267.215 ;
        RECT 3383.220 2267.015 3384.540 2267.045 ;
        RECT 3385.140 2267.215 3386.110 2267.345 ;
        RECT 3385.140 2267.045 3385.940 2267.215 ;
        RECT 3385.140 2267.015 3386.110 2267.045 ;
        RECT 3382.030 2266.555 3383.050 2266.885 ;
        RECT 3383.220 2266.755 3383.390 2267.015 ;
      LAYER li1 ;
        RECT 3383.560 2266.675 3385.770 2266.845 ;
      LAYER li1 ;
        RECT 3385.940 2266.755 3386.110 2267.015 ;
      LAYER li1 ;
        RECT 3384.410 2266.590 3385.290 2266.675 ;
      LAYER li1 ;
        RECT 3382.030 2266.400 3382.200 2266.555 ;
        RECT 3381.320 2266.225 3382.200 2266.400 ;
        RECT 3383.220 2266.505 3383.390 2266.585 ;
        RECT 3383.220 2266.385 3384.190 2266.505 ;
        RECT 3382.420 2266.295 3384.190 2266.385 ;
        RECT 3380.500 2265.835 3380.670 2266.125 ;
      LAYER li1 ;
        RECT 3379.955 2262.390 3380.500 2265.810 ;
      LAYER li1 ;
        RECT 3380.500 2265.625 3380.670 2265.665 ;
        RECT 3380.500 2265.375 3381.150 2265.625 ;
        RECT 3380.670 2265.295 3381.150 2265.375 ;
        RECT 3380.500 2264.915 3380.670 2265.205 ;
        RECT 3380.670 2264.745 3381.150 2264.785 ;
        RECT 3380.500 2264.455 3381.150 2264.745 ;
        RECT 3380.500 2263.995 3380.670 2264.285 ;
        RECT 3380.670 2263.825 3381.150 2263.945 ;
        RECT 3380.500 2263.615 3381.150 2263.825 ;
        RECT 3381.660 2263.775 3381.830 2266.225 ;
        RECT 3382.420 2266.215 3383.220 2266.295 ;
        RECT 3383.390 2266.175 3384.190 2266.295 ;
        RECT 3383.220 2265.835 3383.390 2266.125 ;
      LAYER li1 ;
        RECT 3384.410 2266.005 3384.580 2266.590 ;
        RECT 3383.560 2265.835 3384.580 2266.005 ;
      LAYER li1 ;
        RECT 3383.220 2265.625 3384.190 2265.665 ;
        RECT 3382.420 2265.375 3384.190 2265.625 ;
        RECT 3382.420 2265.295 3383.220 2265.375 ;
        RECT 3383.390 2265.335 3384.190 2265.375 ;
        RECT 3383.220 2264.915 3383.390 2265.205 ;
      LAYER li1 ;
        RECT 3384.410 2265.165 3384.580 2265.835 ;
        RECT 3383.560 2264.995 3384.580 2265.165 ;
      LAYER li1 ;
        RECT 3382.420 2264.745 3383.220 2264.785 ;
        RECT 3383.390 2264.745 3384.190 2264.825 ;
        RECT 3382.420 2264.495 3384.190 2264.745 ;
        RECT 3382.420 2264.455 3383.390 2264.495 ;
      LAYER li1 ;
        RECT 3384.410 2264.325 3384.580 2264.995 ;
      LAYER li1 ;
        RECT 3383.220 2263.995 3383.390 2264.285 ;
      LAYER li1 ;
        RECT 3383.560 2264.155 3384.580 2264.325 ;
      LAYER li1 ;
        RECT 3382.420 2263.825 3383.220 2263.945 ;
        RECT 3383.390 2263.825 3384.190 2263.905 ;
        RECT 3384.780 2263.895 3384.950 2266.345 ;
      LAYER li1 ;
        RECT 3385.120 2266.005 3385.290 2266.590 ;
      LAYER li1 ;
        RECT 3385.940 2266.505 3386.110 2266.585 ;
        RECT 3385.460 2266.295 3386.110 2266.505 ;
        RECT 3385.460 2266.175 3385.940 2266.295 ;
      LAYER li1 ;
        RECT 3385.120 2265.835 3385.770 2266.005 ;
      LAYER li1 ;
        RECT 3385.940 2265.835 3386.110 2266.125 ;
      LAYER li1 ;
        RECT 3385.120 2265.165 3385.290 2265.835 ;
      LAYER li1 ;
        RECT 3385.460 2265.375 3386.110 2265.665 ;
        RECT 3385.460 2265.335 3385.940 2265.375 ;
      LAYER li1 ;
        RECT 3385.120 2264.995 3385.770 2265.165 ;
        RECT 3385.120 2264.325 3385.290 2264.995 ;
      LAYER li1 ;
        RECT 3385.940 2264.915 3386.110 2265.205 ;
        RECT 3385.460 2264.745 3385.940 2264.825 ;
        RECT 3385.460 2264.495 3386.110 2264.745 ;
        RECT 3385.940 2264.455 3386.110 2264.495 ;
      LAYER li1 ;
        RECT 3385.120 2264.155 3385.770 2264.325 ;
      LAYER li1 ;
        RECT 3385.940 2263.995 3386.110 2264.285 ;
        RECT 3382.420 2263.735 3384.190 2263.825 ;
        RECT 3382.420 2263.615 3383.390 2263.735 ;
        RECT 3380.500 2263.535 3380.670 2263.615 ;
        RECT 3383.220 2263.535 3383.390 2263.615 ;
        RECT 3384.410 2263.720 3385.290 2263.895 ;
        RECT 3384.410 2263.565 3384.580 2263.720 ;
        RECT 3380.500 2263.105 3380.670 2263.365 ;
        RECT 3383.220 2263.105 3383.390 2263.365 ;
        RECT 3383.560 2263.235 3384.580 2263.565 ;
        RECT 3380.500 2263.075 3381.470 2263.105 ;
        RECT 3380.670 2262.905 3381.470 2263.075 ;
        RECT 3380.500 2262.775 3381.470 2262.905 ;
        RECT 3382.070 2263.075 3383.390 2263.105 ;
        RECT 3382.070 2262.905 3383.220 2263.075 ;
        RECT 3383.390 2262.905 3384.190 2263.065 ;
        RECT 3382.070 2262.895 3384.190 2262.905 ;
        RECT 3382.070 2262.775 3383.390 2262.895 ;
        RECT 3380.500 2262.615 3380.670 2262.775 ;
        RECT 3383.220 2262.615 3383.390 2262.775 ;
        RECT 3384.410 2262.725 3384.580 2263.235 ;
        RECT 3377.780 2262.215 3377.950 2262.300 ;
        RECT 3380.500 2262.215 3380.670 2262.445 ;
        RECT 3383.220 2262.215 3383.390 2262.445 ;
        RECT 3383.560 2262.395 3384.580 2262.725 ;
        RECT 3385.120 2263.485 3385.290 2263.720 ;
        RECT 3385.460 2263.825 3385.940 2263.985 ;
        RECT 3385.460 2263.655 3386.110 2263.825 ;
        RECT 3385.940 2263.535 3386.110 2263.655 ;
        RECT 3385.120 2263.315 3385.765 2263.485 ;
        RECT 3385.120 2262.645 3385.290 2263.315 ;
        RECT 3385.940 2263.145 3386.110 2263.365 ;
        RECT 3385.460 2263.075 3386.110 2263.145 ;
        RECT 3385.460 2262.905 3385.940 2263.075 ;
        RECT 3385.460 2262.815 3386.110 2262.905 ;
        RECT 3385.120 2262.475 3385.770 2262.645 ;
        RECT 3385.940 2262.615 3386.110 2262.815 ;
        RECT 3385.940 2262.215 3386.110 2262.445 ;
        RECT 3377.780 2262.155 3379.115 2262.215 ;
        RECT 3377.950 2261.985 3379.115 2262.155 ;
        RECT 3377.780 2261.925 3379.115 2261.985 ;
        RECT 3379.775 2262.155 3381.395 2262.215 ;
        RECT 3379.775 2261.985 3380.500 2262.155 ;
        RECT 3380.670 2261.985 3381.395 2262.155 ;
        RECT 3379.775 2261.925 3381.395 2261.985 ;
        RECT 3377.780 2261.840 3377.950 2261.925 ;
      LAYER li1 ;
        RECT 3379.955 2260.170 3380.500 2261.755 ;
      LAYER li1 ;
        RECT 3380.500 2261.695 3380.670 2261.925 ;
        RECT 3380.500 2261.325 3380.670 2261.525 ;
        RECT 3380.840 2261.495 3381.490 2261.665 ;
        RECT 3380.500 2261.235 3381.150 2261.325 ;
        RECT 3380.670 2261.065 3381.150 2261.235 ;
        RECT 3380.500 2260.995 3381.150 2261.065 ;
        RECT 3380.500 2260.775 3380.670 2260.995 ;
        RECT 3381.320 2260.825 3381.490 2261.495 ;
        RECT 3380.845 2260.655 3381.490 2260.825 ;
        RECT 3380.500 2260.485 3380.670 2260.605 ;
        RECT 3380.500 2260.315 3381.150 2260.485 ;
      LAYER li1 ;
        RECT 3379.125 2259.830 3380.500 2260.170 ;
      LAYER li1 ;
        RECT 3380.670 2260.155 3381.150 2260.315 ;
        RECT 3381.320 2260.420 3381.490 2260.655 ;
      LAYER li1 ;
        RECT 3381.660 2260.600 3381.860 2262.190 ;
      LAYER li1 ;
        RECT 3382.055 2262.155 3384.555 2262.215 ;
        RECT 3382.055 2261.985 3383.220 2262.155 ;
        RECT 3383.390 2261.985 3384.555 2262.155 ;
        RECT 3382.055 2261.925 3384.555 2261.985 ;
        RECT 3385.215 2262.155 3386.110 2262.215 ;
        RECT 3385.215 2261.985 3385.940 2262.155 ;
        RECT 3385.215 2261.925 3386.110 2261.985 ;
        RECT 3382.030 2261.415 3383.050 2261.745 ;
        RECT 3383.220 2261.695 3383.390 2261.925 ;
        RECT 3385.940 2261.695 3386.110 2261.925 ;
        RECT 3382.030 2260.905 3382.200 2261.415 ;
        RECT 3383.220 2261.365 3383.390 2261.525 ;
        RECT 3385.940 2261.365 3386.110 2261.525 ;
        RECT 3383.220 2261.245 3384.540 2261.365 ;
        RECT 3382.420 2261.235 3384.540 2261.245 ;
        RECT 3382.420 2261.075 3383.220 2261.235 ;
        RECT 3383.390 2261.065 3384.540 2261.235 ;
        RECT 3383.220 2261.035 3384.540 2261.065 ;
        RECT 3385.140 2261.235 3386.110 2261.365 ;
        RECT 3385.140 2261.065 3385.940 2261.235 ;
        RECT 3385.140 2261.035 3386.110 2261.065 ;
        RECT 3382.030 2260.575 3383.050 2260.905 ;
        RECT 3383.220 2260.775 3383.390 2261.035 ;
      LAYER li1 ;
        RECT 3383.560 2260.695 3385.770 2260.865 ;
      LAYER li1 ;
        RECT 3385.940 2260.775 3386.110 2261.035 ;
      LAYER li1 ;
        RECT 3384.410 2260.610 3385.290 2260.695 ;
      LAYER li1 ;
        RECT 3382.030 2260.420 3382.200 2260.575 ;
        RECT 3381.320 2260.245 3382.200 2260.420 ;
        RECT 3383.220 2260.525 3383.390 2260.605 ;
        RECT 3383.220 2260.405 3384.190 2260.525 ;
        RECT 3382.420 2260.315 3384.190 2260.405 ;
        RECT 3380.500 2259.855 3380.670 2260.145 ;
      LAYER li1 ;
        RECT 3379.955 2256.410 3380.500 2259.830 ;
      LAYER li1 ;
        RECT 3380.500 2259.645 3380.670 2259.685 ;
        RECT 3380.500 2259.395 3381.150 2259.645 ;
        RECT 3380.670 2259.315 3381.150 2259.395 ;
        RECT 3380.500 2258.935 3380.670 2259.225 ;
        RECT 3380.670 2258.765 3381.150 2258.805 ;
        RECT 3380.500 2258.475 3381.150 2258.765 ;
        RECT 3380.500 2258.015 3380.670 2258.305 ;
        RECT 3380.670 2257.845 3381.150 2257.965 ;
        RECT 3380.500 2257.635 3381.150 2257.845 ;
        RECT 3381.660 2257.795 3381.830 2260.245 ;
        RECT 3382.420 2260.235 3383.220 2260.315 ;
        RECT 3383.390 2260.195 3384.190 2260.315 ;
        RECT 3383.220 2259.855 3383.390 2260.145 ;
      LAYER li1 ;
        RECT 3384.410 2260.025 3384.580 2260.610 ;
        RECT 3383.560 2259.855 3384.580 2260.025 ;
      LAYER li1 ;
        RECT 3383.220 2259.645 3384.190 2259.685 ;
        RECT 3382.420 2259.395 3384.190 2259.645 ;
        RECT 3382.420 2259.315 3383.220 2259.395 ;
        RECT 3383.390 2259.355 3384.190 2259.395 ;
        RECT 3383.220 2258.935 3383.390 2259.225 ;
      LAYER li1 ;
        RECT 3384.410 2259.185 3384.580 2259.855 ;
        RECT 3383.560 2259.015 3384.580 2259.185 ;
      LAYER li1 ;
        RECT 3382.420 2258.765 3383.220 2258.805 ;
        RECT 3383.390 2258.765 3384.190 2258.845 ;
        RECT 3382.420 2258.515 3384.190 2258.765 ;
        RECT 3382.420 2258.475 3383.390 2258.515 ;
      LAYER li1 ;
        RECT 3384.410 2258.345 3384.580 2259.015 ;
      LAYER li1 ;
        RECT 3383.220 2258.015 3383.390 2258.305 ;
      LAYER li1 ;
        RECT 3383.560 2258.175 3384.580 2258.345 ;
      LAYER li1 ;
        RECT 3382.420 2257.845 3383.220 2257.965 ;
        RECT 3383.390 2257.845 3384.190 2257.925 ;
        RECT 3384.780 2257.915 3384.950 2260.365 ;
      LAYER li1 ;
        RECT 3385.120 2260.025 3385.290 2260.610 ;
      LAYER li1 ;
        RECT 3385.940 2260.525 3386.110 2260.605 ;
        RECT 3385.460 2260.315 3386.110 2260.525 ;
        RECT 3385.460 2260.195 3385.940 2260.315 ;
      LAYER li1 ;
        RECT 3385.120 2259.855 3385.770 2260.025 ;
      LAYER li1 ;
        RECT 3385.940 2259.855 3386.110 2260.145 ;
      LAYER li1 ;
        RECT 3385.120 2259.185 3385.290 2259.855 ;
      LAYER li1 ;
        RECT 3385.460 2259.395 3386.110 2259.685 ;
        RECT 3385.460 2259.355 3385.940 2259.395 ;
      LAYER li1 ;
        RECT 3385.120 2259.015 3385.770 2259.185 ;
        RECT 3385.120 2258.345 3385.290 2259.015 ;
      LAYER li1 ;
        RECT 3385.940 2258.935 3386.110 2259.225 ;
        RECT 3385.460 2258.765 3385.940 2258.845 ;
        RECT 3385.460 2258.515 3386.110 2258.765 ;
        RECT 3385.940 2258.475 3386.110 2258.515 ;
      LAYER li1 ;
        RECT 3385.120 2258.175 3385.770 2258.345 ;
      LAYER li1 ;
        RECT 3385.940 2258.015 3386.110 2258.305 ;
        RECT 3382.420 2257.755 3384.190 2257.845 ;
        RECT 3382.420 2257.635 3383.390 2257.755 ;
        RECT 3380.500 2257.555 3380.670 2257.635 ;
        RECT 3383.220 2257.555 3383.390 2257.635 ;
        RECT 3384.410 2257.740 3385.290 2257.915 ;
        RECT 3384.410 2257.585 3384.580 2257.740 ;
        RECT 3380.500 2257.125 3380.670 2257.385 ;
        RECT 3383.220 2257.125 3383.390 2257.385 ;
        RECT 3383.560 2257.255 3384.580 2257.585 ;
        RECT 3380.500 2257.095 3381.470 2257.125 ;
        RECT 3380.670 2256.925 3381.470 2257.095 ;
        RECT 3380.500 2256.795 3381.470 2256.925 ;
        RECT 3382.070 2257.095 3383.390 2257.125 ;
        RECT 3382.070 2256.925 3383.220 2257.095 ;
        RECT 3383.390 2256.925 3384.190 2257.085 ;
        RECT 3382.070 2256.915 3384.190 2256.925 ;
        RECT 3382.070 2256.795 3383.390 2256.915 ;
        RECT 3380.500 2256.635 3380.670 2256.795 ;
        RECT 3383.220 2256.635 3383.390 2256.795 ;
        RECT 3384.410 2256.745 3384.580 2257.255 ;
        RECT 3377.780 2256.235 3377.950 2256.320 ;
        RECT 3380.500 2256.235 3380.670 2256.465 ;
        RECT 3383.220 2256.235 3383.390 2256.465 ;
        RECT 3383.560 2256.415 3384.580 2256.745 ;
        RECT 3385.120 2257.505 3385.290 2257.740 ;
        RECT 3385.460 2257.845 3385.940 2258.005 ;
        RECT 3385.460 2257.675 3386.110 2257.845 ;
        RECT 3385.940 2257.555 3386.110 2257.675 ;
        RECT 3385.120 2257.335 3385.765 2257.505 ;
        RECT 3385.120 2256.665 3385.290 2257.335 ;
        RECT 3385.940 2257.165 3386.110 2257.385 ;
        RECT 3385.460 2257.095 3386.110 2257.165 ;
        RECT 3385.460 2256.925 3385.940 2257.095 ;
        RECT 3385.460 2256.835 3386.110 2256.925 ;
        RECT 3385.120 2256.495 3385.770 2256.665 ;
        RECT 3385.940 2256.635 3386.110 2256.835 ;
        RECT 3385.940 2256.235 3386.110 2256.465 ;
        RECT 3377.780 2256.175 3379.115 2256.235 ;
        RECT 3377.950 2256.005 3379.115 2256.175 ;
        RECT 3377.780 2255.945 3379.115 2256.005 ;
        RECT 3379.775 2256.175 3381.395 2256.235 ;
        RECT 3379.775 2256.005 3380.500 2256.175 ;
        RECT 3380.670 2256.005 3381.395 2256.175 ;
        RECT 3379.775 2255.945 3381.395 2256.005 ;
        RECT 3377.780 2255.860 3377.950 2255.945 ;
      LAYER li1 ;
        RECT 3379.955 2254.190 3380.500 2255.775 ;
      LAYER li1 ;
        RECT 3380.500 2255.715 3380.670 2255.945 ;
        RECT 3380.500 2255.345 3380.670 2255.545 ;
        RECT 3380.840 2255.515 3381.490 2255.685 ;
        RECT 3380.500 2255.255 3381.150 2255.345 ;
        RECT 3380.670 2255.085 3381.150 2255.255 ;
        RECT 3380.500 2255.015 3381.150 2255.085 ;
        RECT 3380.500 2254.795 3380.670 2255.015 ;
        RECT 3381.320 2254.845 3381.490 2255.515 ;
        RECT 3380.845 2254.675 3381.490 2254.845 ;
        RECT 3380.500 2254.505 3380.670 2254.625 ;
        RECT 3380.500 2254.335 3381.150 2254.505 ;
      LAYER li1 ;
        RECT 3379.125 2253.850 3380.500 2254.190 ;
      LAYER li1 ;
        RECT 3380.670 2254.175 3381.150 2254.335 ;
        RECT 3381.320 2254.440 3381.490 2254.675 ;
      LAYER li1 ;
        RECT 3381.660 2254.620 3381.860 2256.210 ;
      LAYER li1 ;
        RECT 3382.055 2256.175 3384.555 2256.235 ;
        RECT 3382.055 2256.005 3383.220 2256.175 ;
        RECT 3383.390 2256.005 3384.555 2256.175 ;
        RECT 3382.055 2255.945 3384.555 2256.005 ;
        RECT 3385.215 2256.175 3386.110 2256.235 ;
        RECT 3385.215 2256.005 3385.940 2256.175 ;
        RECT 3385.215 2255.945 3386.110 2256.005 ;
        RECT 3382.030 2255.435 3383.050 2255.765 ;
        RECT 3383.220 2255.715 3383.390 2255.945 ;
        RECT 3385.940 2255.715 3386.110 2255.945 ;
        RECT 3382.030 2254.925 3382.200 2255.435 ;
        RECT 3383.220 2255.385 3383.390 2255.545 ;
        RECT 3385.940 2255.385 3386.110 2255.545 ;
        RECT 3383.220 2255.265 3384.540 2255.385 ;
        RECT 3382.420 2255.255 3384.540 2255.265 ;
        RECT 3382.420 2255.095 3383.220 2255.255 ;
        RECT 3383.390 2255.085 3384.540 2255.255 ;
        RECT 3383.220 2255.055 3384.540 2255.085 ;
        RECT 3385.140 2255.255 3386.110 2255.385 ;
        RECT 3385.140 2255.085 3385.940 2255.255 ;
        RECT 3385.140 2255.055 3386.110 2255.085 ;
        RECT 3382.030 2254.595 3383.050 2254.925 ;
        RECT 3383.220 2254.795 3383.390 2255.055 ;
      LAYER li1 ;
        RECT 3383.560 2254.715 3385.770 2254.885 ;
      LAYER li1 ;
        RECT 3385.940 2254.795 3386.110 2255.055 ;
      LAYER li1 ;
        RECT 3384.410 2254.630 3385.290 2254.715 ;
      LAYER li1 ;
        RECT 3382.030 2254.440 3382.200 2254.595 ;
        RECT 3381.320 2254.265 3382.200 2254.440 ;
        RECT 3383.220 2254.545 3383.390 2254.625 ;
        RECT 3383.220 2254.425 3384.190 2254.545 ;
        RECT 3382.420 2254.335 3384.190 2254.425 ;
        RECT 3380.500 2253.875 3380.670 2254.165 ;
      LAYER li1 ;
        RECT 3379.955 2250.430 3380.500 2253.850 ;
      LAYER li1 ;
        RECT 3380.500 2253.665 3380.670 2253.705 ;
        RECT 3380.500 2253.415 3381.150 2253.665 ;
        RECT 3380.670 2253.335 3381.150 2253.415 ;
        RECT 3380.500 2252.955 3380.670 2253.245 ;
        RECT 3380.670 2252.785 3381.150 2252.825 ;
        RECT 3380.500 2252.495 3381.150 2252.785 ;
        RECT 3380.500 2252.035 3380.670 2252.325 ;
        RECT 3380.670 2251.865 3381.150 2251.985 ;
        RECT 3380.500 2251.655 3381.150 2251.865 ;
        RECT 3381.660 2251.815 3381.830 2254.265 ;
        RECT 3382.420 2254.255 3383.220 2254.335 ;
        RECT 3383.390 2254.215 3384.190 2254.335 ;
        RECT 3383.220 2253.875 3383.390 2254.165 ;
      LAYER li1 ;
        RECT 3384.410 2254.045 3384.580 2254.630 ;
        RECT 3383.560 2253.875 3384.580 2254.045 ;
      LAYER li1 ;
        RECT 3383.220 2253.665 3384.190 2253.705 ;
        RECT 3382.420 2253.415 3384.190 2253.665 ;
        RECT 3382.420 2253.335 3383.220 2253.415 ;
        RECT 3383.390 2253.375 3384.190 2253.415 ;
        RECT 3383.220 2252.955 3383.390 2253.245 ;
      LAYER li1 ;
        RECT 3384.410 2253.205 3384.580 2253.875 ;
        RECT 3383.560 2253.035 3384.580 2253.205 ;
      LAYER li1 ;
        RECT 3382.420 2252.785 3383.220 2252.825 ;
        RECT 3383.390 2252.785 3384.190 2252.865 ;
        RECT 3382.420 2252.535 3384.190 2252.785 ;
        RECT 3382.420 2252.495 3383.390 2252.535 ;
      LAYER li1 ;
        RECT 3384.410 2252.365 3384.580 2253.035 ;
      LAYER li1 ;
        RECT 3383.220 2252.035 3383.390 2252.325 ;
      LAYER li1 ;
        RECT 3383.560 2252.195 3384.580 2252.365 ;
      LAYER li1 ;
        RECT 3382.420 2251.865 3383.220 2251.985 ;
        RECT 3383.390 2251.865 3384.190 2251.945 ;
        RECT 3384.780 2251.935 3384.950 2254.385 ;
      LAYER li1 ;
        RECT 3385.120 2254.045 3385.290 2254.630 ;
      LAYER li1 ;
        RECT 3385.940 2254.545 3386.110 2254.625 ;
        RECT 3385.460 2254.335 3386.110 2254.545 ;
        RECT 3385.460 2254.215 3385.940 2254.335 ;
      LAYER li1 ;
        RECT 3385.120 2253.875 3385.770 2254.045 ;
      LAYER li1 ;
        RECT 3385.940 2253.875 3386.110 2254.165 ;
      LAYER li1 ;
        RECT 3385.120 2253.205 3385.290 2253.875 ;
      LAYER li1 ;
        RECT 3385.460 2253.415 3386.110 2253.705 ;
        RECT 3385.460 2253.375 3385.940 2253.415 ;
      LAYER li1 ;
        RECT 3385.120 2253.035 3385.770 2253.205 ;
        RECT 3385.120 2252.365 3385.290 2253.035 ;
      LAYER li1 ;
        RECT 3385.940 2252.955 3386.110 2253.245 ;
        RECT 3385.460 2252.785 3385.940 2252.865 ;
        RECT 3385.460 2252.535 3386.110 2252.785 ;
        RECT 3385.940 2252.495 3386.110 2252.535 ;
      LAYER li1 ;
        RECT 3385.120 2252.195 3385.770 2252.365 ;
      LAYER li1 ;
        RECT 3385.940 2252.035 3386.110 2252.325 ;
        RECT 3382.420 2251.775 3384.190 2251.865 ;
        RECT 3382.420 2251.655 3383.390 2251.775 ;
        RECT 3380.500 2251.575 3380.670 2251.655 ;
        RECT 3383.220 2251.575 3383.390 2251.655 ;
        RECT 3384.410 2251.760 3385.290 2251.935 ;
        RECT 3384.410 2251.605 3384.580 2251.760 ;
        RECT 3380.500 2251.145 3380.670 2251.405 ;
        RECT 3383.220 2251.145 3383.390 2251.405 ;
        RECT 3383.560 2251.275 3384.580 2251.605 ;
        RECT 3380.500 2251.115 3381.470 2251.145 ;
        RECT 3380.670 2250.945 3381.470 2251.115 ;
        RECT 3380.500 2250.815 3381.470 2250.945 ;
        RECT 3382.070 2251.115 3383.390 2251.145 ;
        RECT 3382.070 2250.945 3383.220 2251.115 ;
        RECT 3383.390 2250.945 3384.190 2251.105 ;
        RECT 3382.070 2250.935 3384.190 2250.945 ;
        RECT 3382.070 2250.815 3383.390 2250.935 ;
        RECT 3380.500 2250.655 3380.670 2250.815 ;
        RECT 3383.220 2250.655 3383.390 2250.815 ;
        RECT 3384.410 2250.765 3384.580 2251.275 ;
        RECT 3377.780 2250.255 3377.950 2250.340 ;
        RECT 3380.500 2250.255 3380.670 2250.485 ;
        RECT 3383.220 2250.255 3383.390 2250.485 ;
        RECT 3383.560 2250.435 3384.580 2250.765 ;
        RECT 3385.120 2251.525 3385.290 2251.760 ;
        RECT 3385.460 2251.865 3385.940 2252.025 ;
        RECT 3385.460 2251.695 3386.110 2251.865 ;
        RECT 3385.940 2251.575 3386.110 2251.695 ;
        RECT 3385.120 2251.355 3385.765 2251.525 ;
        RECT 3385.120 2250.685 3385.290 2251.355 ;
        RECT 3385.940 2251.185 3386.110 2251.405 ;
        RECT 3385.460 2251.115 3386.110 2251.185 ;
        RECT 3385.460 2250.945 3385.940 2251.115 ;
        RECT 3385.460 2250.855 3386.110 2250.945 ;
        RECT 3385.120 2250.515 3385.770 2250.685 ;
        RECT 3385.940 2250.655 3386.110 2250.855 ;
        RECT 3385.940 2250.255 3386.110 2250.485 ;
        RECT 3377.780 2250.195 3379.115 2250.255 ;
        RECT 3377.950 2250.025 3379.115 2250.195 ;
        RECT 3377.780 2249.965 3379.115 2250.025 ;
        RECT 3379.775 2250.195 3381.395 2250.255 ;
        RECT 3379.775 2250.025 3380.500 2250.195 ;
        RECT 3380.670 2250.025 3381.395 2250.195 ;
        RECT 3379.775 2249.965 3381.395 2250.025 ;
        RECT 3377.780 2249.880 3377.950 2249.965 ;
      LAYER li1 ;
        RECT 3379.955 2248.210 3380.500 2249.795 ;
      LAYER li1 ;
        RECT 3380.500 2249.735 3380.670 2249.965 ;
        RECT 3380.500 2249.365 3380.670 2249.565 ;
        RECT 3380.840 2249.535 3381.490 2249.705 ;
        RECT 3380.500 2249.275 3381.150 2249.365 ;
        RECT 3380.670 2249.105 3381.150 2249.275 ;
        RECT 3380.500 2249.035 3381.150 2249.105 ;
        RECT 3380.500 2248.815 3380.670 2249.035 ;
        RECT 3381.320 2248.865 3381.490 2249.535 ;
        RECT 3380.845 2248.695 3381.490 2248.865 ;
        RECT 3380.500 2248.525 3380.670 2248.645 ;
        RECT 3380.500 2248.355 3381.150 2248.525 ;
      LAYER li1 ;
        RECT 3379.125 2247.870 3380.500 2248.210 ;
      LAYER li1 ;
        RECT 3380.670 2248.195 3381.150 2248.355 ;
        RECT 3381.320 2248.460 3381.490 2248.695 ;
      LAYER li1 ;
        RECT 3381.660 2248.640 3381.860 2250.230 ;
      LAYER li1 ;
        RECT 3382.055 2250.195 3384.555 2250.255 ;
        RECT 3382.055 2250.025 3383.220 2250.195 ;
        RECT 3383.390 2250.025 3384.555 2250.195 ;
        RECT 3382.055 2249.965 3384.555 2250.025 ;
        RECT 3385.215 2250.195 3386.110 2250.255 ;
        RECT 3385.215 2250.025 3385.940 2250.195 ;
        RECT 3385.215 2249.965 3386.110 2250.025 ;
        RECT 3382.030 2249.455 3383.050 2249.785 ;
        RECT 3383.220 2249.735 3383.390 2249.965 ;
        RECT 3385.940 2249.735 3386.110 2249.965 ;
        RECT 3382.030 2248.945 3382.200 2249.455 ;
        RECT 3383.220 2249.405 3383.390 2249.565 ;
        RECT 3385.940 2249.405 3386.110 2249.565 ;
        RECT 3383.220 2249.285 3384.540 2249.405 ;
        RECT 3382.420 2249.275 3384.540 2249.285 ;
        RECT 3382.420 2249.115 3383.220 2249.275 ;
        RECT 3383.390 2249.105 3384.540 2249.275 ;
        RECT 3383.220 2249.075 3384.540 2249.105 ;
        RECT 3385.140 2249.275 3386.110 2249.405 ;
        RECT 3385.140 2249.105 3385.940 2249.275 ;
        RECT 3385.140 2249.075 3386.110 2249.105 ;
        RECT 3382.030 2248.615 3383.050 2248.945 ;
        RECT 3383.220 2248.815 3383.390 2249.075 ;
      LAYER li1 ;
        RECT 3383.560 2248.735 3385.770 2248.905 ;
      LAYER li1 ;
        RECT 3385.940 2248.815 3386.110 2249.075 ;
      LAYER li1 ;
        RECT 3384.410 2248.650 3385.290 2248.735 ;
      LAYER li1 ;
        RECT 3382.030 2248.460 3382.200 2248.615 ;
        RECT 3381.320 2248.285 3382.200 2248.460 ;
        RECT 3383.220 2248.565 3383.390 2248.645 ;
        RECT 3383.220 2248.445 3384.190 2248.565 ;
        RECT 3382.420 2248.355 3384.190 2248.445 ;
        RECT 3380.500 2247.895 3380.670 2248.185 ;
      LAYER li1 ;
        RECT 3379.955 2244.450 3380.500 2247.870 ;
      LAYER li1 ;
        RECT 3380.500 2247.685 3380.670 2247.725 ;
        RECT 3380.500 2247.435 3381.150 2247.685 ;
        RECT 3380.670 2247.355 3381.150 2247.435 ;
        RECT 3380.500 2246.975 3380.670 2247.265 ;
        RECT 3380.670 2246.805 3381.150 2246.845 ;
        RECT 3380.500 2246.515 3381.150 2246.805 ;
        RECT 3380.500 2246.055 3380.670 2246.345 ;
        RECT 3380.670 2245.885 3381.150 2246.005 ;
        RECT 3380.500 2245.675 3381.150 2245.885 ;
        RECT 3381.660 2245.835 3381.830 2248.285 ;
        RECT 3382.420 2248.275 3383.220 2248.355 ;
        RECT 3383.390 2248.235 3384.190 2248.355 ;
        RECT 3383.220 2247.895 3383.390 2248.185 ;
      LAYER li1 ;
        RECT 3384.410 2248.065 3384.580 2248.650 ;
        RECT 3383.560 2247.895 3384.580 2248.065 ;
      LAYER li1 ;
        RECT 3383.220 2247.685 3384.190 2247.725 ;
        RECT 3382.420 2247.435 3384.190 2247.685 ;
        RECT 3382.420 2247.355 3383.220 2247.435 ;
        RECT 3383.390 2247.395 3384.190 2247.435 ;
        RECT 3383.220 2246.975 3383.390 2247.265 ;
      LAYER li1 ;
        RECT 3384.410 2247.225 3384.580 2247.895 ;
        RECT 3383.560 2247.055 3384.580 2247.225 ;
      LAYER li1 ;
        RECT 3382.420 2246.805 3383.220 2246.845 ;
        RECT 3383.390 2246.805 3384.190 2246.885 ;
        RECT 3382.420 2246.555 3384.190 2246.805 ;
        RECT 3382.420 2246.515 3383.390 2246.555 ;
      LAYER li1 ;
        RECT 3384.410 2246.385 3384.580 2247.055 ;
      LAYER li1 ;
        RECT 3383.220 2246.055 3383.390 2246.345 ;
      LAYER li1 ;
        RECT 3383.560 2246.215 3384.580 2246.385 ;
      LAYER li1 ;
        RECT 3382.420 2245.885 3383.220 2246.005 ;
        RECT 3383.390 2245.885 3384.190 2245.965 ;
        RECT 3384.780 2245.955 3384.950 2248.405 ;
      LAYER li1 ;
        RECT 3385.120 2248.065 3385.290 2248.650 ;
      LAYER li1 ;
        RECT 3385.940 2248.565 3386.110 2248.645 ;
        RECT 3385.460 2248.355 3386.110 2248.565 ;
        RECT 3385.460 2248.235 3385.940 2248.355 ;
      LAYER li1 ;
        RECT 3385.120 2247.895 3385.770 2248.065 ;
      LAYER li1 ;
        RECT 3385.940 2247.895 3386.110 2248.185 ;
      LAYER li1 ;
        RECT 3385.120 2247.225 3385.290 2247.895 ;
      LAYER li1 ;
        RECT 3385.460 2247.435 3386.110 2247.725 ;
        RECT 3385.460 2247.395 3385.940 2247.435 ;
      LAYER li1 ;
        RECT 3385.120 2247.055 3385.770 2247.225 ;
        RECT 3385.120 2246.385 3385.290 2247.055 ;
      LAYER li1 ;
        RECT 3385.940 2246.975 3386.110 2247.265 ;
        RECT 3385.460 2246.805 3385.940 2246.885 ;
        RECT 3385.460 2246.555 3386.110 2246.805 ;
        RECT 3385.940 2246.515 3386.110 2246.555 ;
      LAYER li1 ;
        RECT 3385.120 2246.215 3385.770 2246.385 ;
      LAYER li1 ;
        RECT 3385.940 2246.055 3386.110 2246.345 ;
        RECT 3382.420 2245.795 3384.190 2245.885 ;
        RECT 3382.420 2245.675 3383.390 2245.795 ;
        RECT 3380.500 2245.595 3380.670 2245.675 ;
        RECT 3383.220 2245.595 3383.390 2245.675 ;
        RECT 3384.410 2245.780 3385.290 2245.955 ;
        RECT 3384.410 2245.625 3384.580 2245.780 ;
        RECT 3380.500 2245.165 3380.670 2245.425 ;
        RECT 3383.220 2245.165 3383.390 2245.425 ;
        RECT 3383.560 2245.295 3384.580 2245.625 ;
        RECT 3380.500 2245.135 3381.470 2245.165 ;
        RECT 3380.670 2244.965 3381.470 2245.135 ;
        RECT 3380.500 2244.835 3381.470 2244.965 ;
        RECT 3382.070 2245.135 3383.390 2245.165 ;
        RECT 3382.070 2244.965 3383.220 2245.135 ;
        RECT 3383.390 2244.965 3384.190 2245.125 ;
        RECT 3382.070 2244.955 3384.190 2244.965 ;
        RECT 3382.070 2244.835 3383.390 2244.955 ;
        RECT 3380.500 2244.675 3380.670 2244.835 ;
        RECT 3383.220 2244.675 3383.390 2244.835 ;
        RECT 3384.410 2244.785 3384.580 2245.295 ;
        RECT 3377.780 2244.275 3377.950 2244.360 ;
        RECT 3380.500 2244.275 3380.670 2244.505 ;
        RECT 3383.220 2244.275 3383.390 2244.505 ;
        RECT 3383.560 2244.455 3384.580 2244.785 ;
        RECT 3385.120 2245.545 3385.290 2245.780 ;
        RECT 3385.460 2245.885 3385.940 2246.045 ;
        RECT 3385.460 2245.715 3386.110 2245.885 ;
        RECT 3385.940 2245.595 3386.110 2245.715 ;
        RECT 3385.120 2245.375 3385.765 2245.545 ;
        RECT 3385.120 2244.705 3385.290 2245.375 ;
        RECT 3385.940 2245.205 3386.110 2245.425 ;
        RECT 3385.460 2245.135 3386.110 2245.205 ;
        RECT 3385.460 2244.965 3385.940 2245.135 ;
        RECT 3385.460 2244.875 3386.110 2244.965 ;
        RECT 3385.120 2244.535 3385.770 2244.705 ;
        RECT 3385.940 2244.675 3386.110 2244.875 ;
        RECT 3385.940 2244.275 3386.110 2244.505 ;
        RECT 3377.780 2244.215 3379.115 2244.275 ;
        RECT 3377.950 2244.045 3379.115 2244.215 ;
        RECT 3377.780 2243.985 3379.115 2244.045 ;
        RECT 3379.775 2244.215 3381.395 2244.275 ;
        RECT 3379.775 2244.045 3380.500 2244.215 ;
        RECT 3380.670 2244.045 3381.395 2244.215 ;
        RECT 3379.775 2243.985 3381.395 2244.045 ;
        RECT 3377.780 2243.900 3377.950 2243.985 ;
      LAYER li1 ;
        RECT 3379.955 2242.230 3380.500 2243.815 ;
      LAYER li1 ;
        RECT 3380.500 2243.755 3380.670 2243.985 ;
        RECT 3380.500 2243.385 3380.670 2243.585 ;
        RECT 3380.840 2243.555 3381.490 2243.725 ;
        RECT 3380.500 2243.295 3381.150 2243.385 ;
        RECT 3380.670 2243.125 3381.150 2243.295 ;
        RECT 3380.500 2243.055 3381.150 2243.125 ;
        RECT 3380.500 2242.835 3380.670 2243.055 ;
        RECT 3381.320 2242.885 3381.490 2243.555 ;
        RECT 3380.845 2242.715 3381.490 2242.885 ;
        RECT 3380.500 2242.545 3380.670 2242.665 ;
        RECT 3380.500 2242.375 3381.150 2242.545 ;
      LAYER li1 ;
        RECT 3379.125 2241.890 3380.500 2242.230 ;
      LAYER li1 ;
        RECT 3380.670 2242.215 3381.150 2242.375 ;
        RECT 3381.320 2242.480 3381.490 2242.715 ;
      LAYER li1 ;
        RECT 3381.660 2242.660 3381.860 2244.250 ;
      LAYER li1 ;
        RECT 3382.055 2244.215 3384.555 2244.275 ;
        RECT 3382.055 2244.045 3383.220 2244.215 ;
        RECT 3383.390 2244.045 3384.555 2244.215 ;
        RECT 3382.055 2243.985 3384.555 2244.045 ;
        RECT 3385.215 2244.215 3386.110 2244.275 ;
        RECT 3385.215 2244.045 3385.940 2244.215 ;
        RECT 3385.215 2243.985 3386.110 2244.045 ;
        RECT 3382.030 2243.475 3383.050 2243.805 ;
        RECT 3383.220 2243.755 3383.390 2243.985 ;
        RECT 3385.940 2243.755 3386.110 2243.985 ;
        RECT 3382.030 2242.965 3382.200 2243.475 ;
        RECT 3383.220 2243.425 3383.390 2243.585 ;
        RECT 3385.940 2243.425 3386.110 2243.585 ;
        RECT 3383.220 2243.305 3384.540 2243.425 ;
        RECT 3382.420 2243.295 3384.540 2243.305 ;
        RECT 3382.420 2243.135 3383.220 2243.295 ;
        RECT 3383.390 2243.125 3384.540 2243.295 ;
        RECT 3383.220 2243.095 3384.540 2243.125 ;
        RECT 3385.140 2243.295 3386.110 2243.425 ;
        RECT 3385.140 2243.125 3385.940 2243.295 ;
        RECT 3385.140 2243.095 3386.110 2243.125 ;
        RECT 3382.030 2242.635 3383.050 2242.965 ;
        RECT 3383.220 2242.835 3383.390 2243.095 ;
      LAYER li1 ;
        RECT 3383.560 2242.755 3385.770 2242.925 ;
      LAYER li1 ;
        RECT 3385.940 2242.835 3386.110 2243.095 ;
      LAYER li1 ;
        RECT 3384.410 2242.670 3385.290 2242.755 ;
      LAYER li1 ;
        RECT 3382.030 2242.480 3382.200 2242.635 ;
        RECT 3381.320 2242.305 3382.200 2242.480 ;
        RECT 3383.220 2242.585 3383.390 2242.665 ;
        RECT 3383.220 2242.465 3384.190 2242.585 ;
        RECT 3382.420 2242.375 3384.190 2242.465 ;
        RECT 3380.500 2241.915 3380.670 2242.205 ;
      LAYER li1 ;
        RECT 3379.955 2238.470 3380.500 2241.890 ;
      LAYER li1 ;
        RECT 3380.500 2241.705 3380.670 2241.745 ;
        RECT 3380.500 2241.455 3381.150 2241.705 ;
        RECT 3380.670 2241.375 3381.150 2241.455 ;
        RECT 3380.500 2240.995 3380.670 2241.285 ;
        RECT 3380.670 2240.825 3381.150 2240.865 ;
        RECT 3380.500 2240.535 3381.150 2240.825 ;
        RECT 3380.500 2240.075 3380.670 2240.365 ;
        RECT 3380.670 2239.905 3381.150 2240.025 ;
        RECT 3380.500 2239.695 3381.150 2239.905 ;
        RECT 3381.660 2239.855 3381.830 2242.305 ;
        RECT 3382.420 2242.295 3383.220 2242.375 ;
        RECT 3383.390 2242.255 3384.190 2242.375 ;
        RECT 3383.220 2241.915 3383.390 2242.205 ;
      LAYER li1 ;
        RECT 3384.410 2242.085 3384.580 2242.670 ;
        RECT 3383.560 2241.915 3384.580 2242.085 ;
      LAYER li1 ;
        RECT 3383.220 2241.705 3384.190 2241.745 ;
        RECT 3382.420 2241.455 3384.190 2241.705 ;
        RECT 3382.420 2241.375 3383.220 2241.455 ;
        RECT 3383.390 2241.415 3384.190 2241.455 ;
        RECT 3383.220 2240.995 3383.390 2241.285 ;
      LAYER li1 ;
        RECT 3384.410 2241.245 3384.580 2241.915 ;
        RECT 3383.560 2241.075 3384.580 2241.245 ;
      LAYER li1 ;
        RECT 3382.420 2240.825 3383.220 2240.865 ;
        RECT 3383.390 2240.825 3384.190 2240.905 ;
        RECT 3382.420 2240.575 3384.190 2240.825 ;
        RECT 3382.420 2240.535 3383.390 2240.575 ;
      LAYER li1 ;
        RECT 3384.410 2240.405 3384.580 2241.075 ;
      LAYER li1 ;
        RECT 3383.220 2240.075 3383.390 2240.365 ;
      LAYER li1 ;
        RECT 3383.560 2240.235 3384.580 2240.405 ;
      LAYER li1 ;
        RECT 3382.420 2239.905 3383.220 2240.025 ;
        RECT 3383.390 2239.905 3384.190 2239.985 ;
        RECT 3384.780 2239.975 3384.950 2242.425 ;
      LAYER li1 ;
        RECT 3385.120 2242.085 3385.290 2242.670 ;
      LAYER li1 ;
        RECT 3385.940 2242.585 3386.110 2242.665 ;
        RECT 3385.460 2242.375 3386.110 2242.585 ;
        RECT 3385.460 2242.255 3385.940 2242.375 ;
      LAYER li1 ;
        RECT 3385.120 2241.915 3385.770 2242.085 ;
      LAYER li1 ;
        RECT 3385.940 2241.915 3386.110 2242.205 ;
      LAYER li1 ;
        RECT 3385.120 2241.245 3385.290 2241.915 ;
      LAYER li1 ;
        RECT 3385.460 2241.455 3386.110 2241.745 ;
        RECT 3385.460 2241.415 3385.940 2241.455 ;
      LAYER li1 ;
        RECT 3385.120 2241.075 3385.770 2241.245 ;
        RECT 3385.120 2240.405 3385.290 2241.075 ;
      LAYER li1 ;
        RECT 3385.940 2240.995 3386.110 2241.285 ;
        RECT 3385.460 2240.825 3385.940 2240.905 ;
        RECT 3385.460 2240.575 3386.110 2240.825 ;
        RECT 3385.940 2240.535 3386.110 2240.575 ;
      LAYER li1 ;
        RECT 3385.120 2240.235 3385.770 2240.405 ;
      LAYER li1 ;
        RECT 3385.940 2240.075 3386.110 2240.365 ;
        RECT 3382.420 2239.815 3384.190 2239.905 ;
        RECT 3382.420 2239.695 3383.390 2239.815 ;
        RECT 3380.500 2239.615 3380.670 2239.695 ;
        RECT 3383.220 2239.615 3383.390 2239.695 ;
        RECT 3384.410 2239.800 3385.290 2239.975 ;
        RECT 3384.410 2239.645 3384.580 2239.800 ;
        RECT 3380.500 2239.185 3380.670 2239.445 ;
        RECT 3383.220 2239.185 3383.390 2239.445 ;
        RECT 3383.560 2239.315 3384.580 2239.645 ;
        RECT 3380.500 2239.155 3381.470 2239.185 ;
        RECT 3380.670 2238.985 3381.470 2239.155 ;
        RECT 3380.500 2238.855 3381.470 2238.985 ;
        RECT 3382.070 2239.155 3383.390 2239.185 ;
        RECT 3382.070 2238.985 3383.220 2239.155 ;
        RECT 3383.390 2238.985 3384.190 2239.145 ;
        RECT 3382.070 2238.975 3384.190 2238.985 ;
        RECT 3382.070 2238.855 3383.390 2238.975 ;
        RECT 3380.500 2238.695 3380.670 2238.855 ;
        RECT 3383.220 2238.695 3383.390 2238.855 ;
        RECT 3384.410 2238.805 3384.580 2239.315 ;
        RECT 3377.780 2238.295 3377.950 2238.380 ;
        RECT 3380.500 2238.295 3380.670 2238.525 ;
        RECT 3383.220 2238.295 3383.390 2238.525 ;
        RECT 3383.560 2238.475 3384.580 2238.805 ;
        RECT 3385.120 2239.565 3385.290 2239.800 ;
        RECT 3385.460 2239.905 3385.940 2240.065 ;
        RECT 3385.460 2239.735 3386.110 2239.905 ;
        RECT 3385.940 2239.615 3386.110 2239.735 ;
        RECT 3385.120 2239.395 3385.765 2239.565 ;
        RECT 3385.120 2238.725 3385.290 2239.395 ;
        RECT 3385.940 2239.225 3386.110 2239.445 ;
        RECT 3385.460 2239.155 3386.110 2239.225 ;
        RECT 3385.460 2238.985 3385.940 2239.155 ;
        RECT 3385.460 2238.895 3386.110 2238.985 ;
        RECT 3385.120 2238.555 3385.770 2238.725 ;
        RECT 3385.940 2238.695 3386.110 2238.895 ;
        RECT 3385.940 2238.295 3386.110 2238.525 ;
        RECT 3377.780 2238.235 3379.115 2238.295 ;
        RECT 3377.950 2238.065 3379.115 2238.235 ;
        RECT 3377.780 2238.005 3379.115 2238.065 ;
        RECT 3379.775 2238.235 3381.395 2238.295 ;
        RECT 3379.775 2238.065 3380.500 2238.235 ;
        RECT 3380.670 2238.065 3381.395 2238.235 ;
        RECT 3379.775 2238.005 3381.395 2238.065 ;
        RECT 3377.780 2237.920 3377.950 2238.005 ;
      LAYER li1 ;
        RECT 3379.955 2236.250 3380.500 2237.835 ;
      LAYER li1 ;
        RECT 3380.500 2237.775 3380.670 2238.005 ;
        RECT 3380.500 2237.405 3380.670 2237.605 ;
        RECT 3380.840 2237.575 3381.490 2237.745 ;
        RECT 3380.500 2237.315 3381.150 2237.405 ;
        RECT 3380.670 2237.145 3381.150 2237.315 ;
        RECT 3380.500 2237.075 3381.150 2237.145 ;
        RECT 3380.500 2236.855 3380.670 2237.075 ;
        RECT 3381.320 2236.905 3381.490 2237.575 ;
        RECT 3380.845 2236.735 3381.490 2236.905 ;
        RECT 3380.500 2236.565 3380.670 2236.685 ;
        RECT 3380.500 2236.395 3381.150 2236.565 ;
      LAYER li1 ;
        RECT 3379.125 2235.910 3380.500 2236.250 ;
      LAYER li1 ;
        RECT 3380.670 2236.235 3381.150 2236.395 ;
        RECT 3381.320 2236.500 3381.490 2236.735 ;
      LAYER li1 ;
        RECT 3381.660 2236.680 3381.860 2238.270 ;
      LAYER li1 ;
        RECT 3382.055 2238.235 3384.555 2238.295 ;
        RECT 3382.055 2238.065 3383.220 2238.235 ;
        RECT 3383.390 2238.065 3384.555 2238.235 ;
        RECT 3382.055 2238.005 3384.555 2238.065 ;
        RECT 3385.215 2238.235 3386.110 2238.295 ;
        RECT 3385.215 2238.065 3385.940 2238.235 ;
        RECT 3385.215 2238.005 3386.110 2238.065 ;
        RECT 3382.030 2237.495 3383.050 2237.825 ;
        RECT 3383.220 2237.775 3383.390 2238.005 ;
        RECT 3385.940 2237.775 3386.110 2238.005 ;
        RECT 3382.030 2236.985 3382.200 2237.495 ;
        RECT 3383.220 2237.445 3383.390 2237.605 ;
        RECT 3385.940 2237.445 3386.110 2237.605 ;
        RECT 3383.220 2237.325 3384.540 2237.445 ;
        RECT 3382.420 2237.315 3384.540 2237.325 ;
        RECT 3382.420 2237.155 3383.220 2237.315 ;
        RECT 3383.390 2237.145 3384.540 2237.315 ;
        RECT 3383.220 2237.115 3384.540 2237.145 ;
        RECT 3385.140 2237.315 3386.110 2237.445 ;
        RECT 3385.140 2237.145 3385.940 2237.315 ;
        RECT 3385.140 2237.115 3386.110 2237.145 ;
        RECT 3382.030 2236.655 3383.050 2236.985 ;
        RECT 3383.220 2236.855 3383.390 2237.115 ;
      LAYER li1 ;
        RECT 3383.560 2236.775 3385.770 2236.945 ;
      LAYER li1 ;
        RECT 3385.940 2236.855 3386.110 2237.115 ;
      LAYER li1 ;
        RECT 3384.410 2236.690 3385.290 2236.775 ;
      LAYER li1 ;
        RECT 3382.030 2236.500 3382.200 2236.655 ;
        RECT 3381.320 2236.325 3382.200 2236.500 ;
        RECT 3383.220 2236.605 3383.390 2236.685 ;
        RECT 3383.220 2236.485 3384.190 2236.605 ;
        RECT 3382.420 2236.395 3384.190 2236.485 ;
        RECT 3380.500 2235.935 3380.670 2236.225 ;
      LAYER li1 ;
        RECT 3379.955 2232.490 3380.500 2235.910 ;
      LAYER li1 ;
        RECT 3380.500 2235.725 3380.670 2235.765 ;
        RECT 3380.500 2235.475 3381.150 2235.725 ;
        RECT 3380.670 2235.395 3381.150 2235.475 ;
        RECT 3380.500 2235.015 3380.670 2235.305 ;
        RECT 3380.670 2234.845 3381.150 2234.885 ;
        RECT 3380.500 2234.555 3381.150 2234.845 ;
        RECT 3380.500 2234.095 3380.670 2234.385 ;
        RECT 3380.670 2233.925 3381.150 2234.045 ;
        RECT 3380.500 2233.715 3381.150 2233.925 ;
        RECT 3381.660 2233.875 3381.830 2236.325 ;
        RECT 3382.420 2236.315 3383.220 2236.395 ;
        RECT 3383.390 2236.275 3384.190 2236.395 ;
        RECT 3383.220 2235.935 3383.390 2236.225 ;
      LAYER li1 ;
        RECT 3384.410 2236.105 3384.580 2236.690 ;
        RECT 3383.560 2235.935 3384.580 2236.105 ;
      LAYER li1 ;
        RECT 3383.220 2235.725 3384.190 2235.765 ;
        RECT 3382.420 2235.475 3384.190 2235.725 ;
        RECT 3382.420 2235.395 3383.220 2235.475 ;
        RECT 3383.390 2235.435 3384.190 2235.475 ;
        RECT 3383.220 2235.015 3383.390 2235.305 ;
      LAYER li1 ;
        RECT 3384.410 2235.265 3384.580 2235.935 ;
        RECT 3383.560 2235.095 3384.580 2235.265 ;
      LAYER li1 ;
        RECT 3382.420 2234.845 3383.220 2234.885 ;
        RECT 3383.390 2234.845 3384.190 2234.925 ;
        RECT 3382.420 2234.595 3384.190 2234.845 ;
        RECT 3382.420 2234.555 3383.390 2234.595 ;
      LAYER li1 ;
        RECT 3384.410 2234.425 3384.580 2235.095 ;
      LAYER li1 ;
        RECT 3383.220 2234.095 3383.390 2234.385 ;
      LAYER li1 ;
        RECT 3383.560 2234.255 3384.580 2234.425 ;
      LAYER li1 ;
        RECT 3382.420 2233.925 3383.220 2234.045 ;
        RECT 3383.390 2233.925 3384.190 2234.005 ;
        RECT 3384.780 2233.995 3384.950 2236.445 ;
      LAYER li1 ;
        RECT 3385.120 2236.105 3385.290 2236.690 ;
      LAYER li1 ;
        RECT 3385.940 2236.605 3386.110 2236.685 ;
        RECT 3385.460 2236.395 3386.110 2236.605 ;
        RECT 3385.460 2236.275 3385.940 2236.395 ;
      LAYER li1 ;
        RECT 3385.120 2235.935 3385.770 2236.105 ;
      LAYER li1 ;
        RECT 3385.940 2235.935 3386.110 2236.225 ;
      LAYER li1 ;
        RECT 3385.120 2235.265 3385.290 2235.935 ;
      LAYER li1 ;
        RECT 3385.460 2235.475 3386.110 2235.765 ;
        RECT 3385.460 2235.435 3385.940 2235.475 ;
      LAYER li1 ;
        RECT 3385.120 2235.095 3385.770 2235.265 ;
        RECT 3385.120 2234.425 3385.290 2235.095 ;
      LAYER li1 ;
        RECT 3385.940 2235.015 3386.110 2235.305 ;
        RECT 3385.460 2234.845 3385.940 2234.925 ;
        RECT 3385.460 2234.595 3386.110 2234.845 ;
        RECT 3385.940 2234.555 3386.110 2234.595 ;
      LAYER li1 ;
        RECT 3385.120 2234.255 3385.770 2234.425 ;
      LAYER li1 ;
        RECT 3385.940 2234.095 3386.110 2234.385 ;
        RECT 3382.420 2233.835 3384.190 2233.925 ;
        RECT 3382.420 2233.715 3383.390 2233.835 ;
        RECT 3380.500 2233.635 3380.670 2233.715 ;
        RECT 3383.220 2233.635 3383.390 2233.715 ;
        RECT 3384.410 2233.820 3385.290 2233.995 ;
        RECT 3384.410 2233.665 3384.580 2233.820 ;
        RECT 3380.500 2233.205 3380.670 2233.465 ;
        RECT 3383.220 2233.205 3383.390 2233.465 ;
        RECT 3383.560 2233.335 3384.580 2233.665 ;
        RECT 3380.500 2233.175 3381.470 2233.205 ;
        RECT 3380.670 2233.005 3381.470 2233.175 ;
        RECT 3380.500 2232.875 3381.470 2233.005 ;
        RECT 3382.070 2233.175 3383.390 2233.205 ;
        RECT 3382.070 2233.005 3383.220 2233.175 ;
        RECT 3383.390 2233.005 3384.190 2233.165 ;
        RECT 3382.070 2232.995 3384.190 2233.005 ;
        RECT 3382.070 2232.875 3383.390 2232.995 ;
        RECT 3380.500 2232.715 3380.670 2232.875 ;
        RECT 3383.220 2232.715 3383.390 2232.875 ;
        RECT 3384.410 2232.825 3384.580 2233.335 ;
        RECT 3377.780 2232.315 3377.950 2232.400 ;
        RECT 3380.500 2232.315 3380.670 2232.545 ;
        RECT 3383.220 2232.315 3383.390 2232.545 ;
        RECT 3383.560 2232.495 3384.580 2232.825 ;
        RECT 3385.120 2233.585 3385.290 2233.820 ;
        RECT 3385.460 2233.925 3385.940 2234.085 ;
        RECT 3385.460 2233.755 3386.110 2233.925 ;
        RECT 3385.940 2233.635 3386.110 2233.755 ;
        RECT 3385.120 2233.415 3385.765 2233.585 ;
        RECT 3385.120 2232.745 3385.290 2233.415 ;
        RECT 3385.940 2233.245 3386.110 2233.465 ;
        RECT 3385.460 2233.175 3386.110 2233.245 ;
        RECT 3385.460 2233.005 3385.940 2233.175 ;
        RECT 3385.460 2232.915 3386.110 2233.005 ;
        RECT 3385.120 2232.575 3385.770 2232.745 ;
        RECT 3385.940 2232.715 3386.110 2232.915 ;
        RECT 3385.940 2232.315 3386.110 2232.545 ;
        RECT 3377.780 2232.255 3379.115 2232.315 ;
        RECT 3377.950 2232.085 3379.115 2232.255 ;
        RECT 3377.780 2232.025 3379.115 2232.085 ;
        RECT 3379.775 2232.255 3381.395 2232.315 ;
        RECT 3379.775 2232.085 3380.500 2232.255 ;
        RECT 3380.670 2232.085 3381.395 2232.255 ;
        RECT 3379.775 2232.025 3381.395 2232.085 ;
        RECT 3382.055 2232.255 3384.555 2232.315 ;
        RECT 3382.055 2232.085 3383.220 2232.255 ;
        RECT 3383.390 2232.085 3384.555 2232.255 ;
        RECT 3382.055 2232.025 3384.555 2232.085 ;
        RECT 3385.215 2232.255 3386.110 2232.315 ;
        RECT 3385.215 2232.085 3385.940 2232.255 ;
        RECT 3385.215 2232.025 3386.110 2232.085 ;
        RECT 3377.780 2231.940 3377.950 2232.025 ;
      LAYER li1 ;
        RECT 3379.955 2230.270 3380.500 2231.855 ;
      LAYER li1 ;
        RECT 3380.500 2231.795 3380.670 2232.025 ;
        RECT 3380.500 2231.425 3380.670 2231.625 ;
        RECT 3380.840 2231.595 3381.490 2231.765 ;
        RECT 3380.500 2231.335 3381.150 2231.425 ;
        RECT 3380.670 2231.165 3381.150 2231.335 ;
        RECT 3380.500 2231.095 3381.150 2231.165 ;
        RECT 3380.500 2230.875 3380.670 2231.095 ;
        RECT 3381.320 2230.925 3381.490 2231.595 ;
        RECT 3380.845 2230.755 3381.490 2230.925 ;
        RECT 3380.500 2230.585 3380.670 2230.705 ;
        RECT 3380.500 2230.415 3381.150 2230.585 ;
      LAYER li1 ;
        RECT 3379.125 2229.930 3380.500 2230.270 ;
      LAYER li1 ;
        RECT 3380.670 2230.255 3381.150 2230.415 ;
        RECT 3381.320 2230.520 3381.490 2230.755 ;
        RECT 3382.030 2231.515 3383.050 2231.845 ;
        RECT 3383.220 2231.795 3383.390 2232.025 ;
        RECT 3385.940 2231.795 3386.110 2232.025 ;
        RECT 3382.030 2231.005 3382.200 2231.515 ;
        RECT 3383.220 2231.465 3383.390 2231.625 ;
        RECT 3385.940 2231.465 3386.110 2231.625 ;
        RECT 3383.220 2231.345 3384.540 2231.465 ;
        RECT 3382.420 2231.335 3384.540 2231.345 ;
        RECT 3382.420 2231.175 3383.220 2231.335 ;
        RECT 3383.390 2231.165 3384.540 2231.335 ;
        RECT 3383.220 2231.135 3384.540 2231.165 ;
        RECT 3385.140 2231.335 3386.110 2231.465 ;
        RECT 3385.140 2231.165 3385.940 2231.335 ;
        RECT 3385.140 2231.135 3386.110 2231.165 ;
        RECT 3382.030 2230.675 3383.050 2231.005 ;
        RECT 3383.220 2230.875 3383.390 2231.135 ;
        RECT 3385.940 2230.875 3386.110 2231.135 ;
        RECT 3382.030 2230.520 3382.200 2230.675 ;
        RECT 3381.320 2230.345 3382.200 2230.520 ;
        RECT 3383.220 2230.625 3383.390 2230.705 ;
        RECT 3385.940 2230.625 3386.110 2230.705 ;
        RECT 3383.220 2230.505 3384.190 2230.625 ;
        RECT 3382.420 2230.415 3384.190 2230.505 ;
        RECT 3380.500 2229.955 3380.670 2230.245 ;
      LAYER li1 ;
        RECT 3379.955 2226.510 3380.500 2229.930 ;
      LAYER li1 ;
        RECT 3380.500 2229.745 3380.670 2229.785 ;
        RECT 3380.500 2229.495 3381.150 2229.745 ;
        RECT 3380.670 2229.415 3381.150 2229.495 ;
        RECT 3380.500 2229.035 3380.670 2229.325 ;
        RECT 3380.670 2228.865 3381.150 2228.905 ;
        RECT 3380.500 2228.575 3381.150 2228.865 ;
        RECT 3380.500 2228.115 3380.670 2228.405 ;
        RECT 3380.670 2227.945 3381.150 2228.065 ;
        RECT 3380.500 2227.735 3381.150 2227.945 ;
        RECT 3381.660 2227.895 3381.830 2230.345 ;
        RECT 3382.420 2230.335 3383.220 2230.415 ;
        RECT 3383.390 2230.295 3384.190 2230.415 ;
        RECT 3383.220 2229.955 3383.390 2230.245 ;
        RECT 3383.220 2229.745 3384.190 2229.785 ;
        RECT 3382.420 2229.495 3384.190 2229.745 ;
        RECT 3382.420 2229.415 3383.220 2229.495 ;
        RECT 3383.390 2229.455 3384.190 2229.495 ;
        RECT 3383.220 2229.035 3383.390 2229.325 ;
        RECT 3382.420 2228.865 3383.220 2228.905 ;
        RECT 3383.390 2228.865 3384.190 2228.945 ;
        RECT 3382.420 2228.615 3384.190 2228.865 ;
        RECT 3382.420 2228.575 3383.390 2228.615 ;
        RECT 3383.220 2228.115 3383.390 2228.405 ;
        RECT 3382.420 2227.945 3383.220 2228.065 ;
        RECT 3383.390 2227.945 3384.190 2228.025 ;
        RECT 3384.780 2228.015 3384.950 2230.465 ;
        RECT 3385.460 2230.415 3386.110 2230.625 ;
        RECT 3385.460 2230.295 3385.940 2230.415 ;
        RECT 3385.940 2229.955 3386.110 2230.245 ;
        RECT 3385.460 2229.495 3386.110 2229.785 ;
        RECT 3385.460 2229.455 3385.940 2229.495 ;
        RECT 3385.940 2229.035 3386.110 2229.325 ;
        RECT 3385.460 2228.865 3385.940 2228.945 ;
        RECT 3385.460 2228.615 3386.110 2228.865 ;
        RECT 3385.940 2228.575 3386.110 2228.615 ;
        RECT 3385.940 2228.115 3386.110 2228.405 ;
        RECT 3382.420 2227.855 3384.190 2227.945 ;
        RECT 3382.420 2227.735 3383.390 2227.855 ;
        RECT 3380.500 2227.655 3380.670 2227.735 ;
        RECT 3383.220 2227.655 3383.390 2227.735 ;
        RECT 3384.410 2227.840 3385.290 2228.015 ;
        RECT 3384.410 2227.685 3384.580 2227.840 ;
        RECT 3380.500 2227.225 3380.670 2227.485 ;
        RECT 3383.220 2227.225 3383.390 2227.485 ;
        RECT 3383.560 2227.355 3384.580 2227.685 ;
        RECT 3380.500 2227.195 3381.470 2227.225 ;
        RECT 3380.670 2227.025 3381.470 2227.195 ;
        RECT 3380.500 2226.895 3381.470 2227.025 ;
        RECT 3382.070 2227.195 3383.390 2227.225 ;
        RECT 3382.070 2227.025 3383.220 2227.195 ;
        RECT 3383.390 2227.025 3384.190 2227.185 ;
        RECT 3382.070 2227.015 3384.190 2227.025 ;
        RECT 3382.070 2226.895 3383.390 2227.015 ;
        RECT 3380.500 2226.735 3380.670 2226.895 ;
        RECT 3383.220 2226.735 3383.390 2226.895 ;
        RECT 3384.410 2226.845 3384.580 2227.355 ;
        RECT 3377.780 2226.335 3377.950 2226.420 ;
        RECT 3380.500 2226.335 3380.670 2226.565 ;
        RECT 3383.220 2226.335 3383.390 2226.565 ;
        RECT 3383.560 2226.515 3384.580 2226.845 ;
        RECT 3385.120 2227.605 3385.290 2227.840 ;
        RECT 3385.460 2227.945 3385.940 2228.105 ;
        RECT 3385.460 2227.775 3386.110 2227.945 ;
        RECT 3385.940 2227.655 3386.110 2227.775 ;
        RECT 3385.120 2227.435 3385.765 2227.605 ;
        RECT 3385.120 2226.765 3385.290 2227.435 ;
        RECT 3385.940 2227.265 3386.110 2227.485 ;
        RECT 3385.460 2227.195 3386.110 2227.265 ;
        RECT 3385.460 2227.025 3385.940 2227.195 ;
        RECT 3385.460 2226.935 3386.110 2227.025 ;
        RECT 3385.120 2226.595 3385.770 2226.765 ;
        RECT 3385.940 2226.735 3386.110 2226.935 ;
        RECT 3385.940 2226.335 3386.110 2226.565 ;
        RECT 3377.780 2226.275 3379.115 2226.335 ;
        RECT 3377.950 2226.105 3379.115 2226.275 ;
        RECT 3377.780 2226.045 3379.115 2226.105 ;
        RECT 3379.775 2226.275 3381.395 2226.335 ;
        RECT 3379.775 2226.105 3380.500 2226.275 ;
        RECT 3380.670 2226.105 3381.395 2226.275 ;
        RECT 3379.775 2226.045 3381.395 2226.105 ;
        RECT 3382.055 2226.275 3384.555 2226.335 ;
        RECT 3382.055 2226.105 3383.220 2226.275 ;
        RECT 3383.390 2226.105 3384.555 2226.275 ;
        RECT 3382.055 2226.045 3384.555 2226.105 ;
        RECT 3385.215 2226.275 3386.110 2226.335 ;
        RECT 3385.215 2226.105 3385.940 2226.275 ;
        RECT 3385.215 2226.045 3386.110 2226.105 ;
        RECT 3377.780 2225.960 3377.950 2226.045 ;
      LAYER li1 ;
        RECT 3379.955 2224.290 3380.500 2225.875 ;
      LAYER li1 ;
        RECT 3380.500 2225.815 3380.670 2226.045 ;
        RECT 3380.500 2225.445 3380.670 2225.645 ;
        RECT 3380.840 2225.615 3381.490 2225.785 ;
        RECT 3380.500 2225.355 3381.150 2225.445 ;
        RECT 3380.670 2225.185 3381.150 2225.355 ;
        RECT 3380.500 2225.115 3381.150 2225.185 ;
        RECT 3380.500 2224.895 3380.670 2225.115 ;
        RECT 3381.320 2224.945 3381.490 2225.615 ;
        RECT 3380.845 2224.775 3381.490 2224.945 ;
        RECT 3380.500 2224.605 3380.670 2224.725 ;
        RECT 3380.500 2224.435 3381.150 2224.605 ;
      LAYER li1 ;
        RECT 3379.125 2223.950 3380.500 2224.290 ;
      LAYER li1 ;
        RECT 3380.670 2224.275 3381.150 2224.435 ;
        RECT 3381.320 2224.540 3381.490 2224.775 ;
        RECT 3382.030 2225.535 3383.050 2225.865 ;
        RECT 3383.220 2225.815 3383.390 2226.045 ;
        RECT 3385.940 2225.815 3386.110 2226.045 ;
        RECT 3382.030 2225.025 3382.200 2225.535 ;
        RECT 3383.220 2225.485 3383.390 2225.645 ;
        RECT 3385.940 2225.485 3386.110 2225.645 ;
        RECT 3383.220 2225.365 3384.540 2225.485 ;
        RECT 3382.420 2225.355 3384.540 2225.365 ;
        RECT 3382.420 2225.195 3383.220 2225.355 ;
        RECT 3383.390 2225.185 3384.540 2225.355 ;
        RECT 3383.220 2225.155 3384.540 2225.185 ;
        RECT 3385.140 2225.355 3386.110 2225.485 ;
        RECT 3385.140 2225.185 3385.940 2225.355 ;
        RECT 3385.140 2225.155 3386.110 2225.185 ;
        RECT 3382.030 2224.695 3383.050 2225.025 ;
        RECT 3383.220 2224.895 3383.390 2225.155 ;
        RECT 3385.940 2224.895 3386.110 2225.155 ;
        RECT 3382.030 2224.540 3382.200 2224.695 ;
        RECT 3381.320 2224.365 3382.200 2224.540 ;
        RECT 3383.220 2224.645 3383.390 2224.725 ;
        RECT 3385.940 2224.645 3386.110 2224.725 ;
        RECT 3383.220 2224.525 3384.190 2224.645 ;
        RECT 3382.420 2224.435 3384.190 2224.525 ;
        RECT 3380.500 2223.975 3380.670 2224.265 ;
      LAYER li1 ;
        RECT 3379.955 2220.530 3380.500 2223.950 ;
      LAYER li1 ;
        RECT 3380.500 2223.765 3380.670 2223.805 ;
        RECT 3380.500 2223.515 3381.150 2223.765 ;
        RECT 3380.670 2223.435 3381.150 2223.515 ;
        RECT 3380.500 2223.055 3380.670 2223.345 ;
        RECT 3380.670 2222.885 3381.150 2222.925 ;
        RECT 3380.500 2222.595 3381.150 2222.885 ;
        RECT 3380.500 2222.135 3380.670 2222.425 ;
        RECT 3380.670 2221.965 3381.150 2222.085 ;
        RECT 3380.500 2221.755 3381.150 2221.965 ;
        RECT 3381.660 2221.915 3381.830 2224.365 ;
        RECT 3382.420 2224.355 3383.220 2224.435 ;
        RECT 3383.390 2224.315 3384.190 2224.435 ;
        RECT 3383.220 2223.975 3383.390 2224.265 ;
        RECT 3383.220 2223.765 3384.190 2223.805 ;
        RECT 3382.420 2223.515 3384.190 2223.765 ;
        RECT 3382.420 2223.435 3383.220 2223.515 ;
        RECT 3383.390 2223.475 3384.190 2223.515 ;
        RECT 3383.220 2223.055 3383.390 2223.345 ;
        RECT 3382.420 2222.885 3383.220 2222.925 ;
        RECT 3383.390 2222.885 3384.190 2222.965 ;
        RECT 3382.420 2222.635 3384.190 2222.885 ;
        RECT 3382.420 2222.595 3383.390 2222.635 ;
        RECT 3383.220 2222.135 3383.390 2222.425 ;
        RECT 3382.420 2221.965 3383.220 2222.085 ;
        RECT 3383.390 2221.965 3384.190 2222.045 ;
        RECT 3384.780 2222.035 3384.950 2224.485 ;
        RECT 3385.460 2224.435 3386.110 2224.645 ;
        RECT 3385.460 2224.315 3385.940 2224.435 ;
        RECT 3385.940 2223.975 3386.110 2224.265 ;
        RECT 3385.460 2223.515 3386.110 2223.805 ;
        RECT 3385.460 2223.475 3385.940 2223.515 ;
        RECT 3385.940 2223.055 3386.110 2223.345 ;
        RECT 3385.460 2222.885 3385.940 2222.965 ;
        RECT 3385.460 2222.635 3386.110 2222.885 ;
        RECT 3385.940 2222.595 3386.110 2222.635 ;
        RECT 3385.940 2222.135 3386.110 2222.425 ;
        RECT 3382.420 2221.875 3384.190 2221.965 ;
        RECT 3382.420 2221.755 3383.390 2221.875 ;
        RECT 3380.500 2221.675 3380.670 2221.755 ;
        RECT 3383.220 2221.675 3383.390 2221.755 ;
        RECT 3384.410 2221.860 3385.290 2222.035 ;
        RECT 3384.410 2221.705 3384.580 2221.860 ;
        RECT 3380.500 2221.245 3380.670 2221.505 ;
        RECT 3383.220 2221.245 3383.390 2221.505 ;
        RECT 3383.560 2221.375 3384.580 2221.705 ;
        RECT 3380.500 2221.215 3381.470 2221.245 ;
        RECT 3380.670 2221.045 3381.470 2221.215 ;
        RECT 3380.500 2220.915 3381.470 2221.045 ;
        RECT 3382.070 2221.215 3383.390 2221.245 ;
        RECT 3382.070 2221.045 3383.220 2221.215 ;
        RECT 3383.390 2221.045 3384.190 2221.205 ;
        RECT 3382.070 2221.035 3384.190 2221.045 ;
        RECT 3382.070 2220.915 3383.390 2221.035 ;
        RECT 3380.500 2220.755 3380.670 2220.915 ;
        RECT 3383.220 2220.755 3383.390 2220.915 ;
        RECT 3384.410 2220.865 3384.580 2221.375 ;
        RECT 3377.780 2220.355 3377.950 2220.440 ;
        RECT 3380.500 2220.355 3380.670 2220.585 ;
        RECT 3383.220 2220.355 3383.390 2220.585 ;
        RECT 3383.560 2220.535 3384.580 2220.865 ;
        RECT 3385.120 2221.625 3385.290 2221.860 ;
        RECT 3385.460 2221.965 3385.940 2222.125 ;
        RECT 3385.460 2221.795 3386.110 2221.965 ;
        RECT 3385.940 2221.675 3386.110 2221.795 ;
        RECT 3385.120 2221.455 3385.765 2221.625 ;
        RECT 3385.120 2220.785 3385.290 2221.455 ;
        RECT 3385.940 2221.285 3386.110 2221.505 ;
        RECT 3385.460 2221.215 3386.110 2221.285 ;
        RECT 3385.460 2221.045 3385.940 2221.215 ;
        RECT 3385.460 2220.955 3386.110 2221.045 ;
        RECT 3385.120 2220.615 3385.770 2220.785 ;
        RECT 3385.940 2220.755 3386.110 2220.955 ;
        RECT 3385.940 2220.355 3386.110 2220.585 ;
        RECT 3377.780 2220.295 3379.115 2220.355 ;
        RECT 3377.950 2220.125 3379.115 2220.295 ;
        RECT 3377.780 2220.065 3379.115 2220.125 ;
        RECT 3379.775 2220.295 3381.395 2220.355 ;
        RECT 3379.775 2220.125 3380.500 2220.295 ;
        RECT 3380.670 2220.125 3381.395 2220.295 ;
        RECT 3379.775 2220.065 3381.395 2220.125 ;
        RECT 3382.055 2220.295 3384.555 2220.355 ;
        RECT 3382.055 2220.125 3383.220 2220.295 ;
        RECT 3383.390 2220.125 3384.555 2220.295 ;
        RECT 3382.055 2220.065 3384.555 2220.125 ;
        RECT 3385.215 2220.295 3386.110 2220.355 ;
        RECT 3385.215 2220.125 3385.940 2220.295 ;
        RECT 3385.215 2220.065 3386.110 2220.125 ;
        RECT 3377.780 2219.980 3377.950 2220.065 ;
      LAYER li1 ;
        RECT 3379.955 2218.310 3380.500 2219.895 ;
      LAYER li1 ;
        RECT 3380.500 2219.835 3380.670 2220.065 ;
        RECT 3380.500 2219.465 3380.670 2219.665 ;
        RECT 3380.840 2219.635 3381.490 2219.805 ;
        RECT 3380.500 2219.375 3381.150 2219.465 ;
        RECT 3380.670 2219.205 3381.150 2219.375 ;
        RECT 3380.500 2219.135 3381.150 2219.205 ;
        RECT 3380.500 2218.915 3380.670 2219.135 ;
        RECT 3381.320 2218.965 3381.490 2219.635 ;
        RECT 3380.845 2218.795 3381.490 2218.965 ;
        RECT 3380.500 2218.625 3380.670 2218.745 ;
        RECT 3380.500 2218.455 3381.150 2218.625 ;
      LAYER li1 ;
        RECT 3379.125 2217.970 3380.500 2218.310 ;
      LAYER li1 ;
        RECT 3380.670 2218.295 3381.150 2218.455 ;
        RECT 3381.320 2218.560 3381.490 2218.795 ;
        RECT 3382.030 2219.555 3383.050 2219.885 ;
        RECT 3383.220 2219.835 3383.390 2220.065 ;
        RECT 3385.940 2219.835 3386.110 2220.065 ;
        RECT 3382.030 2219.045 3382.200 2219.555 ;
        RECT 3383.220 2219.505 3383.390 2219.665 ;
        RECT 3385.940 2219.505 3386.110 2219.665 ;
        RECT 3383.220 2219.385 3384.540 2219.505 ;
        RECT 3382.420 2219.375 3384.540 2219.385 ;
        RECT 3382.420 2219.215 3383.220 2219.375 ;
        RECT 3383.390 2219.205 3384.540 2219.375 ;
        RECT 3383.220 2219.175 3384.540 2219.205 ;
        RECT 3385.140 2219.375 3386.110 2219.505 ;
        RECT 3385.140 2219.205 3385.940 2219.375 ;
        RECT 3385.140 2219.175 3386.110 2219.205 ;
        RECT 3382.030 2218.715 3383.050 2219.045 ;
        RECT 3383.220 2218.915 3383.390 2219.175 ;
        RECT 3385.940 2218.915 3386.110 2219.175 ;
        RECT 3382.030 2218.560 3382.200 2218.715 ;
        RECT 3381.320 2218.385 3382.200 2218.560 ;
        RECT 3383.220 2218.665 3383.390 2218.745 ;
        RECT 3385.940 2218.665 3386.110 2218.745 ;
        RECT 3383.220 2218.545 3384.190 2218.665 ;
        RECT 3382.420 2218.455 3384.190 2218.545 ;
        RECT 3380.500 2217.995 3380.670 2218.285 ;
      LAYER li1 ;
        RECT 3379.955 2214.550 3380.500 2217.970 ;
      LAYER li1 ;
        RECT 3380.500 2217.785 3380.670 2217.825 ;
        RECT 3380.500 2217.535 3381.150 2217.785 ;
        RECT 3380.670 2217.455 3381.150 2217.535 ;
        RECT 3380.500 2217.075 3380.670 2217.365 ;
        RECT 3380.670 2216.905 3381.150 2216.945 ;
        RECT 3380.500 2216.615 3381.150 2216.905 ;
        RECT 3380.500 2216.155 3380.670 2216.445 ;
        RECT 3380.670 2215.985 3381.150 2216.105 ;
        RECT 3380.500 2215.775 3381.150 2215.985 ;
        RECT 3381.660 2215.935 3381.830 2218.385 ;
        RECT 3382.420 2218.375 3383.220 2218.455 ;
        RECT 3383.390 2218.335 3384.190 2218.455 ;
        RECT 3383.220 2217.995 3383.390 2218.285 ;
        RECT 3383.220 2217.785 3384.190 2217.825 ;
        RECT 3382.420 2217.535 3384.190 2217.785 ;
        RECT 3382.420 2217.455 3383.220 2217.535 ;
        RECT 3383.390 2217.495 3384.190 2217.535 ;
        RECT 3383.220 2217.075 3383.390 2217.365 ;
        RECT 3382.420 2216.905 3383.220 2216.945 ;
        RECT 3383.390 2216.905 3384.190 2216.985 ;
        RECT 3382.420 2216.655 3384.190 2216.905 ;
        RECT 3382.420 2216.615 3383.390 2216.655 ;
        RECT 3383.220 2216.155 3383.390 2216.445 ;
        RECT 3382.420 2215.985 3383.220 2216.105 ;
        RECT 3383.390 2215.985 3384.190 2216.065 ;
        RECT 3384.780 2216.055 3384.950 2218.505 ;
        RECT 3385.460 2218.455 3386.110 2218.665 ;
        RECT 3385.460 2218.335 3385.940 2218.455 ;
        RECT 3385.940 2217.995 3386.110 2218.285 ;
        RECT 3385.460 2217.535 3386.110 2217.825 ;
        RECT 3385.460 2217.495 3385.940 2217.535 ;
        RECT 3385.940 2217.075 3386.110 2217.365 ;
        RECT 3385.460 2216.905 3385.940 2216.985 ;
        RECT 3385.460 2216.655 3386.110 2216.905 ;
        RECT 3385.940 2216.615 3386.110 2216.655 ;
        RECT 3385.940 2216.155 3386.110 2216.445 ;
        RECT 3382.420 2215.895 3384.190 2215.985 ;
        RECT 3382.420 2215.775 3383.390 2215.895 ;
        RECT 3380.500 2215.695 3380.670 2215.775 ;
        RECT 3383.220 2215.695 3383.390 2215.775 ;
        RECT 3384.410 2215.880 3385.290 2216.055 ;
        RECT 3384.410 2215.725 3384.580 2215.880 ;
        RECT 3380.500 2215.265 3380.670 2215.525 ;
        RECT 3383.220 2215.265 3383.390 2215.525 ;
        RECT 3383.560 2215.395 3384.580 2215.725 ;
        RECT 3380.500 2215.235 3381.470 2215.265 ;
        RECT 3380.670 2215.065 3381.470 2215.235 ;
        RECT 3380.500 2214.935 3381.470 2215.065 ;
        RECT 3382.070 2215.235 3383.390 2215.265 ;
        RECT 3382.070 2215.065 3383.220 2215.235 ;
        RECT 3383.390 2215.065 3384.190 2215.225 ;
        RECT 3382.070 2215.055 3384.190 2215.065 ;
        RECT 3382.070 2214.935 3383.390 2215.055 ;
        RECT 3380.500 2214.775 3380.670 2214.935 ;
        RECT 3383.220 2214.775 3383.390 2214.935 ;
        RECT 3384.410 2214.885 3384.580 2215.395 ;
        RECT 3377.780 2214.375 3377.950 2214.460 ;
        RECT 3380.500 2214.375 3380.670 2214.605 ;
        RECT 3383.220 2214.375 3383.390 2214.605 ;
        RECT 3383.560 2214.555 3384.580 2214.885 ;
        RECT 3385.120 2215.645 3385.290 2215.880 ;
        RECT 3385.460 2215.985 3385.940 2216.145 ;
        RECT 3385.460 2215.815 3386.110 2215.985 ;
        RECT 3385.940 2215.695 3386.110 2215.815 ;
        RECT 3385.120 2215.475 3385.765 2215.645 ;
        RECT 3385.120 2214.805 3385.290 2215.475 ;
        RECT 3385.940 2215.305 3386.110 2215.525 ;
        RECT 3385.460 2215.235 3386.110 2215.305 ;
        RECT 3385.460 2215.065 3385.940 2215.235 ;
        RECT 3385.460 2214.975 3386.110 2215.065 ;
        RECT 3385.120 2214.635 3385.770 2214.805 ;
        RECT 3385.940 2214.775 3386.110 2214.975 ;
        RECT 3385.940 2214.375 3386.110 2214.605 ;
        RECT 3377.780 2214.315 3379.115 2214.375 ;
        RECT 3377.950 2214.145 3379.115 2214.315 ;
        RECT 3377.780 2214.085 3379.115 2214.145 ;
        RECT 3379.775 2214.315 3381.395 2214.375 ;
        RECT 3379.775 2214.145 3380.500 2214.315 ;
        RECT 3380.670 2214.145 3381.395 2214.315 ;
        RECT 3379.775 2214.085 3381.395 2214.145 ;
        RECT 3382.055 2214.315 3384.555 2214.375 ;
        RECT 3382.055 2214.145 3383.220 2214.315 ;
        RECT 3383.390 2214.145 3384.555 2214.315 ;
        RECT 3382.055 2214.085 3384.555 2214.145 ;
        RECT 3385.215 2214.315 3386.110 2214.375 ;
        RECT 3385.215 2214.145 3385.940 2214.315 ;
        RECT 3385.215 2214.085 3386.110 2214.145 ;
        RECT 3377.780 2214.000 3377.950 2214.085 ;
      LAYER li1 ;
        RECT 3379.955 2212.330 3380.500 2213.915 ;
      LAYER li1 ;
        RECT 3380.500 2213.855 3380.670 2214.085 ;
        RECT 3380.500 2213.485 3380.670 2213.685 ;
        RECT 3380.840 2213.655 3381.490 2213.825 ;
        RECT 3380.500 2213.395 3381.150 2213.485 ;
        RECT 3380.670 2213.225 3381.150 2213.395 ;
        RECT 3380.500 2213.155 3381.150 2213.225 ;
        RECT 3380.500 2212.935 3380.670 2213.155 ;
        RECT 3381.320 2212.985 3381.490 2213.655 ;
        RECT 3380.845 2212.815 3381.490 2212.985 ;
        RECT 3380.500 2212.645 3380.670 2212.765 ;
        RECT 3380.500 2212.475 3381.150 2212.645 ;
      LAYER li1 ;
        RECT 3379.125 2211.990 3380.500 2212.330 ;
      LAYER li1 ;
        RECT 3380.670 2212.315 3381.150 2212.475 ;
        RECT 3381.320 2212.580 3381.490 2212.815 ;
        RECT 3382.030 2213.575 3383.050 2213.905 ;
        RECT 3383.220 2213.855 3383.390 2214.085 ;
        RECT 3385.940 2213.855 3386.110 2214.085 ;
        RECT 3382.030 2213.065 3382.200 2213.575 ;
        RECT 3383.220 2213.525 3383.390 2213.685 ;
        RECT 3385.940 2213.525 3386.110 2213.685 ;
        RECT 3383.220 2213.405 3384.540 2213.525 ;
        RECT 3382.420 2213.395 3384.540 2213.405 ;
        RECT 3382.420 2213.235 3383.220 2213.395 ;
        RECT 3383.390 2213.225 3384.540 2213.395 ;
        RECT 3383.220 2213.195 3384.540 2213.225 ;
        RECT 3385.140 2213.395 3386.110 2213.525 ;
        RECT 3385.140 2213.225 3385.940 2213.395 ;
        RECT 3385.140 2213.195 3386.110 2213.225 ;
        RECT 3382.030 2212.735 3383.050 2213.065 ;
        RECT 3383.220 2212.935 3383.390 2213.195 ;
        RECT 3385.940 2212.935 3386.110 2213.195 ;
        RECT 3382.030 2212.580 3382.200 2212.735 ;
        RECT 3381.320 2212.405 3382.200 2212.580 ;
        RECT 3383.220 2212.685 3383.390 2212.765 ;
        RECT 3385.940 2212.685 3386.110 2212.765 ;
        RECT 3383.220 2212.565 3384.190 2212.685 ;
        RECT 3382.420 2212.475 3384.190 2212.565 ;
        RECT 3380.500 2212.015 3380.670 2212.305 ;
      LAYER li1 ;
        RECT 3379.955 2208.570 3380.500 2211.990 ;
      LAYER li1 ;
        RECT 3380.500 2211.805 3380.670 2211.845 ;
        RECT 3380.500 2211.555 3381.150 2211.805 ;
        RECT 3380.670 2211.475 3381.150 2211.555 ;
        RECT 3380.500 2211.095 3380.670 2211.385 ;
        RECT 3380.670 2210.925 3381.150 2210.965 ;
        RECT 3380.500 2210.635 3381.150 2210.925 ;
        RECT 3380.500 2210.175 3380.670 2210.465 ;
        RECT 3380.670 2210.005 3381.150 2210.125 ;
        RECT 3380.500 2209.795 3381.150 2210.005 ;
        RECT 3381.660 2209.955 3381.830 2212.405 ;
        RECT 3382.420 2212.395 3383.220 2212.475 ;
        RECT 3383.390 2212.355 3384.190 2212.475 ;
        RECT 3383.220 2212.015 3383.390 2212.305 ;
        RECT 3383.220 2211.805 3384.190 2211.845 ;
        RECT 3382.420 2211.555 3384.190 2211.805 ;
        RECT 3382.420 2211.475 3383.220 2211.555 ;
        RECT 3383.390 2211.515 3384.190 2211.555 ;
        RECT 3383.220 2211.095 3383.390 2211.385 ;
        RECT 3382.420 2210.925 3383.220 2210.965 ;
        RECT 3383.390 2210.925 3384.190 2211.005 ;
        RECT 3382.420 2210.675 3384.190 2210.925 ;
        RECT 3382.420 2210.635 3383.390 2210.675 ;
        RECT 3383.220 2210.175 3383.390 2210.465 ;
        RECT 3382.420 2210.005 3383.220 2210.125 ;
        RECT 3383.390 2210.005 3384.190 2210.085 ;
        RECT 3384.780 2210.075 3384.950 2212.525 ;
        RECT 3385.460 2212.475 3386.110 2212.685 ;
        RECT 3385.460 2212.355 3385.940 2212.475 ;
        RECT 3385.940 2212.015 3386.110 2212.305 ;
        RECT 3385.460 2211.555 3386.110 2211.845 ;
        RECT 3385.460 2211.515 3385.940 2211.555 ;
        RECT 3385.940 2211.095 3386.110 2211.385 ;
        RECT 3385.460 2210.925 3385.940 2211.005 ;
        RECT 3385.460 2210.675 3386.110 2210.925 ;
        RECT 3385.940 2210.635 3386.110 2210.675 ;
        RECT 3385.940 2210.175 3386.110 2210.465 ;
        RECT 3382.420 2209.915 3384.190 2210.005 ;
        RECT 3382.420 2209.795 3383.390 2209.915 ;
        RECT 3380.500 2209.715 3380.670 2209.795 ;
        RECT 3383.220 2209.715 3383.390 2209.795 ;
        RECT 3384.410 2209.900 3385.290 2210.075 ;
        RECT 3384.410 2209.745 3384.580 2209.900 ;
        RECT 3380.500 2209.285 3380.670 2209.545 ;
        RECT 3383.220 2209.285 3383.390 2209.545 ;
        RECT 3383.560 2209.415 3384.580 2209.745 ;
        RECT 3380.500 2209.255 3381.470 2209.285 ;
        RECT 3380.670 2209.085 3381.470 2209.255 ;
        RECT 3380.500 2208.955 3381.470 2209.085 ;
        RECT 3382.070 2209.255 3383.390 2209.285 ;
        RECT 3382.070 2209.085 3383.220 2209.255 ;
        RECT 3383.390 2209.085 3384.190 2209.245 ;
        RECT 3382.070 2209.075 3384.190 2209.085 ;
        RECT 3382.070 2208.955 3383.390 2209.075 ;
        RECT 3380.500 2208.795 3380.670 2208.955 ;
        RECT 3383.220 2208.795 3383.390 2208.955 ;
        RECT 3384.410 2208.905 3384.580 2209.415 ;
        RECT 3377.780 2208.395 3377.950 2208.480 ;
        RECT 3380.500 2208.395 3380.670 2208.625 ;
        RECT 3383.220 2208.395 3383.390 2208.625 ;
        RECT 3383.560 2208.575 3384.580 2208.905 ;
        RECT 3385.120 2209.665 3385.290 2209.900 ;
        RECT 3385.460 2210.005 3385.940 2210.165 ;
        RECT 3385.460 2209.835 3386.110 2210.005 ;
        RECT 3385.940 2209.715 3386.110 2209.835 ;
        RECT 3385.120 2209.495 3385.765 2209.665 ;
        RECT 3385.120 2208.825 3385.290 2209.495 ;
        RECT 3385.940 2209.325 3386.110 2209.545 ;
        RECT 3385.460 2209.255 3386.110 2209.325 ;
        RECT 3385.460 2209.085 3385.940 2209.255 ;
        RECT 3385.460 2208.995 3386.110 2209.085 ;
        RECT 3385.120 2208.655 3385.770 2208.825 ;
        RECT 3385.940 2208.795 3386.110 2208.995 ;
        RECT 3385.940 2208.395 3386.110 2208.625 ;
        RECT 3377.780 2208.335 3379.115 2208.395 ;
        RECT 3377.950 2208.165 3379.115 2208.335 ;
        RECT 3377.780 2208.105 3379.115 2208.165 ;
        RECT 3379.775 2208.335 3381.395 2208.395 ;
        RECT 3379.775 2208.165 3380.500 2208.335 ;
        RECT 3380.670 2208.165 3381.395 2208.335 ;
        RECT 3379.775 2208.105 3381.395 2208.165 ;
        RECT 3382.055 2208.335 3384.555 2208.395 ;
        RECT 3382.055 2208.165 3383.220 2208.335 ;
        RECT 3383.390 2208.165 3384.555 2208.335 ;
        RECT 3382.055 2208.105 3384.555 2208.165 ;
        RECT 3385.215 2208.335 3386.110 2208.395 ;
        RECT 3385.215 2208.165 3385.940 2208.335 ;
        RECT 3385.215 2208.105 3386.110 2208.165 ;
        RECT 3377.780 2208.020 3377.950 2208.105 ;
      LAYER li1 ;
        RECT 3379.955 2206.350 3380.500 2207.935 ;
      LAYER li1 ;
        RECT 3380.500 2207.875 3380.670 2208.105 ;
        RECT 3380.500 2207.505 3380.670 2207.705 ;
        RECT 3380.840 2207.675 3381.490 2207.845 ;
        RECT 3380.500 2207.415 3381.150 2207.505 ;
        RECT 3380.670 2207.245 3381.150 2207.415 ;
        RECT 3380.500 2207.175 3381.150 2207.245 ;
        RECT 3380.500 2206.955 3380.670 2207.175 ;
        RECT 3381.320 2207.005 3381.490 2207.675 ;
        RECT 3380.845 2206.835 3381.490 2207.005 ;
        RECT 3380.500 2206.665 3380.670 2206.785 ;
        RECT 3380.500 2206.495 3381.150 2206.665 ;
      LAYER li1 ;
        RECT 3379.125 2206.010 3380.500 2206.350 ;
      LAYER li1 ;
        RECT 3380.670 2206.335 3381.150 2206.495 ;
        RECT 3381.320 2206.600 3381.490 2206.835 ;
        RECT 3382.030 2207.595 3383.050 2207.925 ;
        RECT 3383.220 2207.875 3383.390 2208.105 ;
        RECT 3385.940 2207.875 3386.110 2208.105 ;
        RECT 3382.030 2207.085 3382.200 2207.595 ;
        RECT 3383.220 2207.545 3383.390 2207.705 ;
        RECT 3385.940 2207.545 3386.110 2207.705 ;
        RECT 3383.220 2207.425 3384.540 2207.545 ;
        RECT 3382.420 2207.415 3384.540 2207.425 ;
        RECT 3382.420 2207.255 3383.220 2207.415 ;
        RECT 3383.390 2207.245 3384.540 2207.415 ;
        RECT 3383.220 2207.215 3384.540 2207.245 ;
        RECT 3385.140 2207.415 3386.110 2207.545 ;
        RECT 3385.140 2207.245 3385.940 2207.415 ;
        RECT 3385.140 2207.215 3386.110 2207.245 ;
        RECT 3382.030 2206.755 3383.050 2207.085 ;
        RECT 3383.220 2206.955 3383.390 2207.215 ;
        RECT 3385.940 2206.955 3386.110 2207.215 ;
        RECT 3382.030 2206.600 3382.200 2206.755 ;
        RECT 3381.320 2206.425 3382.200 2206.600 ;
        RECT 3383.220 2206.705 3383.390 2206.785 ;
        RECT 3385.940 2206.705 3386.110 2206.785 ;
        RECT 3383.220 2206.585 3384.190 2206.705 ;
        RECT 3382.420 2206.495 3384.190 2206.585 ;
        RECT 3380.500 2206.035 3380.670 2206.325 ;
      LAYER li1 ;
        RECT 3379.955 2202.590 3380.500 2206.010 ;
      LAYER li1 ;
        RECT 3380.500 2205.825 3380.670 2205.865 ;
        RECT 3380.500 2205.575 3381.150 2205.825 ;
        RECT 3380.670 2205.495 3381.150 2205.575 ;
        RECT 3380.500 2205.115 3380.670 2205.405 ;
        RECT 3380.670 2204.945 3381.150 2204.985 ;
        RECT 3380.500 2204.655 3381.150 2204.945 ;
        RECT 3380.500 2204.195 3380.670 2204.485 ;
        RECT 3380.670 2204.025 3381.150 2204.145 ;
        RECT 3380.500 2203.815 3381.150 2204.025 ;
        RECT 3381.660 2203.975 3381.830 2206.425 ;
        RECT 3382.420 2206.415 3383.220 2206.495 ;
        RECT 3383.390 2206.375 3384.190 2206.495 ;
        RECT 3383.220 2206.035 3383.390 2206.325 ;
        RECT 3383.220 2205.825 3384.190 2205.865 ;
        RECT 3382.420 2205.575 3384.190 2205.825 ;
        RECT 3382.420 2205.495 3383.220 2205.575 ;
        RECT 3383.390 2205.535 3384.190 2205.575 ;
        RECT 3383.220 2205.115 3383.390 2205.405 ;
        RECT 3382.420 2204.945 3383.220 2204.985 ;
        RECT 3383.390 2204.945 3384.190 2205.025 ;
        RECT 3382.420 2204.695 3384.190 2204.945 ;
        RECT 3382.420 2204.655 3383.390 2204.695 ;
        RECT 3383.220 2204.195 3383.390 2204.485 ;
        RECT 3382.420 2204.025 3383.220 2204.145 ;
        RECT 3383.390 2204.025 3384.190 2204.105 ;
        RECT 3384.780 2204.095 3384.950 2206.545 ;
        RECT 3385.460 2206.495 3386.110 2206.705 ;
        RECT 3385.460 2206.375 3385.940 2206.495 ;
        RECT 3385.940 2206.035 3386.110 2206.325 ;
        RECT 3385.460 2205.575 3386.110 2205.865 ;
        RECT 3385.460 2205.535 3385.940 2205.575 ;
        RECT 3385.940 2205.115 3386.110 2205.405 ;
        RECT 3385.460 2204.945 3385.940 2205.025 ;
        RECT 3385.460 2204.695 3386.110 2204.945 ;
        RECT 3385.940 2204.655 3386.110 2204.695 ;
        RECT 3385.940 2204.195 3386.110 2204.485 ;
        RECT 3382.420 2203.935 3384.190 2204.025 ;
        RECT 3382.420 2203.815 3383.390 2203.935 ;
        RECT 3380.500 2203.735 3380.670 2203.815 ;
        RECT 3383.220 2203.735 3383.390 2203.815 ;
        RECT 3384.410 2203.920 3385.290 2204.095 ;
        RECT 3384.410 2203.765 3384.580 2203.920 ;
        RECT 3380.500 2203.305 3380.670 2203.565 ;
        RECT 3383.220 2203.305 3383.390 2203.565 ;
        RECT 3383.560 2203.435 3384.580 2203.765 ;
        RECT 3380.500 2203.275 3381.470 2203.305 ;
        RECT 3380.670 2203.105 3381.470 2203.275 ;
        RECT 3380.500 2202.975 3381.470 2203.105 ;
        RECT 3382.070 2203.275 3383.390 2203.305 ;
        RECT 3382.070 2203.105 3383.220 2203.275 ;
        RECT 3383.390 2203.105 3384.190 2203.265 ;
        RECT 3382.070 2203.095 3384.190 2203.105 ;
        RECT 3382.070 2202.975 3383.390 2203.095 ;
        RECT 3380.500 2202.815 3380.670 2202.975 ;
        RECT 3383.220 2202.815 3383.390 2202.975 ;
        RECT 3384.410 2202.925 3384.580 2203.435 ;
        RECT 3377.780 2202.415 3377.950 2202.500 ;
        RECT 3380.500 2202.415 3380.670 2202.645 ;
        RECT 3383.220 2202.415 3383.390 2202.645 ;
        RECT 3383.560 2202.595 3384.580 2202.925 ;
        RECT 3385.120 2203.685 3385.290 2203.920 ;
        RECT 3385.460 2204.025 3385.940 2204.185 ;
        RECT 3385.460 2203.855 3386.110 2204.025 ;
        RECT 3385.940 2203.735 3386.110 2203.855 ;
        RECT 3385.120 2203.515 3385.765 2203.685 ;
        RECT 3385.120 2202.845 3385.290 2203.515 ;
        RECT 3385.940 2203.345 3386.110 2203.565 ;
        RECT 3385.460 2203.275 3386.110 2203.345 ;
        RECT 3385.460 2203.105 3385.940 2203.275 ;
        RECT 3385.460 2203.015 3386.110 2203.105 ;
        RECT 3385.120 2202.675 3385.770 2202.845 ;
        RECT 3385.940 2202.815 3386.110 2203.015 ;
        RECT 3385.940 2202.415 3386.110 2202.645 ;
        RECT 3377.780 2202.355 3379.115 2202.415 ;
        RECT 3377.950 2202.185 3379.115 2202.355 ;
        RECT 3377.780 2202.125 3379.115 2202.185 ;
        RECT 3379.775 2202.355 3381.395 2202.415 ;
        RECT 3379.775 2202.185 3380.500 2202.355 ;
        RECT 3380.670 2202.185 3381.395 2202.355 ;
        RECT 3379.775 2202.125 3381.395 2202.185 ;
        RECT 3382.055 2202.355 3384.555 2202.415 ;
        RECT 3382.055 2202.185 3383.220 2202.355 ;
        RECT 3383.390 2202.185 3384.555 2202.355 ;
        RECT 3382.055 2202.125 3384.555 2202.185 ;
        RECT 3385.215 2202.355 3386.110 2202.415 ;
        RECT 3385.215 2202.185 3385.940 2202.355 ;
        RECT 3385.215 2202.125 3386.110 2202.185 ;
        RECT 3377.780 2202.040 3377.950 2202.125 ;
        RECT 3380.500 2202.040 3380.670 2202.125 ;
        RECT 3380.840 2201.695 3381.490 2201.865 ;
        RECT 3380.670 2201.195 3381.150 2201.525 ;
        RECT 3381.320 2201.025 3381.490 2201.695 ;
        RECT 3380.845 2200.855 3381.490 2201.025 ;
        RECT 3380.670 2200.355 3381.150 2200.685 ;
        RECT 3381.320 2200.620 3381.490 2200.855 ;
        RECT 3382.030 2201.615 3383.050 2201.945 ;
        RECT 3383.220 2201.895 3383.390 2202.125 ;
        RECT 3385.940 2201.895 3386.110 2202.125 ;
        RECT 3382.030 2201.105 3382.200 2201.615 ;
        RECT 3383.220 2201.565 3383.390 2201.725 ;
        RECT 3385.940 2201.565 3386.110 2201.725 ;
        RECT 3383.220 2201.445 3384.540 2201.565 ;
        RECT 3382.420 2201.435 3384.540 2201.445 ;
        RECT 3382.420 2201.275 3383.220 2201.435 ;
        RECT 3383.390 2201.265 3384.540 2201.435 ;
        RECT 3383.220 2201.235 3384.540 2201.265 ;
        RECT 3385.140 2201.435 3386.110 2201.565 ;
        RECT 3385.140 2201.265 3385.940 2201.435 ;
        RECT 3385.140 2201.235 3386.110 2201.265 ;
        RECT 3382.030 2200.775 3383.050 2201.105 ;
        RECT 3383.220 2200.975 3383.390 2201.235 ;
        RECT 3385.940 2200.975 3386.110 2201.235 ;
        RECT 3382.030 2200.620 3382.200 2200.775 ;
        RECT 3381.320 2200.445 3382.200 2200.620 ;
        RECT 3383.220 2200.725 3383.390 2200.805 ;
        RECT 3385.940 2200.725 3386.110 2200.805 ;
        RECT 3383.220 2200.605 3384.190 2200.725 ;
        RECT 3382.420 2200.515 3384.190 2200.605 ;
        RECT 3380.670 2199.515 3381.150 2199.845 ;
        RECT 3380.670 2198.675 3381.150 2199.005 ;
        RECT 3380.670 2197.835 3381.150 2198.165 ;
        RECT 3381.660 2197.995 3381.830 2200.445 ;
        RECT 3382.420 2200.435 3383.220 2200.515 ;
        RECT 3383.390 2200.395 3384.190 2200.515 ;
        RECT 3383.220 2200.055 3383.390 2200.345 ;
        RECT 3383.220 2199.845 3384.190 2199.885 ;
        RECT 3382.420 2199.595 3384.190 2199.845 ;
        RECT 3382.420 2199.515 3383.220 2199.595 ;
        RECT 3383.390 2199.555 3384.190 2199.595 ;
        RECT 3383.220 2199.135 3383.390 2199.425 ;
        RECT 3382.420 2198.965 3383.220 2199.005 ;
        RECT 3383.390 2198.965 3384.190 2199.045 ;
        RECT 3382.420 2198.715 3384.190 2198.965 ;
        RECT 3382.420 2198.675 3383.390 2198.715 ;
        RECT 3383.220 2198.215 3383.390 2198.505 ;
        RECT 3382.420 2198.045 3383.220 2198.165 ;
        RECT 3383.390 2198.045 3384.190 2198.125 ;
        RECT 3384.780 2198.115 3384.950 2200.565 ;
        RECT 3385.460 2200.515 3386.110 2200.725 ;
        RECT 3385.460 2200.395 3385.940 2200.515 ;
        RECT 3385.940 2200.055 3386.110 2200.345 ;
        RECT 3385.460 2199.595 3386.110 2199.885 ;
        RECT 3385.460 2199.555 3385.940 2199.595 ;
        RECT 3385.940 2199.135 3386.110 2199.425 ;
        RECT 3385.460 2198.965 3385.940 2199.045 ;
        RECT 3385.460 2198.715 3386.110 2198.965 ;
        RECT 3385.940 2198.675 3386.110 2198.715 ;
        RECT 3385.940 2198.215 3386.110 2198.505 ;
        RECT 3382.420 2197.955 3384.190 2198.045 ;
        RECT 3382.420 2197.835 3383.390 2197.955 ;
        RECT 3383.220 2197.755 3383.390 2197.835 ;
        RECT 3384.410 2197.940 3385.290 2198.115 ;
        RECT 3384.410 2197.785 3384.580 2197.940 ;
        RECT 3383.220 2197.325 3383.390 2197.585 ;
        RECT 3383.560 2197.455 3384.580 2197.785 ;
        RECT 3380.670 2196.995 3381.470 2197.325 ;
        RECT 3382.070 2197.295 3383.390 2197.325 ;
        RECT 3382.070 2197.125 3383.220 2197.295 ;
        RECT 3383.390 2197.125 3384.190 2197.285 ;
        RECT 3382.070 2197.115 3384.190 2197.125 ;
        RECT 3382.070 2196.995 3383.390 2197.115 ;
        RECT 3383.220 2196.835 3383.390 2196.995 ;
        RECT 3384.410 2196.945 3384.580 2197.455 ;
        RECT 3377.780 2196.435 3377.950 2196.520 ;
        RECT 3380.500 2196.435 3380.670 2196.520 ;
        RECT 3383.220 2196.435 3383.390 2196.665 ;
        RECT 3383.560 2196.615 3384.580 2196.945 ;
        RECT 3385.120 2197.705 3385.290 2197.940 ;
        RECT 3385.460 2198.045 3385.940 2198.205 ;
        RECT 3385.460 2197.875 3386.110 2198.045 ;
        RECT 3385.940 2197.755 3386.110 2197.875 ;
        RECT 3385.120 2197.535 3385.765 2197.705 ;
        RECT 3385.120 2196.865 3385.290 2197.535 ;
        RECT 3385.940 2197.365 3386.110 2197.585 ;
        RECT 3385.460 2197.295 3386.110 2197.365 ;
        RECT 3385.460 2197.125 3385.940 2197.295 ;
        RECT 3385.460 2197.035 3386.110 2197.125 ;
        RECT 3385.120 2196.695 3385.770 2196.865 ;
        RECT 3385.940 2196.835 3386.110 2197.035 ;
        RECT 3385.940 2196.435 3386.110 2196.665 ;
        RECT 3377.780 2196.375 3379.115 2196.435 ;
        RECT 3377.950 2196.205 3379.115 2196.375 ;
        RECT 3377.780 2196.145 3379.115 2196.205 ;
        RECT 3379.775 2196.375 3381.395 2196.435 ;
        RECT 3379.775 2196.205 3380.500 2196.375 ;
        RECT 3380.670 2196.205 3381.395 2196.375 ;
        RECT 3379.775 2196.145 3381.395 2196.205 ;
        RECT 3382.055 2196.375 3384.555 2196.435 ;
        RECT 3382.055 2196.205 3383.220 2196.375 ;
        RECT 3383.390 2196.205 3384.555 2196.375 ;
        RECT 3382.055 2196.145 3384.555 2196.205 ;
        RECT 3385.215 2196.375 3386.110 2196.435 ;
        RECT 3385.215 2196.205 3385.940 2196.375 ;
        RECT 3385.215 2196.145 3386.110 2196.205 ;
        RECT 3377.780 2196.060 3377.950 2196.145 ;
        RECT 3380.500 2196.060 3380.670 2196.145 ;
        RECT 3383.220 2196.060 3383.390 2196.145 ;
        RECT 3385.940 2196.060 3386.110 2196.145 ;
        RECT 201.995 1762.980 202.165 1763.065 ;
        RECT 204.715 1762.980 204.885 1763.065 ;
        RECT 207.435 1762.980 207.605 1763.065 ;
        RECT 210.155 1762.980 210.325 1763.065 ;
        RECT 201.995 1762.920 202.890 1762.980 ;
        RECT 202.165 1762.750 202.890 1762.920 ;
        RECT 201.995 1762.690 202.890 1762.750 ;
        RECT 203.550 1762.920 206.050 1762.980 ;
        RECT 203.550 1762.750 204.715 1762.920 ;
        RECT 204.885 1762.750 206.050 1762.920 ;
        RECT 203.550 1762.690 206.050 1762.750 ;
        RECT 201.995 1762.460 202.165 1762.690 ;
        RECT 204.715 1762.460 204.885 1762.690 ;
        RECT 201.995 1762.130 202.165 1762.290 ;
        RECT 204.715 1762.130 204.885 1762.290 ;
        RECT 205.055 1762.180 206.075 1762.510 ;
        RECT 201.995 1762.000 202.965 1762.130 ;
        RECT 202.165 1761.830 202.965 1762.000 ;
        RECT 201.995 1761.800 202.965 1761.830 ;
        RECT 203.565 1762.010 204.885 1762.130 ;
        RECT 203.565 1762.000 205.685 1762.010 ;
        RECT 203.565 1761.830 204.715 1762.000 ;
        RECT 204.885 1761.840 205.685 1762.000 ;
        RECT 203.565 1761.800 204.885 1761.830 ;
        RECT 201.995 1761.540 202.165 1761.800 ;
      LAYER li1 ;
        RECT 202.335 1761.460 204.545 1761.630 ;
      LAYER li1 ;
        RECT 204.715 1761.540 204.885 1761.800 ;
        RECT 205.905 1761.670 206.075 1762.180 ;
      LAYER li1 ;
        RECT 202.815 1761.375 203.695 1761.460 ;
      LAYER li1 ;
        RECT 201.995 1761.290 202.165 1761.370 ;
        RECT 201.995 1761.080 202.645 1761.290 ;
        RECT 202.165 1760.960 202.645 1761.080 ;
        RECT 201.995 1760.620 202.165 1760.910 ;
      LAYER li1 ;
        RECT 202.815 1760.790 202.985 1761.375 ;
        RECT 202.335 1760.620 202.985 1760.790 ;
      LAYER li1 ;
        RECT 201.995 1760.160 202.645 1760.450 ;
        RECT 202.165 1760.120 202.645 1760.160 ;
        RECT 201.995 1759.700 202.165 1759.990 ;
      LAYER li1 ;
        RECT 202.815 1759.950 202.985 1760.620 ;
        RECT 202.335 1759.780 202.985 1759.950 ;
      LAYER li1 ;
        RECT 202.165 1759.530 202.645 1759.610 ;
        RECT 201.995 1759.280 202.645 1759.530 ;
        RECT 201.995 1759.240 202.165 1759.280 ;
      LAYER li1 ;
        RECT 202.815 1759.110 202.985 1759.780 ;
      LAYER li1 ;
        RECT 201.995 1758.780 202.165 1759.070 ;
      LAYER li1 ;
        RECT 202.335 1758.940 202.985 1759.110 ;
      LAYER li1 ;
        RECT 202.165 1758.610 202.645 1758.770 ;
        RECT 203.155 1758.680 203.325 1761.130 ;
      LAYER li1 ;
        RECT 203.525 1760.790 203.695 1761.375 ;
      LAYER li1 ;
        RECT 204.715 1761.290 204.885 1761.370 ;
        RECT 205.055 1761.340 206.075 1761.670 ;
      LAYER li1 ;
        RECT 206.245 1761.365 206.445 1762.955 ;
      LAYER li1 ;
        RECT 206.710 1762.920 208.330 1762.980 ;
        RECT 206.710 1762.750 207.435 1762.920 ;
        RECT 207.605 1762.750 208.330 1762.920 ;
        RECT 206.710 1762.690 208.330 1762.750 ;
        RECT 208.990 1762.920 210.325 1762.980 ;
        RECT 208.990 1762.750 210.155 1762.920 ;
        RECT 208.990 1762.690 210.325 1762.750 ;
        RECT 207.435 1762.605 207.605 1762.690 ;
        RECT 210.155 1762.605 210.325 1762.690 ;
        RECT 206.615 1762.260 207.265 1762.430 ;
        RECT 206.615 1761.590 206.785 1762.260 ;
        RECT 206.955 1761.760 207.435 1762.090 ;
        RECT 206.615 1761.420 207.260 1761.590 ;
        RECT 203.915 1761.170 204.885 1761.290 ;
        RECT 205.905 1761.185 206.075 1761.340 ;
        RECT 206.615 1761.185 206.785 1761.420 ;
        RECT 203.915 1761.080 205.685 1761.170 ;
        RECT 203.915 1760.960 204.715 1761.080 ;
        RECT 204.885 1761.000 205.685 1761.080 ;
        RECT 205.905 1761.010 206.785 1761.185 ;
      LAYER li1 ;
        RECT 203.525 1760.620 204.545 1760.790 ;
      LAYER li1 ;
        RECT 204.715 1760.620 204.885 1760.910 ;
      LAYER li1 ;
        RECT 203.525 1759.950 203.695 1760.620 ;
        RECT 205.055 1760.580 206.075 1760.750 ;
      LAYER li1 ;
        RECT 203.915 1760.410 204.885 1760.450 ;
        RECT 203.915 1760.160 205.685 1760.410 ;
        RECT 203.915 1760.120 204.715 1760.160 ;
        RECT 204.885 1760.080 205.685 1760.160 ;
      LAYER li1 ;
        RECT 203.525 1759.780 204.545 1759.950 ;
        RECT 203.525 1759.110 203.695 1759.780 ;
      LAYER li1 ;
        RECT 204.715 1759.700 204.885 1759.990 ;
      LAYER li1 ;
        RECT 205.905 1759.910 206.075 1760.580 ;
        RECT 205.055 1759.740 206.075 1759.910 ;
      LAYER li1 ;
        RECT 203.915 1759.530 204.715 1759.610 ;
        RECT 204.885 1759.530 205.685 1759.570 ;
        RECT 203.915 1759.280 205.685 1759.530 ;
        RECT 204.715 1759.240 205.685 1759.280 ;
      LAYER li1 ;
        RECT 203.525 1758.940 204.545 1759.110 ;
        RECT 205.905 1759.070 206.075 1759.740 ;
      LAYER li1 ;
        RECT 204.715 1758.780 204.885 1759.070 ;
      LAYER li1 ;
        RECT 205.055 1758.900 206.075 1759.070 ;
      LAYER li1 ;
        RECT 201.995 1758.440 202.645 1758.610 ;
        RECT 202.815 1758.505 203.695 1758.680 ;
        RECT 203.915 1758.610 204.715 1758.690 ;
        RECT 204.885 1758.610 205.685 1758.730 ;
        RECT 203.915 1758.520 205.685 1758.610 ;
        RECT 201.995 1758.320 202.165 1758.440 ;
        RECT 202.815 1758.270 202.985 1758.505 ;
        RECT 203.525 1758.350 203.695 1758.505 ;
        RECT 204.715 1758.400 205.685 1758.520 ;
        RECT 201.995 1757.930 202.165 1758.150 ;
        RECT 202.340 1758.100 202.985 1758.270 ;
        RECT 201.995 1757.860 202.645 1757.930 ;
        RECT 202.165 1757.690 202.645 1757.860 ;
        RECT 201.995 1757.600 202.645 1757.690 ;
        RECT 201.995 1757.400 202.165 1757.600 ;
        RECT 202.815 1757.430 202.985 1758.100 ;
        RECT 202.335 1757.260 202.985 1757.430 ;
        RECT 201.995 1757.000 202.165 1757.230 ;
      LAYER li1 ;
        RECT 203.155 1757.225 203.355 1758.325 ;
      LAYER li1 ;
        RECT 203.525 1758.020 204.545 1758.350 ;
        RECT 204.715 1758.320 204.885 1758.400 ;
      LAYER li1 ;
        RECT 205.905 1758.315 206.075 1758.900 ;
      LAYER li1 ;
        RECT 206.275 1758.560 206.445 1761.010 ;
        RECT 206.955 1760.920 207.435 1761.250 ;
      LAYER li1 ;
        RECT 206.615 1760.580 207.265 1760.750 ;
        RECT 206.615 1759.910 206.785 1760.580 ;
      LAYER li1 ;
        RECT 206.955 1760.080 207.435 1760.410 ;
      LAYER li1 ;
        RECT 206.615 1759.740 207.265 1759.910 ;
        RECT 206.615 1759.070 206.785 1759.740 ;
      LAYER li1 ;
        RECT 206.955 1759.240 207.435 1759.570 ;
      LAYER li1 ;
        RECT 206.615 1758.900 207.265 1759.070 ;
        RECT 206.615 1758.315 206.785 1758.900 ;
      LAYER li1 ;
        RECT 206.955 1758.400 207.435 1758.730 ;
      LAYER li1 ;
        RECT 205.905 1758.230 206.785 1758.315 ;
      LAYER li1 ;
        RECT 203.525 1757.510 203.695 1758.020 ;
        RECT 204.715 1757.890 204.885 1758.150 ;
      LAYER li1 ;
        RECT 205.055 1758.060 207.265 1758.230 ;
      LAYER li1 ;
        RECT 204.715 1757.860 206.035 1757.890 ;
        RECT 203.915 1757.690 204.715 1757.850 ;
        RECT 204.885 1757.690 206.035 1757.860 ;
        RECT 203.915 1757.680 206.035 1757.690 ;
        RECT 204.715 1757.560 206.035 1757.680 ;
        RECT 206.635 1757.560 207.435 1757.890 ;
        RECT 203.525 1757.180 204.545 1757.510 ;
        RECT 204.715 1757.400 204.885 1757.560 ;
        RECT 204.715 1757.000 204.885 1757.230 ;
        RECT 207.435 1757.000 207.605 1757.085 ;
        RECT 210.155 1757.000 210.325 1757.085 ;
        RECT 201.995 1756.940 202.890 1757.000 ;
        RECT 202.165 1756.770 202.890 1756.940 ;
        RECT 201.995 1756.710 202.890 1756.770 ;
        RECT 203.550 1756.940 206.050 1757.000 ;
        RECT 203.550 1756.770 204.715 1756.940 ;
        RECT 204.885 1756.770 206.050 1756.940 ;
        RECT 203.550 1756.710 206.050 1756.770 ;
        RECT 201.995 1756.480 202.165 1756.710 ;
        RECT 204.715 1756.480 204.885 1756.710 ;
        RECT 201.995 1756.150 202.165 1756.310 ;
        RECT 204.715 1756.150 204.885 1756.310 ;
        RECT 205.055 1756.200 206.075 1756.530 ;
        RECT 201.995 1756.020 202.965 1756.150 ;
        RECT 202.165 1755.850 202.965 1756.020 ;
        RECT 201.995 1755.820 202.965 1755.850 ;
        RECT 203.565 1756.030 204.885 1756.150 ;
        RECT 203.565 1756.020 205.685 1756.030 ;
        RECT 203.565 1755.850 204.715 1756.020 ;
        RECT 204.885 1755.860 205.685 1756.020 ;
        RECT 203.565 1755.820 204.885 1755.850 ;
        RECT 201.995 1755.560 202.165 1755.820 ;
      LAYER li1 ;
        RECT 202.335 1755.480 204.545 1755.650 ;
      LAYER li1 ;
        RECT 204.715 1755.560 204.885 1755.820 ;
        RECT 205.905 1755.690 206.075 1756.200 ;
      LAYER li1 ;
        RECT 202.815 1755.395 203.695 1755.480 ;
      LAYER li1 ;
        RECT 201.995 1755.310 202.165 1755.390 ;
        RECT 201.995 1755.100 202.645 1755.310 ;
        RECT 202.165 1754.980 202.645 1755.100 ;
        RECT 201.995 1754.640 202.165 1754.930 ;
      LAYER li1 ;
        RECT 202.815 1754.810 202.985 1755.395 ;
        RECT 202.335 1754.640 202.985 1754.810 ;
      LAYER li1 ;
        RECT 201.995 1754.180 202.645 1754.470 ;
        RECT 202.165 1754.140 202.645 1754.180 ;
        RECT 201.995 1753.720 202.165 1754.010 ;
      LAYER li1 ;
        RECT 202.815 1753.970 202.985 1754.640 ;
        RECT 202.335 1753.800 202.985 1753.970 ;
      LAYER li1 ;
        RECT 202.165 1753.550 202.645 1753.630 ;
        RECT 201.995 1753.300 202.645 1753.550 ;
        RECT 201.995 1753.260 202.165 1753.300 ;
      LAYER li1 ;
        RECT 202.815 1753.130 202.985 1753.800 ;
      LAYER li1 ;
        RECT 201.995 1752.800 202.165 1753.090 ;
      LAYER li1 ;
        RECT 202.335 1752.960 202.985 1753.130 ;
      LAYER li1 ;
        RECT 202.165 1752.630 202.645 1752.790 ;
        RECT 203.155 1752.700 203.325 1755.150 ;
      LAYER li1 ;
        RECT 203.525 1754.810 203.695 1755.395 ;
      LAYER li1 ;
        RECT 204.715 1755.310 204.885 1755.390 ;
        RECT 205.055 1755.360 206.075 1755.690 ;
      LAYER li1 ;
        RECT 206.245 1755.385 206.445 1756.975 ;
      LAYER li1 ;
        RECT 206.710 1756.940 208.330 1757.000 ;
        RECT 206.710 1756.770 207.435 1756.940 ;
        RECT 207.605 1756.770 208.330 1756.940 ;
        RECT 206.710 1756.710 208.330 1756.770 ;
        RECT 208.990 1756.940 210.325 1757.000 ;
        RECT 208.990 1756.770 210.155 1756.940 ;
        RECT 208.990 1756.710 210.325 1756.770 ;
        RECT 207.435 1756.625 207.605 1756.710 ;
        RECT 210.155 1756.625 210.325 1756.710 ;
        RECT 206.615 1756.280 207.265 1756.450 ;
        RECT 206.615 1755.610 206.785 1756.280 ;
        RECT 206.955 1755.780 207.435 1756.110 ;
        RECT 206.615 1755.440 207.260 1755.610 ;
        RECT 203.915 1755.190 204.885 1755.310 ;
        RECT 205.905 1755.205 206.075 1755.360 ;
        RECT 206.615 1755.205 206.785 1755.440 ;
        RECT 203.915 1755.100 205.685 1755.190 ;
        RECT 203.915 1754.980 204.715 1755.100 ;
        RECT 204.885 1755.020 205.685 1755.100 ;
        RECT 205.905 1755.030 206.785 1755.205 ;
      LAYER li1 ;
        RECT 203.525 1754.640 204.545 1754.810 ;
      LAYER li1 ;
        RECT 204.715 1754.640 204.885 1754.930 ;
      LAYER li1 ;
        RECT 203.525 1753.970 203.695 1754.640 ;
        RECT 205.055 1754.600 206.075 1754.770 ;
      LAYER li1 ;
        RECT 203.915 1754.430 204.885 1754.470 ;
        RECT 203.915 1754.180 205.685 1754.430 ;
        RECT 203.915 1754.140 204.715 1754.180 ;
        RECT 204.885 1754.100 205.685 1754.180 ;
      LAYER li1 ;
        RECT 203.525 1753.800 204.545 1753.970 ;
        RECT 203.525 1753.130 203.695 1753.800 ;
      LAYER li1 ;
        RECT 204.715 1753.720 204.885 1754.010 ;
      LAYER li1 ;
        RECT 205.905 1753.930 206.075 1754.600 ;
        RECT 205.055 1753.760 206.075 1753.930 ;
      LAYER li1 ;
        RECT 203.915 1753.550 204.715 1753.630 ;
        RECT 204.885 1753.550 205.685 1753.590 ;
        RECT 203.915 1753.300 205.685 1753.550 ;
        RECT 204.715 1753.260 205.685 1753.300 ;
      LAYER li1 ;
        RECT 203.525 1752.960 204.545 1753.130 ;
        RECT 205.905 1753.090 206.075 1753.760 ;
      LAYER li1 ;
        RECT 204.715 1752.800 204.885 1753.090 ;
      LAYER li1 ;
        RECT 205.055 1752.920 206.075 1753.090 ;
      LAYER li1 ;
        RECT 201.995 1752.460 202.645 1752.630 ;
        RECT 202.815 1752.525 203.695 1752.700 ;
        RECT 203.915 1752.630 204.715 1752.710 ;
        RECT 204.885 1752.630 205.685 1752.750 ;
        RECT 203.915 1752.540 205.685 1752.630 ;
        RECT 201.995 1752.340 202.165 1752.460 ;
        RECT 202.815 1752.290 202.985 1752.525 ;
        RECT 203.525 1752.370 203.695 1752.525 ;
        RECT 204.715 1752.420 205.685 1752.540 ;
        RECT 201.995 1751.950 202.165 1752.170 ;
        RECT 202.340 1752.120 202.985 1752.290 ;
        RECT 201.995 1751.880 202.645 1751.950 ;
        RECT 202.165 1751.710 202.645 1751.880 ;
        RECT 201.995 1751.620 202.645 1751.710 ;
        RECT 201.995 1751.420 202.165 1751.620 ;
        RECT 202.815 1751.450 202.985 1752.120 ;
        RECT 202.335 1751.280 202.985 1751.450 ;
        RECT 201.995 1751.020 202.165 1751.250 ;
      LAYER li1 ;
        RECT 203.155 1751.245 203.355 1752.345 ;
      LAYER li1 ;
        RECT 203.525 1752.040 204.545 1752.370 ;
        RECT 204.715 1752.340 204.885 1752.420 ;
      LAYER li1 ;
        RECT 205.905 1752.335 206.075 1752.920 ;
      LAYER li1 ;
        RECT 206.275 1752.580 206.445 1755.030 ;
        RECT 206.955 1754.940 207.435 1755.270 ;
      LAYER li1 ;
        RECT 206.615 1754.600 207.265 1754.770 ;
        RECT 206.615 1753.930 206.785 1754.600 ;
      LAYER li1 ;
        RECT 206.955 1754.100 207.435 1754.430 ;
      LAYER li1 ;
        RECT 206.615 1753.760 207.265 1753.930 ;
        RECT 206.615 1753.090 206.785 1753.760 ;
      LAYER li1 ;
        RECT 206.955 1753.260 207.435 1753.590 ;
      LAYER li1 ;
        RECT 206.615 1752.920 207.265 1753.090 ;
        RECT 206.615 1752.335 206.785 1752.920 ;
      LAYER li1 ;
        RECT 206.955 1752.420 207.435 1752.750 ;
      LAYER li1 ;
        RECT 205.855 1752.250 206.785 1752.335 ;
      LAYER li1 ;
        RECT 203.525 1751.530 203.695 1752.040 ;
        RECT 204.715 1751.910 204.885 1752.170 ;
      LAYER li1 ;
        RECT 205.055 1752.080 207.265 1752.250 ;
      LAYER li1 ;
        RECT 204.715 1751.880 206.035 1751.910 ;
        RECT 203.915 1751.710 204.715 1751.870 ;
        RECT 204.885 1751.710 206.035 1751.880 ;
        RECT 203.915 1751.700 206.035 1751.710 ;
        RECT 204.715 1751.580 206.035 1751.700 ;
        RECT 206.635 1751.580 207.435 1751.910 ;
        RECT 203.525 1751.200 204.545 1751.530 ;
        RECT 204.715 1751.420 204.885 1751.580 ;
        RECT 204.715 1751.020 204.885 1751.250 ;
        RECT 207.435 1751.020 207.605 1751.105 ;
        RECT 210.155 1751.020 210.325 1751.105 ;
        RECT 201.995 1750.960 202.890 1751.020 ;
        RECT 202.165 1750.790 202.890 1750.960 ;
        RECT 201.995 1750.730 202.890 1750.790 ;
        RECT 203.550 1750.960 206.050 1751.020 ;
        RECT 203.550 1750.790 204.715 1750.960 ;
        RECT 204.885 1750.790 206.050 1750.960 ;
        RECT 203.550 1750.730 206.050 1750.790 ;
        RECT 201.995 1750.500 202.165 1750.730 ;
        RECT 204.715 1750.500 204.885 1750.730 ;
        RECT 201.995 1750.170 202.165 1750.330 ;
        RECT 204.715 1750.170 204.885 1750.330 ;
        RECT 205.055 1750.220 206.075 1750.550 ;
        RECT 201.995 1750.040 202.965 1750.170 ;
        RECT 202.165 1749.870 202.965 1750.040 ;
        RECT 201.995 1749.840 202.965 1749.870 ;
        RECT 203.565 1750.050 204.885 1750.170 ;
        RECT 203.565 1750.040 205.685 1750.050 ;
        RECT 203.565 1749.870 204.715 1750.040 ;
        RECT 204.885 1749.880 205.685 1750.040 ;
        RECT 203.565 1749.840 204.885 1749.870 ;
        RECT 201.995 1749.580 202.165 1749.840 ;
      LAYER li1 ;
        RECT 202.335 1749.500 204.545 1749.670 ;
      LAYER li1 ;
        RECT 204.715 1749.580 204.885 1749.840 ;
        RECT 205.905 1749.710 206.075 1750.220 ;
      LAYER li1 ;
        RECT 202.815 1749.415 203.695 1749.500 ;
      LAYER li1 ;
        RECT 201.995 1749.330 202.165 1749.410 ;
        RECT 201.995 1749.120 202.645 1749.330 ;
        RECT 202.165 1749.000 202.645 1749.120 ;
        RECT 201.995 1748.660 202.165 1748.950 ;
      LAYER li1 ;
        RECT 202.815 1748.830 202.985 1749.415 ;
        RECT 202.335 1748.660 202.985 1748.830 ;
      LAYER li1 ;
        RECT 201.995 1748.200 202.645 1748.490 ;
        RECT 202.165 1748.160 202.645 1748.200 ;
        RECT 201.995 1747.740 202.165 1748.030 ;
      LAYER li1 ;
        RECT 202.815 1747.990 202.985 1748.660 ;
        RECT 202.335 1747.820 202.985 1747.990 ;
      LAYER li1 ;
        RECT 202.165 1747.570 202.645 1747.650 ;
        RECT 201.995 1747.320 202.645 1747.570 ;
        RECT 201.995 1747.280 202.165 1747.320 ;
      LAYER li1 ;
        RECT 202.815 1747.150 202.985 1747.820 ;
      LAYER li1 ;
        RECT 201.995 1746.820 202.165 1747.110 ;
      LAYER li1 ;
        RECT 202.335 1746.980 202.985 1747.150 ;
      LAYER li1 ;
        RECT 202.165 1746.650 202.645 1746.810 ;
        RECT 203.155 1746.720 203.325 1749.170 ;
      LAYER li1 ;
        RECT 203.525 1748.830 203.695 1749.415 ;
      LAYER li1 ;
        RECT 204.715 1749.330 204.885 1749.410 ;
        RECT 205.055 1749.380 206.075 1749.710 ;
      LAYER li1 ;
        RECT 206.245 1749.405 206.445 1750.995 ;
      LAYER li1 ;
        RECT 206.710 1750.960 208.330 1751.020 ;
        RECT 206.710 1750.790 207.435 1750.960 ;
        RECT 207.605 1750.790 208.330 1750.960 ;
        RECT 206.710 1750.730 208.330 1750.790 ;
        RECT 208.990 1750.960 210.325 1751.020 ;
        RECT 208.990 1750.790 210.155 1750.960 ;
        RECT 208.990 1750.730 210.325 1750.790 ;
        RECT 207.435 1750.500 207.605 1750.730 ;
        RECT 206.615 1750.300 207.265 1750.470 ;
        RECT 206.615 1749.630 206.785 1750.300 ;
        RECT 207.435 1750.130 207.605 1750.330 ;
        RECT 207.775 1750.300 208.425 1750.470 ;
        RECT 206.955 1750.040 208.085 1750.130 ;
        RECT 206.955 1749.870 207.435 1750.040 ;
        RECT 207.605 1749.870 208.085 1750.040 ;
        RECT 206.955 1749.800 208.085 1749.870 ;
        RECT 206.615 1749.460 207.260 1749.630 ;
        RECT 207.435 1749.580 207.605 1749.800 ;
        RECT 208.255 1749.630 208.425 1750.300 ;
        RECT 207.780 1749.460 208.425 1749.630 ;
        RECT 203.915 1749.210 204.885 1749.330 ;
        RECT 205.905 1749.225 206.075 1749.380 ;
        RECT 206.615 1749.225 206.785 1749.460 ;
        RECT 207.435 1749.290 207.605 1749.410 ;
        RECT 203.915 1749.120 205.685 1749.210 ;
        RECT 203.915 1749.000 204.715 1749.120 ;
        RECT 204.885 1749.040 205.685 1749.120 ;
        RECT 205.905 1749.050 206.785 1749.225 ;
        RECT 206.955 1749.120 208.085 1749.290 ;
      LAYER li1 ;
        RECT 203.525 1748.660 204.545 1748.830 ;
      LAYER li1 ;
        RECT 204.715 1748.660 204.885 1748.950 ;
      LAYER li1 ;
        RECT 203.525 1747.990 203.695 1748.660 ;
        RECT 205.055 1748.620 206.075 1748.790 ;
      LAYER li1 ;
        RECT 203.915 1748.450 204.885 1748.490 ;
        RECT 203.915 1748.200 205.685 1748.450 ;
        RECT 203.915 1748.160 204.715 1748.200 ;
        RECT 204.885 1748.120 205.685 1748.200 ;
      LAYER li1 ;
        RECT 203.525 1747.820 204.545 1747.990 ;
        RECT 203.525 1747.150 203.695 1747.820 ;
      LAYER li1 ;
        RECT 204.715 1747.740 204.885 1748.030 ;
      LAYER li1 ;
        RECT 205.905 1747.950 206.075 1748.620 ;
        RECT 205.055 1747.780 206.075 1747.950 ;
      LAYER li1 ;
        RECT 203.915 1747.570 204.715 1747.650 ;
        RECT 204.885 1747.570 205.685 1747.610 ;
        RECT 203.915 1747.320 205.685 1747.570 ;
        RECT 204.715 1747.280 205.685 1747.320 ;
      LAYER li1 ;
        RECT 203.525 1746.980 204.545 1747.150 ;
        RECT 205.905 1747.110 206.075 1747.780 ;
      LAYER li1 ;
        RECT 204.715 1746.820 204.885 1747.110 ;
      LAYER li1 ;
        RECT 205.055 1746.940 206.075 1747.110 ;
      LAYER li1 ;
        RECT 201.995 1746.480 202.645 1746.650 ;
        RECT 202.815 1746.545 203.695 1746.720 ;
        RECT 203.915 1746.650 204.715 1746.730 ;
        RECT 204.885 1746.650 205.685 1746.770 ;
        RECT 203.915 1746.560 205.685 1746.650 ;
        RECT 201.995 1746.360 202.165 1746.480 ;
        RECT 202.815 1746.310 202.985 1746.545 ;
        RECT 203.525 1746.390 203.695 1746.545 ;
        RECT 204.715 1746.440 205.685 1746.560 ;
        RECT 201.995 1745.970 202.165 1746.190 ;
        RECT 202.340 1746.140 202.985 1746.310 ;
        RECT 201.995 1745.900 202.645 1745.970 ;
        RECT 202.165 1745.730 202.645 1745.900 ;
        RECT 201.995 1745.640 202.645 1745.730 ;
        RECT 201.995 1745.440 202.165 1745.640 ;
        RECT 202.815 1745.470 202.985 1746.140 ;
        RECT 202.335 1745.300 202.985 1745.470 ;
        RECT 201.995 1745.040 202.165 1745.270 ;
      LAYER li1 ;
        RECT 203.155 1745.265 203.355 1746.365 ;
      LAYER li1 ;
        RECT 203.525 1746.060 204.545 1746.390 ;
        RECT 204.715 1746.360 204.885 1746.440 ;
      LAYER li1 ;
        RECT 205.905 1746.355 206.075 1746.940 ;
      LAYER li1 ;
        RECT 206.275 1746.600 206.445 1749.050 ;
        RECT 206.955 1748.960 207.435 1749.120 ;
        RECT 207.605 1748.960 208.085 1749.120 ;
        RECT 208.255 1749.225 208.425 1749.460 ;
      LAYER li1 ;
        RECT 208.595 1749.405 208.795 1750.505 ;
      LAYER li1 ;
        RECT 208.965 1750.220 209.985 1750.550 ;
        RECT 210.155 1750.500 210.325 1750.730 ;
        RECT 208.965 1749.710 209.135 1750.220 ;
        RECT 210.155 1750.050 210.325 1750.330 ;
        RECT 209.355 1750.040 210.325 1750.050 ;
        RECT 209.355 1749.880 210.155 1750.040 ;
        RECT 208.965 1749.380 209.985 1749.710 ;
        RECT 210.155 1749.580 210.325 1749.870 ;
        RECT 208.965 1749.225 209.135 1749.380 ;
        RECT 208.255 1749.050 209.135 1749.225 ;
        RECT 210.155 1749.210 210.325 1749.410 ;
        RECT 209.355 1749.120 210.325 1749.210 ;
      LAYER li1 ;
        RECT 206.615 1748.620 207.265 1748.790 ;
      LAYER li1 ;
        RECT 207.435 1748.660 207.605 1748.950 ;
      LAYER li1 ;
        RECT 207.775 1748.620 208.425 1748.790 ;
        RECT 206.615 1747.950 206.785 1748.620 ;
      LAYER li1 ;
        RECT 207.435 1748.450 207.605 1748.490 ;
        RECT 206.955 1748.200 208.085 1748.450 ;
        RECT 206.955 1748.120 207.435 1748.200 ;
        RECT 207.605 1748.120 208.085 1748.200 ;
      LAYER li1 ;
        RECT 206.615 1747.780 207.265 1747.950 ;
        RECT 206.615 1747.110 206.785 1747.780 ;
      LAYER li1 ;
        RECT 207.435 1747.740 207.605 1748.030 ;
      LAYER li1 ;
        RECT 208.255 1747.950 208.425 1748.620 ;
        RECT 207.775 1747.780 208.425 1747.950 ;
      LAYER li1 ;
        RECT 206.955 1747.570 207.435 1747.610 ;
        RECT 207.605 1747.570 208.085 1747.610 ;
        RECT 206.955 1747.280 208.085 1747.570 ;
      LAYER li1 ;
        RECT 208.255 1747.110 208.425 1747.780 ;
        RECT 206.615 1746.940 207.265 1747.110 ;
        RECT 206.615 1746.355 206.785 1746.940 ;
      LAYER li1 ;
        RECT 207.435 1746.820 207.605 1747.110 ;
      LAYER li1 ;
        RECT 207.775 1746.940 208.425 1747.110 ;
      LAYER li1 ;
        RECT 206.955 1746.650 207.435 1746.770 ;
        RECT 207.605 1746.650 208.085 1746.770 ;
        RECT 206.955 1746.440 208.085 1746.650 ;
        RECT 207.435 1746.360 207.605 1746.440 ;
      LAYER li1 ;
        RECT 205.905 1746.270 206.785 1746.355 ;
        RECT 208.255 1746.355 208.425 1746.940 ;
      LAYER li1 ;
        RECT 208.595 1746.600 208.765 1749.050 ;
        RECT 209.355 1749.040 210.155 1749.120 ;
      LAYER li1 ;
        RECT 208.965 1748.620 209.985 1748.790 ;
      LAYER li1 ;
        RECT 210.155 1748.660 210.325 1748.950 ;
      LAYER li1 ;
        RECT 208.965 1747.950 209.135 1748.620 ;
      LAYER li1 ;
        RECT 210.155 1748.450 210.325 1748.490 ;
        RECT 209.355 1748.200 210.325 1748.450 ;
        RECT 209.355 1748.120 210.155 1748.200 ;
      LAYER li1 ;
        RECT 208.965 1747.780 209.985 1747.950 ;
        RECT 208.965 1747.110 209.135 1747.780 ;
      LAYER li1 ;
        RECT 210.155 1747.740 210.325 1748.030 ;
        RECT 209.355 1747.570 210.155 1747.610 ;
        RECT 209.355 1747.280 210.325 1747.570 ;
      LAYER li1 ;
        RECT 208.965 1746.940 209.985 1747.110 ;
        RECT 208.965 1746.355 209.135 1746.940 ;
      LAYER li1 ;
        RECT 210.155 1746.820 210.325 1747.110 ;
        RECT 209.355 1746.650 210.155 1746.770 ;
        RECT 209.355 1746.440 210.325 1746.650 ;
        RECT 210.155 1746.360 210.325 1746.440 ;
      LAYER li1 ;
        RECT 208.255 1746.270 209.135 1746.355 ;
      LAYER li1 ;
        RECT 203.525 1745.550 203.695 1746.060 ;
        RECT 204.715 1745.930 204.885 1746.190 ;
      LAYER li1 ;
        RECT 205.055 1746.100 207.265 1746.270 ;
      LAYER li1 ;
        RECT 207.435 1745.930 207.605 1746.190 ;
      LAYER li1 ;
        RECT 207.775 1746.100 209.985 1746.270 ;
      LAYER li1 ;
        RECT 210.155 1745.930 210.325 1746.190 ;
        RECT 204.715 1745.900 206.035 1745.930 ;
        RECT 203.915 1745.730 204.715 1745.890 ;
        RECT 204.885 1745.730 206.035 1745.900 ;
        RECT 203.915 1745.720 206.035 1745.730 ;
        RECT 204.715 1745.600 206.035 1745.720 ;
        RECT 206.635 1745.900 208.405 1745.930 ;
        RECT 206.635 1745.730 207.435 1745.900 ;
        RECT 207.605 1745.730 208.405 1745.900 ;
        RECT 206.635 1745.600 208.405 1745.730 ;
        RECT 209.005 1745.900 210.325 1745.930 ;
        RECT 209.005 1745.730 210.155 1745.900 ;
        RECT 209.005 1745.600 210.325 1745.730 ;
        RECT 203.525 1745.220 204.545 1745.550 ;
        RECT 204.715 1745.440 204.885 1745.600 ;
        RECT 207.435 1745.440 207.605 1745.600 ;
        RECT 210.155 1745.440 210.325 1745.600 ;
        RECT 204.715 1745.040 204.885 1745.270 ;
        RECT 207.435 1745.040 207.605 1745.270 ;
        RECT 210.155 1745.040 210.325 1745.270 ;
        RECT 201.995 1744.980 202.890 1745.040 ;
        RECT 202.165 1744.810 202.890 1744.980 ;
        RECT 201.995 1744.750 202.890 1744.810 ;
        RECT 203.550 1744.980 206.050 1745.040 ;
        RECT 203.550 1744.810 204.715 1744.980 ;
        RECT 204.885 1744.810 206.050 1744.980 ;
        RECT 203.550 1744.750 206.050 1744.810 ;
        RECT 201.995 1744.520 202.165 1744.750 ;
        RECT 204.715 1744.520 204.885 1744.750 ;
        RECT 201.995 1744.190 202.165 1744.350 ;
        RECT 204.715 1744.190 204.885 1744.350 ;
        RECT 205.055 1744.240 206.075 1744.570 ;
        RECT 201.995 1744.060 202.965 1744.190 ;
        RECT 202.165 1743.890 202.965 1744.060 ;
        RECT 201.995 1743.860 202.965 1743.890 ;
        RECT 203.565 1744.070 204.885 1744.190 ;
        RECT 203.565 1744.060 205.685 1744.070 ;
        RECT 203.565 1743.890 204.715 1744.060 ;
        RECT 204.885 1743.900 205.685 1744.060 ;
        RECT 203.565 1743.860 204.885 1743.890 ;
        RECT 201.995 1743.600 202.165 1743.860 ;
      LAYER li1 ;
        RECT 202.335 1743.520 204.545 1743.690 ;
      LAYER li1 ;
        RECT 204.715 1743.600 204.885 1743.860 ;
        RECT 205.905 1743.730 206.075 1744.240 ;
      LAYER li1 ;
        RECT 202.815 1743.435 203.695 1743.520 ;
      LAYER li1 ;
        RECT 201.995 1743.350 202.165 1743.430 ;
        RECT 201.995 1743.140 202.645 1743.350 ;
        RECT 202.165 1743.020 202.645 1743.140 ;
        RECT 201.995 1742.680 202.165 1742.970 ;
      LAYER li1 ;
        RECT 202.815 1742.850 202.985 1743.435 ;
        RECT 202.335 1742.680 202.985 1742.850 ;
      LAYER li1 ;
        RECT 201.995 1742.220 202.645 1742.510 ;
        RECT 202.165 1742.180 202.645 1742.220 ;
        RECT 201.995 1741.760 202.165 1742.050 ;
      LAYER li1 ;
        RECT 202.815 1742.010 202.985 1742.680 ;
        RECT 202.335 1741.840 202.985 1742.010 ;
      LAYER li1 ;
        RECT 202.165 1741.590 202.645 1741.670 ;
        RECT 201.995 1741.340 202.645 1741.590 ;
        RECT 201.995 1741.300 202.165 1741.340 ;
      LAYER li1 ;
        RECT 202.815 1741.170 202.985 1741.840 ;
      LAYER li1 ;
        RECT 201.995 1740.840 202.165 1741.130 ;
      LAYER li1 ;
        RECT 202.335 1741.000 202.985 1741.170 ;
      LAYER li1 ;
        RECT 202.165 1740.670 202.645 1740.830 ;
        RECT 203.155 1740.740 203.325 1743.190 ;
      LAYER li1 ;
        RECT 203.525 1742.850 203.695 1743.435 ;
      LAYER li1 ;
        RECT 204.715 1743.350 204.885 1743.430 ;
        RECT 205.055 1743.400 206.075 1743.730 ;
      LAYER li1 ;
        RECT 206.245 1743.425 206.445 1745.015 ;
      LAYER li1 ;
        RECT 206.710 1744.980 208.330 1745.040 ;
        RECT 206.710 1744.810 207.435 1744.980 ;
        RECT 207.605 1744.810 208.330 1744.980 ;
        RECT 206.710 1744.750 208.330 1744.810 ;
        RECT 208.990 1744.980 210.325 1745.040 ;
        RECT 208.990 1744.810 210.155 1744.980 ;
        RECT 208.990 1744.750 210.325 1744.810 ;
        RECT 207.435 1744.665 207.605 1744.750 ;
        RECT 210.155 1744.665 210.325 1744.750 ;
        RECT 206.615 1744.320 207.265 1744.490 ;
        RECT 206.615 1743.650 206.785 1744.320 ;
        RECT 206.955 1743.820 207.435 1744.150 ;
        RECT 206.615 1743.480 207.260 1743.650 ;
        RECT 203.915 1743.230 204.885 1743.350 ;
        RECT 205.905 1743.245 206.075 1743.400 ;
        RECT 206.615 1743.245 206.785 1743.480 ;
        RECT 203.915 1743.140 205.685 1743.230 ;
        RECT 203.915 1743.020 204.715 1743.140 ;
        RECT 204.885 1743.060 205.685 1743.140 ;
        RECT 205.905 1743.070 206.785 1743.245 ;
      LAYER li1 ;
        RECT 203.525 1742.680 204.545 1742.850 ;
      LAYER li1 ;
        RECT 204.715 1742.680 204.885 1742.970 ;
      LAYER li1 ;
        RECT 203.525 1742.010 203.695 1742.680 ;
        RECT 205.055 1742.640 206.075 1742.810 ;
      LAYER li1 ;
        RECT 203.915 1742.470 204.885 1742.510 ;
        RECT 203.915 1742.220 205.685 1742.470 ;
        RECT 203.915 1742.180 204.715 1742.220 ;
        RECT 204.885 1742.140 205.685 1742.220 ;
      LAYER li1 ;
        RECT 203.525 1741.840 204.545 1742.010 ;
        RECT 203.525 1741.170 203.695 1741.840 ;
      LAYER li1 ;
        RECT 204.715 1741.760 204.885 1742.050 ;
      LAYER li1 ;
        RECT 205.905 1741.970 206.075 1742.640 ;
        RECT 205.055 1741.800 206.075 1741.970 ;
      LAYER li1 ;
        RECT 203.915 1741.590 204.715 1741.670 ;
        RECT 204.885 1741.590 205.685 1741.630 ;
        RECT 203.915 1741.340 205.685 1741.590 ;
        RECT 204.715 1741.300 205.685 1741.340 ;
      LAYER li1 ;
        RECT 203.525 1741.000 204.545 1741.170 ;
        RECT 205.905 1741.130 206.075 1741.800 ;
      LAYER li1 ;
        RECT 204.715 1740.840 204.885 1741.130 ;
      LAYER li1 ;
        RECT 205.055 1740.960 206.075 1741.130 ;
      LAYER li1 ;
        RECT 201.995 1740.500 202.645 1740.670 ;
        RECT 202.815 1740.565 203.695 1740.740 ;
        RECT 203.915 1740.670 204.715 1740.750 ;
        RECT 204.885 1740.670 205.685 1740.790 ;
        RECT 203.915 1740.580 205.685 1740.670 ;
        RECT 201.995 1740.380 202.165 1740.500 ;
        RECT 202.815 1740.330 202.985 1740.565 ;
        RECT 203.525 1740.410 203.695 1740.565 ;
        RECT 204.715 1740.460 205.685 1740.580 ;
        RECT 201.995 1739.990 202.165 1740.210 ;
        RECT 202.340 1740.160 202.985 1740.330 ;
        RECT 201.995 1739.920 202.645 1739.990 ;
        RECT 202.165 1739.750 202.645 1739.920 ;
        RECT 201.995 1739.660 202.645 1739.750 ;
        RECT 201.995 1739.460 202.165 1739.660 ;
        RECT 202.815 1739.490 202.985 1740.160 ;
        RECT 202.335 1739.320 202.985 1739.490 ;
        RECT 201.995 1739.060 202.165 1739.290 ;
      LAYER li1 ;
        RECT 203.155 1739.285 203.355 1740.385 ;
      LAYER li1 ;
        RECT 203.525 1740.080 204.545 1740.410 ;
        RECT 204.715 1740.380 204.885 1740.460 ;
      LAYER li1 ;
        RECT 205.905 1740.375 206.075 1740.960 ;
      LAYER li1 ;
        RECT 206.275 1740.620 206.445 1743.070 ;
        RECT 206.955 1742.980 207.435 1743.310 ;
      LAYER li1 ;
        RECT 206.615 1742.640 207.265 1742.810 ;
        RECT 206.615 1741.970 206.785 1742.640 ;
      LAYER li1 ;
        RECT 206.955 1742.140 207.435 1742.470 ;
      LAYER li1 ;
        RECT 206.615 1741.800 207.265 1741.970 ;
        RECT 206.615 1741.130 206.785 1741.800 ;
      LAYER li1 ;
        RECT 206.955 1741.300 207.435 1741.630 ;
      LAYER li1 ;
        RECT 206.615 1740.960 207.265 1741.130 ;
        RECT 206.615 1740.375 206.785 1740.960 ;
      LAYER li1 ;
        RECT 206.955 1740.460 207.435 1740.790 ;
      LAYER li1 ;
        RECT 205.905 1740.290 206.785 1740.375 ;
      LAYER li1 ;
        RECT 203.525 1739.570 203.695 1740.080 ;
        RECT 204.715 1739.950 204.885 1740.210 ;
      LAYER li1 ;
        RECT 205.055 1740.120 207.265 1740.290 ;
      LAYER li1 ;
        RECT 204.715 1739.920 206.035 1739.950 ;
        RECT 203.915 1739.750 204.715 1739.910 ;
        RECT 204.885 1739.750 206.035 1739.920 ;
        RECT 203.915 1739.740 206.035 1739.750 ;
        RECT 204.715 1739.620 206.035 1739.740 ;
        RECT 206.635 1739.620 207.435 1739.950 ;
        RECT 203.525 1739.240 204.545 1739.570 ;
        RECT 204.715 1739.460 204.885 1739.620 ;
        RECT 204.715 1739.060 204.885 1739.290 ;
        RECT 207.435 1739.060 207.605 1739.145 ;
        RECT 210.155 1739.060 210.325 1739.145 ;
        RECT 201.995 1739.000 202.890 1739.060 ;
        RECT 202.165 1738.830 202.890 1739.000 ;
        RECT 201.995 1738.770 202.890 1738.830 ;
        RECT 203.550 1739.000 206.050 1739.060 ;
        RECT 203.550 1738.830 204.715 1739.000 ;
        RECT 204.885 1738.830 206.050 1739.000 ;
        RECT 203.550 1738.770 206.050 1738.830 ;
        RECT 201.995 1738.540 202.165 1738.770 ;
        RECT 204.715 1738.540 204.885 1738.770 ;
        RECT 201.995 1738.210 202.165 1738.370 ;
        RECT 204.715 1738.210 204.885 1738.370 ;
        RECT 205.055 1738.260 206.075 1738.590 ;
        RECT 201.995 1738.080 202.965 1738.210 ;
        RECT 202.165 1737.910 202.965 1738.080 ;
        RECT 201.995 1737.880 202.965 1737.910 ;
        RECT 203.565 1738.090 204.885 1738.210 ;
        RECT 203.565 1738.080 205.685 1738.090 ;
        RECT 203.565 1737.910 204.715 1738.080 ;
        RECT 204.885 1737.920 205.685 1738.080 ;
        RECT 203.565 1737.880 204.885 1737.910 ;
        RECT 201.995 1737.620 202.165 1737.880 ;
      LAYER li1 ;
        RECT 202.335 1737.540 204.545 1737.710 ;
      LAYER li1 ;
        RECT 204.715 1737.620 204.885 1737.880 ;
        RECT 205.905 1737.750 206.075 1738.260 ;
      LAYER li1 ;
        RECT 202.815 1737.455 203.695 1737.540 ;
      LAYER li1 ;
        RECT 201.995 1737.370 202.165 1737.450 ;
        RECT 201.995 1737.160 202.645 1737.370 ;
        RECT 202.165 1737.040 202.645 1737.160 ;
        RECT 201.995 1736.700 202.165 1736.990 ;
      LAYER li1 ;
        RECT 202.815 1736.870 202.985 1737.455 ;
        RECT 202.335 1736.700 202.985 1736.870 ;
      LAYER li1 ;
        RECT 201.995 1736.240 202.645 1736.530 ;
        RECT 202.165 1736.200 202.645 1736.240 ;
        RECT 201.995 1735.780 202.165 1736.070 ;
      LAYER li1 ;
        RECT 202.815 1736.030 202.985 1736.700 ;
        RECT 202.335 1735.860 202.985 1736.030 ;
      LAYER li1 ;
        RECT 202.165 1735.610 202.645 1735.690 ;
        RECT 201.995 1735.360 202.645 1735.610 ;
        RECT 201.995 1735.320 202.165 1735.360 ;
      LAYER li1 ;
        RECT 202.815 1735.190 202.985 1735.860 ;
      LAYER li1 ;
        RECT 201.995 1734.860 202.165 1735.150 ;
      LAYER li1 ;
        RECT 202.335 1735.020 202.985 1735.190 ;
      LAYER li1 ;
        RECT 202.165 1734.690 202.645 1734.850 ;
        RECT 203.155 1734.760 203.325 1737.210 ;
      LAYER li1 ;
        RECT 203.525 1736.870 203.695 1737.455 ;
      LAYER li1 ;
        RECT 204.715 1737.370 204.885 1737.450 ;
        RECT 205.055 1737.420 206.075 1737.750 ;
      LAYER li1 ;
        RECT 206.245 1737.445 206.445 1739.035 ;
      LAYER li1 ;
        RECT 206.710 1739.000 208.330 1739.060 ;
        RECT 206.710 1738.830 207.435 1739.000 ;
        RECT 207.605 1738.830 208.330 1739.000 ;
        RECT 206.710 1738.770 208.330 1738.830 ;
        RECT 208.990 1739.000 210.325 1739.060 ;
        RECT 208.990 1738.830 210.155 1739.000 ;
        RECT 208.990 1738.770 210.325 1738.830 ;
        RECT 207.435 1738.685 207.605 1738.770 ;
        RECT 210.155 1738.685 210.325 1738.770 ;
        RECT 206.615 1738.340 207.265 1738.510 ;
        RECT 206.615 1737.670 206.785 1738.340 ;
        RECT 206.955 1737.840 207.435 1738.170 ;
        RECT 206.615 1737.500 207.260 1737.670 ;
        RECT 203.915 1737.250 204.885 1737.370 ;
        RECT 205.905 1737.265 206.075 1737.420 ;
        RECT 206.615 1737.265 206.785 1737.500 ;
        RECT 203.915 1737.160 205.685 1737.250 ;
        RECT 203.915 1737.040 204.715 1737.160 ;
        RECT 204.885 1737.080 205.685 1737.160 ;
        RECT 205.905 1737.090 206.785 1737.265 ;
      LAYER li1 ;
        RECT 203.525 1736.700 204.545 1736.870 ;
      LAYER li1 ;
        RECT 204.715 1736.700 204.885 1736.990 ;
      LAYER li1 ;
        RECT 203.525 1736.030 203.695 1736.700 ;
        RECT 205.055 1736.660 206.075 1736.830 ;
      LAYER li1 ;
        RECT 203.915 1736.490 204.885 1736.530 ;
        RECT 203.915 1736.240 205.685 1736.490 ;
        RECT 203.915 1736.200 204.715 1736.240 ;
        RECT 204.885 1736.160 205.685 1736.240 ;
      LAYER li1 ;
        RECT 203.525 1735.860 204.545 1736.030 ;
        RECT 203.525 1735.190 203.695 1735.860 ;
      LAYER li1 ;
        RECT 204.715 1735.780 204.885 1736.070 ;
      LAYER li1 ;
        RECT 205.905 1735.990 206.075 1736.660 ;
        RECT 205.055 1735.820 206.075 1735.990 ;
      LAYER li1 ;
        RECT 203.915 1735.610 204.715 1735.690 ;
        RECT 204.885 1735.610 205.685 1735.650 ;
        RECT 203.915 1735.360 205.685 1735.610 ;
        RECT 204.715 1735.320 205.685 1735.360 ;
      LAYER li1 ;
        RECT 203.525 1735.020 204.545 1735.190 ;
        RECT 205.905 1735.150 206.075 1735.820 ;
      LAYER li1 ;
        RECT 204.715 1734.860 204.885 1735.150 ;
      LAYER li1 ;
        RECT 205.055 1734.980 206.075 1735.150 ;
      LAYER li1 ;
        RECT 201.995 1734.520 202.645 1734.690 ;
        RECT 202.815 1734.585 203.695 1734.760 ;
        RECT 203.915 1734.690 204.715 1734.770 ;
        RECT 204.885 1734.690 205.685 1734.810 ;
        RECT 203.915 1734.600 205.685 1734.690 ;
        RECT 201.995 1734.400 202.165 1734.520 ;
        RECT 202.815 1734.350 202.985 1734.585 ;
        RECT 203.525 1734.430 203.695 1734.585 ;
        RECT 204.715 1734.480 205.685 1734.600 ;
        RECT 201.995 1734.010 202.165 1734.230 ;
        RECT 202.340 1734.180 202.985 1734.350 ;
        RECT 201.995 1733.940 202.645 1734.010 ;
        RECT 202.165 1733.770 202.645 1733.940 ;
        RECT 201.995 1733.680 202.645 1733.770 ;
        RECT 201.995 1733.480 202.165 1733.680 ;
        RECT 202.815 1733.510 202.985 1734.180 ;
        RECT 202.335 1733.340 202.985 1733.510 ;
        RECT 201.995 1733.080 202.165 1733.310 ;
      LAYER li1 ;
        RECT 203.155 1733.305 203.355 1734.405 ;
      LAYER li1 ;
        RECT 203.525 1734.100 204.545 1734.430 ;
        RECT 204.715 1734.400 204.885 1734.480 ;
      LAYER li1 ;
        RECT 205.905 1734.395 206.075 1734.980 ;
      LAYER li1 ;
        RECT 206.275 1734.640 206.445 1737.090 ;
        RECT 206.955 1737.000 207.435 1737.330 ;
      LAYER li1 ;
        RECT 206.615 1736.660 207.265 1736.830 ;
        RECT 206.615 1735.990 206.785 1736.660 ;
      LAYER li1 ;
        RECT 206.955 1736.160 207.435 1736.490 ;
      LAYER li1 ;
        RECT 206.615 1735.820 207.265 1735.990 ;
        RECT 206.615 1735.150 206.785 1735.820 ;
      LAYER li1 ;
        RECT 206.955 1735.320 207.435 1735.650 ;
      LAYER li1 ;
        RECT 206.615 1734.980 207.265 1735.150 ;
        RECT 206.615 1734.395 206.785 1734.980 ;
      LAYER li1 ;
        RECT 206.955 1734.480 207.435 1734.810 ;
      LAYER li1 ;
        RECT 205.905 1734.310 206.785 1734.395 ;
      LAYER li1 ;
        RECT 203.525 1733.590 203.695 1734.100 ;
        RECT 204.715 1733.970 204.885 1734.230 ;
      LAYER li1 ;
        RECT 205.055 1734.140 207.265 1734.310 ;
      LAYER li1 ;
        RECT 204.715 1733.940 206.035 1733.970 ;
        RECT 203.915 1733.770 204.715 1733.930 ;
        RECT 204.885 1733.770 206.035 1733.940 ;
        RECT 203.915 1733.760 206.035 1733.770 ;
        RECT 204.715 1733.640 206.035 1733.760 ;
        RECT 206.635 1733.640 207.435 1733.970 ;
        RECT 203.525 1733.260 204.545 1733.590 ;
        RECT 204.715 1733.480 204.885 1733.640 ;
        RECT 204.715 1733.080 204.885 1733.310 ;
        RECT 207.435 1733.080 207.605 1733.165 ;
        RECT 210.155 1733.080 210.325 1733.165 ;
        RECT 201.995 1733.020 202.890 1733.080 ;
        RECT 202.165 1732.850 202.890 1733.020 ;
        RECT 201.995 1732.790 202.890 1732.850 ;
        RECT 203.550 1733.020 206.050 1733.080 ;
        RECT 203.550 1732.850 204.715 1733.020 ;
        RECT 204.885 1732.850 206.050 1733.020 ;
        RECT 203.550 1732.790 206.050 1732.850 ;
        RECT 201.995 1732.560 202.165 1732.790 ;
        RECT 204.715 1732.560 204.885 1732.790 ;
        RECT 201.995 1732.230 202.165 1732.390 ;
        RECT 204.715 1732.230 204.885 1732.390 ;
        RECT 205.055 1732.280 206.075 1732.610 ;
        RECT 201.995 1732.100 202.965 1732.230 ;
        RECT 202.165 1731.930 202.965 1732.100 ;
        RECT 201.995 1731.900 202.965 1731.930 ;
        RECT 203.565 1732.110 204.885 1732.230 ;
        RECT 203.565 1732.100 205.685 1732.110 ;
        RECT 203.565 1731.930 204.715 1732.100 ;
        RECT 204.885 1731.940 205.685 1732.100 ;
        RECT 203.565 1731.900 204.885 1731.930 ;
        RECT 201.995 1731.640 202.165 1731.900 ;
      LAYER li1 ;
        RECT 202.335 1731.560 204.545 1731.730 ;
      LAYER li1 ;
        RECT 204.715 1731.640 204.885 1731.900 ;
        RECT 205.905 1731.770 206.075 1732.280 ;
      LAYER li1 ;
        RECT 202.815 1731.475 203.695 1731.560 ;
      LAYER li1 ;
        RECT 201.995 1731.390 202.165 1731.470 ;
        RECT 201.995 1731.180 202.645 1731.390 ;
        RECT 202.165 1731.060 202.645 1731.180 ;
        RECT 201.995 1730.720 202.165 1731.010 ;
      LAYER li1 ;
        RECT 202.815 1730.890 202.985 1731.475 ;
        RECT 202.335 1730.720 202.985 1730.890 ;
      LAYER li1 ;
        RECT 201.995 1730.260 202.645 1730.550 ;
        RECT 202.165 1730.220 202.645 1730.260 ;
        RECT 201.995 1729.800 202.165 1730.090 ;
      LAYER li1 ;
        RECT 202.815 1730.050 202.985 1730.720 ;
        RECT 202.335 1729.880 202.985 1730.050 ;
      LAYER li1 ;
        RECT 202.165 1729.630 202.645 1729.710 ;
        RECT 201.995 1729.380 202.645 1729.630 ;
        RECT 201.995 1729.340 202.165 1729.380 ;
      LAYER li1 ;
        RECT 202.815 1729.210 202.985 1729.880 ;
      LAYER li1 ;
        RECT 201.995 1728.880 202.165 1729.170 ;
      LAYER li1 ;
        RECT 202.335 1729.040 202.985 1729.210 ;
      LAYER li1 ;
        RECT 202.165 1728.710 202.645 1728.870 ;
        RECT 203.155 1728.780 203.325 1731.230 ;
      LAYER li1 ;
        RECT 203.525 1730.890 203.695 1731.475 ;
      LAYER li1 ;
        RECT 204.715 1731.390 204.885 1731.470 ;
        RECT 205.055 1731.440 206.075 1731.770 ;
      LAYER li1 ;
        RECT 206.245 1731.465 206.445 1733.055 ;
      LAYER li1 ;
        RECT 206.710 1733.020 208.330 1733.080 ;
        RECT 206.710 1732.850 207.435 1733.020 ;
        RECT 207.605 1732.850 208.330 1733.020 ;
        RECT 206.710 1732.790 208.330 1732.850 ;
        RECT 208.990 1733.020 210.325 1733.080 ;
        RECT 208.990 1732.850 210.155 1733.020 ;
        RECT 208.990 1732.790 210.325 1732.850 ;
        RECT 207.435 1732.705 207.605 1732.790 ;
        RECT 210.155 1732.705 210.325 1732.790 ;
        RECT 206.615 1732.360 207.265 1732.530 ;
        RECT 206.615 1731.690 206.785 1732.360 ;
        RECT 206.955 1731.860 207.435 1732.190 ;
        RECT 206.615 1731.520 207.260 1731.690 ;
        RECT 203.915 1731.270 204.885 1731.390 ;
        RECT 205.905 1731.285 206.075 1731.440 ;
        RECT 206.615 1731.285 206.785 1731.520 ;
        RECT 203.915 1731.180 205.685 1731.270 ;
        RECT 203.915 1731.060 204.715 1731.180 ;
        RECT 204.885 1731.100 205.685 1731.180 ;
        RECT 205.905 1731.110 206.785 1731.285 ;
      LAYER li1 ;
        RECT 203.525 1730.720 204.545 1730.890 ;
      LAYER li1 ;
        RECT 204.715 1730.720 204.885 1731.010 ;
      LAYER li1 ;
        RECT 203.525 1730.050 203.695 1730.720 ;
        RECT 205.055 1730.680 206.075 1730.850 ;
      LAYER li1 ;
        RECT 203.915 1730.510 204.885 1730.550 ;
        RECT 203.915 1730.260 205.685 1730.510 ;
        RECT 203.915 1730.220 204.715 1730.260 ;
        RECT 204.885 1730.180 205.685 1730.260 ;
      LAYER li1 ;
        RECT 203.525 1729.880 204.545 1730.050 ;
        RECT 203.525 1729.210 203.695 1729.880 ;
      LAYER li1 ;
        RECT 204.715 1729.800 204.885 1730.090 ;
      LAYER li1 ;
        RECT 205.905 1730.010 206.075 1730.680 ;
        RECT 205.055 1729.840 206.075 1730.010 ;
      LAYER li1 ;
        RECT 203.915 1729.630 204.715 1729.710 ;
        RECT 204.885 1729.630 205.685 1729.670 ;
        RECT 203.915 1729.380 205.685 1729.630 ;
        RECT 204.715 1729.340 205.685 1729.380 ;
      LAYER li1 ;
        RECT 203.525 1729.040 204.545 1729.210 ;
        RECT 205.905 1729.170 206.075 1729.840 ;
      LAYER li1 ;
        RECT 204.715 1728.880 204.885 1729.170 ;
      LAYER li1 ;
        RECT 205.055 1729.000 206.075 1729.170 ;
      LAYER li1 ;
        RECT 201.995 1728.540 202.645 1728.710 ;
        RECT 202.815 1728.605 203.695 1728.780 ;
        RECT 203.915 1728.710 204.715 1728.790 ;
        RECT 204.885 1728.710 205.685 1728.830 ;
        RECT 203.915 1728.620 205.685 1728.710 ;
        RECT 201.995 1728.420 202.165 1728.540 ;
        RECT 202.815 1728.370 202.985 1728.605 ;
        RECT 203.525 1728.450 203.695 1728.605 ;
        RECT 204.715 1728.500 205.685 1728.620 ;
        RECT 201.995 1728.030 202.165 1728.250 ;
        RECT 202.340 1728.200 202.985 1728.370 ;
        RECT 201.995 1727.960 202.645 1728.030 ;
        RECT 202.165 1727.790 202.645 1727.960 ;
        RECT 201.995 1727.700 202.645 1727.790 ;
        RECT 201.995 1727.500 202.165 1727.700 ;
        RECT 202.815 1727.530 202.985 1728.200 ;
        RECT 202.335 1727.360 202.985 1727.530 ;
        RECT 201.995 1727.100 202.165 1727.330 ;
      LAYER li1 ;
        RECT 203.155 1727.325 203.355 1728.425 ;
      LAYER li1 ;
        RECT 203.525 1728.120 204.545 1728.450 ;
        RECT 204.715 1728.420 204.885 1728.500 ;
      LAYER li1 ;
        RECT 205.905 1728.415 206.075 1729.000 ;
      LAYER li1 ;
        RECT 206.275 1728.660 206.445 1731.110 ;
        RECT 206.955 1731.020 207.435 1731.350 ;
      LAYER li1 ;
        RECT 206.615 1730.680 207.265 1730.850 ;
        RECT 206.615 1730.010 206.785 1730.680 ;
      LAYER li1 ;
        RECT 206.955 1730.180 207.435 1730.510 ;
      LAYER li1 ;
        RECT 206.615 1729.840 207.265 1730.010 ;
        RECT 206.615 1729.170 206.785 1729.840 ;
      LAYER li1 ;
        RECT 206.955 1729.340 207.435 1729.670 ;
      LAYER li1 ;
        RECT 206.615 1729.000 207.265 1729.170 ;
        RECT 206.615 1728.415 206.785 1729.000 ;
      LAYER li1 ;
        RECT 206.955 1728.500 207.435 1728.830 ;
      LAYER li1 ;
        RECT 205.905 1728.330 206.785 1728.415 ;
      LAYER li1 ;
        RECT 203.525 1727.610 203.695 1728.120 ;
        RECT 204.715 1727.990 204.885 1728.250 ;
      LAYER li1 ;
        RECT 205.055 1728.160 207.265 1728.330 ;
      LAYER li1 ;
        RECT 204.715 1727.960 206.035 1727.990 ;
        RECT 203.915 1727.790 204.715 1727.950 ;
        RECT 204.885 1727.790 206.035 1727.960 ;
        RECT 203.915 1727.780 206.035 1727.790 ;
        RECT 204.715 1727.660 206.035 1727.780 ;
        RECT 206.635 1727.660 207.435 1727.990 ;
        RECT 203.525 1727.280 204.545 1727.610 ;
        RECT 204.715 1727.500 204.885 1727.660 ;
        RECT 204.715 1727.100 204.885 1727.330 ;
        RECT 207.435 1727.100 207.605 1727.185 ;
        RECT 210.155 1727.100 210.325 1727.185 ;
        RECT 201.995 1727.040 202.890 1727.100 ;
        RECT 202.165 1726.870 202.890 1727.040 ;
        RECT 201.995 1726.810 202.890 1726.870 ;
        RECT 203.550 1727.040 206.050 1727.100 ;
        RECT 203.550 1726.870 204.715 1727.040 ;
        RECT 204.885 1726.870 206.050 1727.040 ;
        RECT 203.550 1726.810 206.050 1726.870 ;
        RECT 201.995 1726.580 202.165 1726.810 ;
        RECT 204.715 1726.580 204.885 1726.810 ;
        RECT 201.995 1726.250 202.165 1726.410 ;
        RECT 204.715 1726.250 204.885 1726.410 ;
        RECT 205.055 1726.300 206.075 1726.630 ;
        RECT 201.995 1726.120 202.965 1726.250 ;
        RECT 202.165 1725.950 202.965 1726.120 ;
        RECT 201.995 1725.920 202.965 1725.950 ;
        RECT 203.565 1726.130 204.885 1726.250 ;
        RECT 203.565 1726.120 205.685 1726.130 ;
        RECT 203.565 1725.950 204.715 1726.120 ;
        RECT 204.885 1725.960 205.685 1726.120 ;
        RECT 203.565 1725.920 204.885 1725.950 ;
        RECT 201.995 1725.660 202.165 1725.920 ;
      LAYER li1 ;
        RECT 202.335 1725.580 204.545 1725.750 ;
      LAYER li1 ;
        RECT 204.715 1725.660 204.885 1725.920 ;
        RECT 205.905 1725.790 206.075 1726.300 ;
      LAYER li1 ;
        RECT 202.815 1725.495 203.695 1725.580 ;
      LAYER li1 ;
        RECT 201.995 1725.410 202.165 1725.490 ;
        RECT 201.995 1725.200 202.645 1725.410 ;
        RECT 202.165 1725.080 202.645 1725.200 ;
        RECT 201.995 1724.740 202.165 1725.030 ;
      LAYER li1 ;
        RECT 202.815 1724.910 202.985 1725.495 ;
        RECT 202.335 1724.740 202.985 1724.910 ;
      LAYER li1 ;
        RECT 201.995 1724.280 202.645 1724.570 ;
        RECT 202.165 1724.240 202.645 1724.280 ;
        RECT 201.995 1723.820 202.165 1724.110 ;
      LAYER li1 ;
        RECT 202.815 1724.070 202.985 1724.740 ;
        RECT 202.335 1723.900 202.985 1724.070 ;
      LAYER li1 ;
        RECT 202.165 1723.650 202.645 1723.730 ;
        RECT 201.995 1723.400 202.645 1723.650 ;
        RECT 201.995 1723.360 202.165 1723.400 ;
      LAYER li1 ;
        RECT 202.815 1723.230 202.985 1723.900 ;
      LAYER li1 ;
        RECT 201.995 1722.900 202.165 1723.190 ;
      LAYER li1 ;
        RECT 202.335 1723.060 202.985 1723.230 ;
      LAYER li1 ;
        RECT 202.165 1722.730 202.645 1722.890 ;
        RECT 203.155 1722.800 203.325 1725.250 ;
      LAYER li1 ;
        RECT 203.525 1724.910 203.695 1725.495 ;
      LAYER li1 ;
        RECT 204.715 1725.410 204.885 1725.490 ;
        RECT 205.055 1725.460 206.075 1725.790 ;
      LAYER li1 ;
        RECT 206.245 1725.485 206.445 1727.075 ;
      LAYER li1 ;
        RECT 206.710 1727.040 208.330 1727.100 ;
        RECT 206.710 1726.870 207.435 1727.040 ;
        RECT 207.605 1726.870 208.330 1727.040 ;
        RECT 206.710 1726.810 208.330 1726.870 ;
        RECT 208.990 1727.040 210.325 1727.100 ;
        RECT 208.990 1726.870 210.155 1727.040 ;
        RECT 208.990 1726.810 210.325 1726.870 ;
        RECT 207.435 1726.725 207.605 1726.810 ;
        RECT 210.155 1726.725 210.325 1726.810 ;
        RECT 206.615 1726.380 207.265 1726.550 ;
        RECT 206.615 1725.710 206.785 1726.380 ;
        RECT 206.955 1725.880 207.435 1726.210 ;
        RECT 206.615 1725.540 207.260 1725.710 ;
        RECT 203.915 1725.290 204.885 1725.410 ;
        RECT 205.905 1725.305 206.075 1725.460 ;
        RECT 206.615 1725.305 206.785 1725.540 ;
        RECT 203.915 1725.200 205.685 1725.290 ;
        RECT 203.915 1725.080 204.715 1725.200 ;
        RECT 204.885 1725.120 205.685 1725.200 ;
        RECT 205.905 1725.130 206.785 1725.305 ;
      LAYER li1 ;
        RECT 203.525 1724.740 204.545 1724.910 ;
      LAYER li1 ;
        RECT 204.715 1724.740 204.885 1725.030 ;
      LAYER li1 ;
        RECT 203.525 1724.070 203.695 1724.740 ;
        RECT 205.055 1724.700 206.075 1724.870 ;
      LAYER li1 ;
        RECT 203.915 1724.530 204.885 1724.570 ;
        RECT 203.915 1724.280 205.685 1724.530 ;
        RECT 203.915 1724.240 204.715 1724.280 ;
        RECT 204.885 1724.200 205.685 1724.280 ;
      LAYER li1 ;
        RECT 203.525 1723.900 204.545 1724.070 ;
        RECT 203.525 1723.230 203.695 1723.900 ;
      LAYER li1 ;
        RECT 204.715 1723.820 204.885 1724.110 ;
      LAYER li1 ;
        RECT 205.905 1724.030 206.075 1724.700 ;
        RECT 205.055 1723.860 206.075 1724.030 ;
      LAYER li1 ;
        RECT 203.915 1723.650 204.715 1723.730 ;
        RECT 204.885 1723.650 205.685 1723.690 ;
        RECT 203.915 1723.400 205.685 1723.650 ;
        RECT 204.715 1723.360 205.685 1723.400 ;
      LAYER li1 ;
        RECT 203.525 1723.060 204.545 1723.230 ;
        RECT 205.905 1723.190 206.075 1723.860 ;
      LAYER li1 ;
        RECT 204.715 1722.900 204.885 1723.190 ;
      LAYER li1 ;
        RECT 205.055 1723.020 206.075 1723.190 ;
      LAYER li1 ;
        RECT 201.995 1722.560 202.645 1722.730 ;
        RECT 202.815 1722.625 203.695 1722.800 ;
        RECT 203.915 1722.730 204.715 1722.810 ;
        RECT 204.885 1722.730 205.685 1722.850 ;
        RECT 203.915 1722.640 205.685 1722.730 ;
        RECT 201.995 1722.440 202.165 1722.560 ;
        RECT 202.815 1722.390 202.985 1722.625 ;
        RECT 203.525 1722.470 203.695 1722.625 ;
        RECT 204.715 1722.520 205.685 1722.640 ;
        RECT 201.995 1722.050 202.165 1722.270 ;
        RECT 202.340 1722.220 202.985 1722.390 ;
        RECT 201.995 1721.980 202.645 1722.050 ;
        RECT 202.165 1721.810 202.645 1721.980 ;
        RECT 201.995 1721.720 202.645 1721.810 ;
        RECT 201.995 1721.520 202.165 1721.720 ;
        RECT 202.815 1721.550 202.985 1722.220 ;
        RECT 202.335 1721.380 202.985 1721.550 ;
        RECT 201.995 1721.120 202.165 1721.350 ;
      LAYER li1 ;
        RECT 203.155 1721.345 203.355 1722.445 ;
      LAYER li1 ;
        RECT 203.525 1722.140 204.545 1722.470 ;
        RECT 204.715 1722.440 204.885 1722.520 ;
      LAYER li1 ;
        RECT 205.905 1722.435 206.075 1723.020 ;
      LAYER li1 ;
        RECT 206.275 1722.680 206.445 1725.130 ;
        RECT 206.955 1725.040 207.435 1725.370 ;
      LAYER li1 ;
        RECT 206.615 1724.700 207.265 1724.870 ;
        RECT 206.615 1724.030 206.785 1724.700 ;
      LAYER li1 ;
        RECT 206.955 1724.200 207.435 1724.530 ;
      LAYER li1 ;
        RECT 206.615 1723.860 207.265 1724.030 ;
        RECT 206.615 1723.190 206.785 1723.860 ;
      LAYER li1 ;
        RECT 206.955 1723.360 207.435 1723.690 ;
      LAYER li1 ;
        RECT 206.615 1723.020 207.265 1723.190 ;
        RECT 206.615 1722.435 206.785 1723.020 ;
      LAYER li1 ;
        RECT 206.955 1722.520 207.435 1722.850 ;
      LAYER li1 ;
        RECT 205.905 1722.350 206.785 1722.435 ;
      LAYER li1 ;
        RECT 203.525 1721.630 203.695 1722.140 ;
        RECT 204.715 1722.010 204.885 1722.270 ;
      LAYER li1 ;
        RECT 205.055 1722.180 207.265 1722.350 ;
      LAYER li1 ;
        RECT 204.715 1721.980 206.035 1722.010 ;
        RECT 203.915 1721.810 204.715 1721.970 ;
        RECT 204.885 1721.810 206.035 1721.980 ;
        RECT 203.915 1721.800 206.035 1721.810 ;
        RECT 204.715 1721.680 206.035 1721.800 ;
        RECT 206.635 1721.680 207.435 1722.010 ;
        RECT 203.525 1721.300 204.545 1721.630 ;
        RECT 204.715 1721.520 204.885 1721.680 ;
        RECT 204.715 1721.120 204.885 1721.350 ;
        RECT 207.435 1721.120 207.605 1721.205 ;
        RECT 210.155 1721.120 210.325 1721.205 ;
        RECT 201.995 1721.060 202.890 1721.120 ;
        RECT 202.165 1720.890 202.890 1721.060 ;
        RECT 201.995 1720.830 202.890 1720.890 ;
        RECT 203.550 1721.060 206.050 1721.120 ;
        RECT 203.550 1720.890 204.715 1721.060 ;
        RECT 204.885 1720.890 206.050 1721.060 ;
        RECT 203.550 1720.830 206.050 1720.890 ;
        RECT 201.995 1720.600 202.165 1720.830 ;
        RECT 204.715 1720.600 204.885 1720.830 ;
        RECT 201.995 1720.270 202.165 1720.430 ;
        RECT 204.715 1720.270 204.885 1720.430 ;
        RECT 205.055 1720.320 206.075 1720.650 ;
        RECT 201.995 1720.140 202.965 1720.270 ;
        RECT 202.165 1719.970 202.965 1720.140 ;
        RECT 201.995 1719.940 202.965 1719.970 ;
        RECT 203.565 1720.150 204.885 1720.270 ;
        RECT 203.565 1720.140 205.685 1720.150 ;
        RECT 203.565 1719.970 204.715 1720.140 ;
        RECT 204.885 1719.980 205.685 1720.140 ;
        RECT 203.565 1719.940 204.885 1719.970 ;
        RECT 201.995 1719.680 202.165 1719.940 ;
      LAYER li1 ;
        RECT 202.335 1719.600 204.545 1719.770 ;
      LAYER li1 ;
        RECT 204.715 1719.680 204.885 1719.940 ;
        RECT 205.905 1719.810 206.075 1720.320 ;
      LAYER li1 ;
        RECT 202.815 1719.515 203.695 1719.600 ;
      LAYER li1 ;
        RECT 201.995 1719.430 202.165 1719.510 ;
        RECT 201.995 1719.220 202.645 1719.430 ;
        RECT 202.165 1719.100 202.645 1719.220 ;
        RECT 201.995 1718.760 202.165 1719.050 ;
      LAYER li1 ;
        RECT 202.815 1718.930 202.985 1719.515 ;
        RECT 202.335 1718.760 202.985 1718.930 ;
      LAYER li1 ;
        RECT 201.995 1718.300 202.645 1718.590 ;
        RECT 202.165 1718.260 202.645 1718.300 ;
        RECT 201.995 1717.840 202.165 1718.130 ;
      LAYER li1 ;
        RECT 202.815 1718.090 202.985 1718.760 ;
        RECT 202.335 1717.920 202.985 1718.090 ;
      LAYER li1 ;
        RECT 202.165 1717.670 202.645 1717.750 ;
        RECT 201.995 1717.420 202.645 1717.670 ;
        RECT 201.995 1717.380 202.165 1717.420 ;
      LAYER li1 ;
        RECT 202.815 1717.250 202.985 1717.920 ;
      LAYER li1 ;
        RECT 201.995 1716.920 202.165 1717.210 ;
      LAYER li1 ;
        RECT 202.335 1717.080 202.985 1717.250 ;
      LAYER li1 ;
        RECT 202.165 1716.750 202.645 1716.910 ;
        RECT 203.155 1716.820 203.325 1719.270 ;
      LAYER li1 ;
        RECT 203.525 1718.930 203.695 1719.515 ;
      LAYER li1 ;
        RECT 204.715 1719.430 204.885 1719.510 ;
        RECT 205.055 1719.480 206.075 1719.810 ;
      LAYER li1 ;
        RECT 206.245 1719.505 206.445 1721.095 ;
      LAYER li1 ;
        RECT 206.710 1721.060 208.330 1721.120 ;
        RECT 206.710 1720.890 207.435 1721.060 ;
        RECT 207.605 1720.890 208.330 1721.060 ;
        RECT 206.710 1720.830 208.330 1720.890 ;
        RECT 208.990 1721.060 210.325 1721.120 ;
        RECT 208.990 1720.890 210.155 1721.060 ;
        RECT 208.990 1720.830 210.325 1720.890 ;
        RECT 207.435 1720.745 207.605 1720.830 ;
        RECT 210.155 1720.745 210.325 1720.830 ;
        RECT 206.615 1720.400 207.265 1720.570 ;
        RECT 206.615 1719.730 206.785 1720.400 ;
        RECT 206.955 1719.900 207.435 1720.230 ;
        RECT 206.615 1719.560 207.260 1719.730 ;
        RECT 203.915 1719.310 204.885 1719.430 ;
        RECT 205.905 1719.325 206.075 1719.480 ;
        RECT 206.615 1719.325 206.785 1719.560 ;
        RECT 203.915 1719.220 205.685 1719.310 ;
        RECT 203.915 1719.100 204.715 1719.220 ;
        RECT 204.885 1719.140 205.685 1719.220 ;
        RECT 205.905 1719.150 206.785 1719.325 ;
      LAYER li1 ;
        RECT 203.525 1718.760 204.545 1718.930 ;
      LAYER li1 ;
        RECT 204.715 1718.760 204.885 1719.050 ;
      LAYER li1 ;
        RECT 203.525 1718.090 203.695 1718.760 ;
        RECT 205.055 1718.720 206.075 1718.890 ;
      LAYER li1 ;
        RECT 203.915 1718.550 204.885 1718.590 ;
        RECT 203.915 1718.300 205.685 1718.550 ;
        RECT 203.915 1718.260 204.715 1718.300 ;
        RECT 204.885 1718.220 205.685 1718.300 ;
      LAYER li1 ;
        RECT 203.525 1717.920 204.545 1718.090 ;
        RECT 203.525 1717.250 203.695 1717.920 ;
      LAYER li1 ;
        RECT 204.715 1717.840 204.885 1718.130 ;
      LAYER li1 ;
        RECT 205.905 1718.050 206.075 1718.720 ;
        RECT 205.055 1717.880 206.075 1718.050 ;
      LAYER li1 ;
        RECT 203.915 1717.670 204.715 1717.750 ;
        RECT 204.885 1717.670 205.685 1717.710 ;
        RECT 203.915 1717.420 205.685 1717.670 ;
        RECT 204.715 1717.380 205.685 1717.420 ;
      LAYER li1 ;
        RECT 203.525 1717.080 204.545 1717.250 ;
        RECT 205.905 1717.210 206.075 1717.880 ;
      LAYER li1 ;
        RECT 204.715 1716.920 204.885 1717.210 ;
      LAYER li1 ;
        RECT 205.055 1717.040 206.075 1717.210 ;
      LAYER li1 ;
        RECT 201.995 1716.580 202.645 1716.750 ;
        RECT 202.815 1716.645 203.695 1716.820 ;
        RECT 203.915 1716.750 204.715 1716.830 ;
        RECT 204.885 1716.750 205.685 1716.870 ;
        RECT 203.915 1716.660 205.685 1716.750 ;
        RECT 201.995 1716.460 202.165 1716.580 ;
        RECT 202.815 1716.410 202.985 1716.645 ;
        RECT 203.525 1716.490 203.695 1716.645 ;
        RECT 204.715 1716.540 205.685 1716.660 ;
        RECT 201.995 1716.070 202.165 1716.290 ;
        RECT 202.340 1716.240 202.985 1716.410 ;
        RECT 201.995 1716.000 202.645 1716.070 ;
        RECT 202.165 1715.830 202.645 1716.000 ;
        RECT 201.995 1715.740 202.645 1715.830 ;
        RECT 201.995 1715.540 202.165 1715.740 ;
        RECT 202.815 1715.570 202.985 1716.240 ;
        RECT 202.335 1715.400 202.985 1715.570 ;
        RECT 201.995 1715.140 202.165 1715.370 ;
      LAYER li1 ;
        RECT 203.155 1715.365 203.355 1716.465 ;
      LAYER li1 ;
        RECT 203.525 1716.160 204.545 1716.490 ;
        RECT 204.715 1716.460 204.885 1716.540 ;
      LAYER li1 ;
        RECT 205.905 1716.455 206.075 1717.040 ;
      LAYER li1 ;
        RECT 206.275 1716.700 206.445 1719.150 ;
        RECT 206.955 1719.060 207.435 1719.390 ;
      LAYER li1 ;
        RECT 206.615 1718.720 207.265 1718.890 ;
        RECT 206.615 1718.050 206.785 1718.720 ;
      LAYER li1 ;
        RECT 206.955 1718.220 207.435 1718.550 ;
      LAYER li1 ;
        RECT 206.615 1717.880 207.265 1718.050 ;
        RECT 206.615 1717.210 206.785 1717.880 ;
      LAYER li1 ;
        RECT 206.955 1717.380 207.435 1717.710 ;
      LAYER li1 ;
        RECT 206.615 1717.040 207.265 1717.210 ;
        RECT 206.615 1716.455 206.785 1717.040 ;
      LAYER li1 ;
        RECT 206.955 1716.540 207.435 1716.870 ;
      LAYER li1 ;
        RECT 205.905 1716.370 206.785 1716.455 ;
      LAYER li1 ;
        RECT 203.525 1715.650 203.695 1716.160 ;
        RECT 204.715 1716.030 204.885 1716.290 ;
      LAYER li1 ;
        RECT 205.055 1716.200 207.265 1716.370 ;
      LAYER li1 ;
        RECT 204.715 1716.000 206.035 1716.030 ;
        RECT 203.915 1715.830 204.715 1715.990 ;
        RECT 204.885 1715.830 206.035 1716.000 ;
        RECT 203.915 1715.820 206.035 1715.830 ;
        RECT 204.715 1715.700 206.035 1715.820 ;
        RECT 206.635 1715.700 207.435 1716.030 ;
        RECT 203.525 1715.320 204.545 1715.650 ;
        RECT 204.715 1715.540 204.885 1715.700 ;
        RECT 204.715 1715.140 204.885 1715.370 ;
        RECT 207.435 1715.140 207.605 1715.225 ;
        RECT 210.155 1715.140 210.325 1715.225 ;
        RECT 201.995 1715.080 202.890 1715.140 ;
        RECT 202.165 1714.910 202.890 1715.080 ;
        RECT 201.995 1714.850 202.890 1714.910 ;
        RECT 203.550 1715.080 206.050 1715.140 ;
        RECT 203.550 1714.910 204.715 1715.080 ;
        RECT 204.885 1714.910 206.050 1715.080 ;
        RECT 203.550 1714.850 206.050 1714.910 ;
        RECT 201.995 1714.620 202.165 1714.850 ;
        RECT 204.715 1714.620 204.885 1714.850 ;
        RECT 201.995 1714.290 202.165 1714.450 ;
        RECT 204.715 1714.290 204.885 1714.450 ;
        RECT 205.055 1714.340 206.075 1714.670 ;
        RECT 201.995 1714.160 202.965 1714.290 ;
        RECT 202.165 1713.990 202.965 1714.160 ;
        RECT 201.995 1713.960 202.965 1713.990 ;
        RECT 203.565 1714.170 204.885 1714.290 ;
        RECT 203.565 1714.160 205.685 1714.170 ;
        RECT 203.565 1713.990 204.715 1714.160 ;
        RECT 204.885 1714.000 205.685 1714.160 ;
        RECT 203.565 1713.960 204.885 1713.990 ;
        RECT 201.995 1713.700 202.165 1713.960 ;
      LAYER li1 ;
        RECT 202.335 1713.620 204.545 1713.790 ;
      LAYER li1 ;
        RECT 204.715 1713.700 204.885 1713.960 ;
        RECT 205.905 1713.830 206.075 1714.340 ;
      LAYER li1 ;
        RECT 202.815 1713.535 203.695 1713.620 ;
      LAYER li1 ;
        RECT 201.995 1713.450 202.165 1713.530 ;
        RECT 201.995 1713.240 202.645 1713.450 ;
        RECT 202.165 1713.120 202.645 1713.240 ;
        RECT 201.995 1712.780 202.165 1713.070 ;
      LAYER li1 ;
        RECT 202.815 1712.950 202.985 1713.535 ;
        RECT 202.335 1712.780 202.985 1712.950 ;
      LAYER li1 ;
        RECT 201.995 1712.320 202.645 1712.610 ;
        RECT 202.165 1712.280 202.645 1712.320 ;
        RECT 201.995 1711.860 202.165 1712.150 ;
      LAYER li1 ;
        RECT 202.815 1712.110 202.985 1712.780 ;
        RECT 202.335 1711.940 202.985 1712.110 ;
      LAYER li1 ;
        RECT 202.165 1711.690 202.645 1711.770 ;
        RECT 201.995 1711.440 202.645 1711.690 ;
        RECT 201.995 1711.400 202.165 1711.440 ;
      LAYER li1 ;
        RECT 202.815 1711.270 202.985 1711.940 ;
      LAYER li1 ;
        RECT 201.995 1710.940 202.165 1711.230 ;
      LAYER li1 ;
        RECT 202.335 1711.100 202.985 1711.270 ;
      LAYER li1 ;
        RECT 202.165 1710.770 202.645 1710.930 ;
        RECT 203.155 1710.840 203.325 1713.290 ;
      LAYER li1 ;
        RECT 203.525 1712.950 203.695 1713.535 ;
      LAYER li1 ;
        RECT 204.715 1713.450 204.885 1713.530 ;
        RECT 205.055 1713.500 206.075 1713.830 ;
      LAYER li1 ;
        RECT 206.245 1713.525 206.445 1715.115 ;
      LAYER li1 ;
        RECT 206.710 1715.080 208.330 1715.140 ;
        RECT 206.710 1714.910 207.435 1715.080 ;
        RECT 207.605 1714.910 208.330 1715.080 ;
        RECT 206.710 1714.850 208.330 1714.910 ;
        RECT 208.990 1715.080 210.325 1715.140 ;
        RECT 208.990 1714.910 210.155 1715.080 ;
        RECT 208.990 1714.850 210.325 1714.910 ;
        RECT 207.435 1714.765 207.605 1714.850 ;
        RECT 210.155 1714.765 210.325 1714.850 ;
        RECT 206.615 1714.420 207.265 1714.590 ;
        RECT 206.615 1713.750 206.785 1714.420 ;
        RECT 206.955 1713.920 207.435 1714.250 ;
        RECT 206.615 1713.580 207.260 1713.750 ;
        RECT 203.915 1713.330 204.885 1713.450 ;
        RECT 205.905 1713.345 206.075 1713.500 ;
        RECT 206.615 1713.345 206.785 1713.580 ;
        RECT 203.915 1713.240 205.685 1713.330 ;
        RECT 203.915 1713.120 204.715 1713.240 ;
        RECT 204.885 1713.160 205.685 1713.240 ;
        RECT 205.905 1713.170 206.785 1713.345 ;
      LAYER li1 ;
        RECT 203.525 1712.780 204.545 1712.950 ;
      LAYER li1 ;
        RECT 204.715 1712.780 204.885 1713.070 ;
      LAYER li1 ;
        RECT 203.525 1712.110 203.695 1712.780 ;
        RECT 205.055 1712.740 206.075 1712.910 ;
      LAYER li1 ;
        RECT 203.915 1712.570 204.885 1712.610 ;
        RECT 203.915 1712.320 205.685 1712.570 ;
        RECT 203.915 1712.280 204.715 1712.320 ;
        RECT 204.885 1712.240 205.685 1712.320 ;
      LAYER li1 ;
        RECT 203.525 1711.940 204.545 1712.110 ;
        RECT 203.525 1711.270 203.695 1711.940 ;
      LAYER li1 ;
        RECT 204.715 1711.860 204.885 1712.150 ;
      LAYER li1 ;
        RECT 205.905 1712.070 206.075 1712.740 ;
        RECT 205.055 1711.900 206.075 1712.070 ;
      LAYER li1 ;
        RECT 203.915 1711.690 204.715 1711.770 ;
        RECT 204.885 1711.690 205.685 1711.730 ;
        RECT 203.915 1711.440 205.685 1711.690 ;
        RECT 204.715 1711.400 205.685 1711.440 ;
      LAYER li1 ;
        RECT 203.525 1711.100 204.545 1711.270 ;
        RECT 205.905 1711.230 206.075 1711.900 ;
      LAYER li1 ;
        RECT 204.715 1710.940 204.885 1711.230 ;
      LAYER li1 ;
        RECT 205.055 1711.060 206.075 1711.230 ;
      LAYER li1 ;
        RECT 201.995 1710.600 202.645 1710.770 ;
        RECT 202.815 1710.665 203.695 1710.840 ;
        RECT 203.915 1710.770 204.715 1710.850 ;
        RECT 204.885 1710.770 205.685 1710.890 ;
        RECT 203.915 1710.680 205.685 1710.770 ;
        RECT 201.995 1710.480 202.165 1710.600 ;
        RECT 202.815 1710.430 202.985 1710.665 ;
        RECT 203.525 1710.510 203.695 1710.665 ;
        RECT 204.715 1710.560 205.685 1710.680 ;
        RECT 201.995 1710.090 202.165 1710.310 ;
        RECT 202.340 1710.260 202.985 1710.430 ;
        RECT 201.995 1710.020 202.645 1710.090 ;
        RECT 202.165 1709.850 202.645 1710.020 ;
        RECT 201.995 1709.760 202.645 1709.850 ;
        RECT 201.995 1709.560 202.165 1709.760 ;
        RECT 202.815 1709.590 202.985 1710.260 ;
        RECT 202.335 1709.420 202.985 1709.590 ;
        RECT 201.995 1709.160 202.165 1709.390 ;
      LAYER li1 ;
        RECT 203.155 1709.385 203.355 1710.485 ;
      LAYER li1 ;
        RECT 203.525 1710.180 204.545 1710.510 ;
        RECT 204.715 1710.480 204.885 1710.560 ;
      LAYER li1 ;
        RECT 205.905 1710.475 206.075 1711.060 ;
      LAYER li1 ;
        RECT 206.275 1710.720 206.445 1713.170 ;
        RECT 206.955 1713.080 207.435 1713.410 ;
      LAYER li1 ;
        RECT 206.615 1712.740 207.265 1712.910 ;
        RECT 206.615 1712.070 206.785 1712.740 ;
      LAYER li1 ;
        RECT 206.955 1712.240 207.435 1712.570 ;
      LAYER li1 ;
        RECT 206.615 1711.900 207.265 1712.070 ;
        RECT 206.615 1711.230 206.785 1711.900 ;
      LAYER li1 ;
        RECT 206.955 1711.400 207.435 1711.730 ;
      LAYER li1 ;
        RECT 206.615 1711.060 207.265 1711.230 ;
        RECT 206.615 1710.475 206.785 1711.060 ;
      LAYER li1 ;
        RECT 206.955 1710.560 207.435 1710.890 ;
      LAYER li1 ;
        RECT 205.905 1710.390 206.785 1710.475 ;
      LAYER li1 ;
        RECT 203.525 1709.670 203.695 1710.180 ;
        RECT 204.715 1710.050 204.885 1710.310 ;
      LAYER li1 ;
        RECT 205.055 1710.220 207.265 1710.390 ;
      LAYER li1 ;
        RECT 204.715 1710.020 206.035 1710.050 ;
        RECT 203.915 1709.850 204.715 1710.010 ;
        RECT 204.885 1709.850 206.035 1710.020 ;
        RECT 203.915 1709.840 206.035 1709.850 ;
        RECT 204.715 1709.720 206.035 1709.840 ;
        RECT 206.635 1709.720 207.435 1710.050 ;
        RECT 203.525 1709.340 204.545 1709.670 ;
        RECT 204.715 1709.560 204.885 1709.720 ;
        RECT 204.715 1709.160 204.885 1709.390 ;
        RECT 207.435 1709.160 207.605 1709.245 ;
        RECT 210.155 1709.160 210.325 1709.245 ;
        RECT 201.995 1709.100 202.890 1709.160 ;
        RECT 202.165 1708.930 202.890 1709.100 ;
        RECT 201.995 1708.870 202.890 1708.930 ;
        RECT 203.550 1709.100 206.050 1709.160 ;
        RECT 203.550 1708.930 204.715 1709.100 ;
        RECT 204.885 1708.930 206.050 1709.100 ;
        RECT 203.550 1708.870 206.050 1708.930 ;
        RECT 201.995 1708.640 202.165 1708.870 ;
        RECT 204.715 1708.640 204.885 1708.870 ;
        RECT 201.995 1708.310 202.165 1708.470 ;
        RECT 204.715 1708.310 204.885 1708.470 ;
        RECT 205.055 1708.360 206.075 1708.690 ;
        RECT 201.995 1708.180 202.965 1708.310 ;
        RECT 202.165 1708.010 202.965 1708.180 ;
        RECT 201.995 1707.980 202.965 1708.010 ;
        RECT 203.565 1708.190 204.885 1708.310 ;
        RECT 203.565 1708.180 205.685 1708.190 ;
        RECT 203.565 1708.010 204.715 1708.180 ;
        RECT 204.885 1708.020 205.685 1708.180 ;
        RECT 203.565 1707.980 204.885 1708.010 ;
        RECT 201.995 1707.720 202.165 1707.980 ;
      LAYER li1 ;
        RECT 202.335 1707.640 204.545 1707.810 ;
      LAYER li1 ;
        RECT 204.715 1707.720 204.885 1707.980 ;
        RECT 205.905 1707.850 206.075 1708.360 ;
      LAYER li1 ;
        RECT 202.815 1707.555 203.695 1707.640 ;
      LAYER li1 ;
        RECT 201.995 1707.470 202.165 1707.550 ;
        RECT 201.995 1707.260 202.645 1707.470 ;
        RECT 202.165 1707.140 202.645 1707.260 ;
        RECT 201.995 1706.800 202.165 1707.090 ;
      LAYER li1 ;
        RECT 202.815 1706.970 202.985 1707.555 ;
        RECT 202.335 1706.800 202.985 1706.970 ;
      LAYER li1 ;
        RECT 201.995 1706.340 202.645 1706.630 ;
        RECT 202.165 1706.300 202.645 1706.340 ;
        RECT 201.995 1705.880 202.165 1706.170 ;
      LAYER li1 ;
        RECT 202.815 1706.130 202.985 1706.800 ;
        RECT 202.335 1705.960 202.985 1706.130 ;
      LAYER li1 ;
        RECT 202.165 1705.710 202.645 1705.790 ;
        RECT 201.995 1705.460 202.645 1705.710 ;
        RECT 201.995 1705.420 202.165 1705.460 ;
      LAYER li1 ;
        RECT 202.815 1705.290 202.985 1705.960 ;
      LAYER li1 ;
        RECT 201.995 1704.960 202.165 1705.250 ;
      LAYER li1 ;
        RECT 202.335 1705.120 202.985 1705.290 ;
      LAYER li1 ;
        RECT 202.165 1704.790 202.645 1704.950 ;
        RECT 203.155 1704.860 203.325 1707.310 ;
      LAYER li1 ;
        RECT 203.525 1706.970 203.695 1707.555 ;
      LAYER li1 ;
        RECT 204.715 1707.470 204.885 1707.550 ;
        RECT 205.055 1707.520 206.075 1707.850 ;
      LAYER li1 ;
        RECT 206.245 1707.545 206.445 1709.135 ;
      LAYER li1 ;
        RECT 206.710 1709.100 208.330 1709.160 ;
        RECT 206.710 1708.930 207.435 1709.100 ;
        RECT 207.605 1708.930 208.330 1709.100 ;
        RECT 206.710 1708.870 208.330 1708.930 ;
        RECT 208.990 1709.100 210.325 1709.160 ;
        RECT 208.990 1708.930 210.155 1709.100 ;
        RECT 208.990 1708.870 210.325 1708.930 ;
        RECT 207.435 1708.785 207.605 1708.870 ;
        RECT 210.155 1708.785 210.325 1708.870 ;
        RECT 206.615 1708.440 207.265 1708.610 ;
        RECT 206.615 1707.770 206.785 1708.440 ;
        RECT 206.955 1707.940 207.435 1708.270 ;
        RECT 206.615 1707.600 207.260 1707.770 ;
        RECT 203.915 1707.350 204.885 1707.470 ;
        RECT 205.905 1707.365 206.075 1707.520 ;
        RECT 206.615 1707.365 206.785 1707.600 ;
        RECT 203.915 1707.260 205.685 1707.350 ;
        RECT 203.915 1707.140 204.715 1707.260 ;
        RECT 204.885 1707.180 205.685 1707.260 ;
        RECT 205.905 1707.190 206.785 1707.365 ;
      LAYER li1 ;
        RECT 203.525 1706.800 204.545 1706.970 ;
      LAYER li1 ;
        RECT 204.715 1706.800 204.885 1707.090 ;
      LAYER li1 ;
        RECT 203.525 1706.130 203.695 1706.800 ;
        RECT 205.055 1706.760 206.075 1706.930 ;
      LAYER li1 ;
        RECT 203.915 1706.590 204.885 1706.630 ;
        RECT 203.915 1706.340 205.685 1706.590 ;
        RECT 203.915 1706.300 204.715 1706.340 ;
        RECT 204.885 1706.260 205.685 1706.340 ;
      LAYER li1 ;
        RECT 203.525 1705.960 204.545 1706.130 ;
        RECT 203.525 1705.290 203.695 1705.960 ;
      LAYER li1 ;
        RECT 204.715 1705.880 204.885 1706.170 ;
      LAYER li1 ;
        RECT 205.905 1706.090 206.075 1706.760 ;
        RECT 205.055 1705.920 206.075 1706.090 ;
      LAYER li1 ;
        RECT 203.915 1705.710 204.715 1705.790 ;
        RECT 204.885 1705.710 205.685 1705.750 ;
        RECT 203.915 1705.460 205.685 1705.710 ;
        RECT 204.715 1705.420 205.685 1705.460 ;
      LAYER li1 ;
        RECT 203.525 1705.120 204.545 1705.290 ;
        RECT 205.905 1705.250 206.075 1705.920 ;
      LAYER li1 ;
        RECT 204.715 1704.960 204.885 1705.250 ;
      LAYER li1 ;
        RECT 205.055 1705.080 206.075 1705.250 ;
      LAYER li1 ;
        RECT 201.995 1704.620 202.645 1704.790 ;
        RECT 202.815 1704.685 203.695 1704.860 ;
        RECT 203.915 1704.790 204.715 1704.870 ;
        RECT 204.885 1704.790 205.685 1704.910 ;
        RECT 203.915 1704.700 205.685 1704.790 ;
        RECT 201.995 1704.500 202.165 1704.620 ;
        RECT 202.815 1704.450 202.985 1704.685 ;
        RECT 203.525 1704.530 203.695 1704.685 ;
        RECT 204.715 1704.580 205.685 1704.700 ;
        RECT 201.995 1704.110 202.165 1704.330 ;
        RECT 202.340 1704.280 202.985 1704.450 ;
        RECT 201.995 1704.040 202.645 1704.110 ;
        RECT 202.165 1703.870 202.645 1704.040 ;
        RECT 201.995 1703.780 202.645 1703.870 ;
        RECT 201.995 1703.580 202.165 1703.780 ;
        RECT 202.815 1703.610 202.985 1704.280 ;
        RECT 202.335 1703.440 202.985 1703.610 ;
        RECT 201.995 1703.180 202.165 1703.410 ;
      LAYER li1 ;
        RECT 203.155 1703.405 203.355 1704.505 ;
      LAYER li1 ;
        RECT 203.525 1704.200 204.545 1704.530 ;
        RECT 204.715 1704.500 204.885 1704.580 ;
      LAYER li1 ;
        RECT 205.905 1704.495 206.075 1705.080 ;
      LAYER li1 ;
        RECT 206.275 1704.740 206.445 1707.190 ;
        RECT 206.955 1707.100 207.435 1707.430 ;
      LAYER li1 ;
        RECT 206.615 1706.760 207.265 1706.930 ;
        RECT 206.615 1706.090 206.785 1706.760 ;
      LAYER li1 ;
        RECT 206.955 1706.260 207.435 1706.590 ;
      LAYER li1 ;
        RECT 206.615 1705.920 207.265 1706.090 ;
        RECT 206.615 1705.250 206.785 1705.920 ;
      LAYER li1 ;
        RECT 206.955 1705.420 207.435 1705.750 ;
      LAYER li1 ;
        RECT 206.615 1705.080 207.265 1705.250 ;
        RECT 206.615 1704.495 206.785 1705.080 ;
      LAYER li1 ;
        RECT 206.955 1704.580 207.435 1704.910 ;
      LAYER li1 ;
        RECT 205.905 1704.410 206.785 1704.495 ;
      LAYER li1 ;
        RECT 203.525 1703.690 203.695 1704.200 ;
        RECT 204.715 1704.070 204.885 1704.330 ;
      LAYER li1 ;
        RECT 205.055 1704.240 207.265 1704.410 ;
      LAYER li1 ;
        RECT 204.715 1704.040 206.035 1704.070 ;
        RECT 203.915 1703.870 204.715 1704.030 ;
        RECT 204.885 1703.870 206.035 1704.040 ;
        RECT 203.915 1703.860 206.035 1703.870 ;
        RECT 204.715 1703.740 206.035 1703.860 ;
        RECT 206.635 1703.740 207.435 1704.070 ;
        RECT 203.525 1703.360 204.545 1703.690 ;
        RECT 204.715 1703.580 204.885 1703.740 ;
        RECT 204.715 1703.180 204.885 1703.410 ;
        RECT 207.435 1703.180 207.605 1703.265 ;
        RECT 210.155 1703.180 210.325 1703.265 ;
        RECT 201.995 1703.120 202.890 1703.180 ;
        RECT 202.165 1702.950 202.890 1703.120 ;
        RECT 201.995 1702.890 202.890 1702.950 ;
        RECT 203.550 1703.120 206.050 1703.180 ;
        RECT 203.550 1702.950 204.715 1703.120 ;
        RECT 204.885 1702.950 206.050 1703.120 ;
        RECT 203.550 1702.890 206.050 1702.950 ;
        RECT 201.995 1702.660 202.165 1702.890 ;
        RECT 204.715 1702.660 204.885 1702.890 ;
        RECT 201.995 1702.330 202.165 1702.490 ;
        RECT 204.715 1702.330 204.885 1702.490 ;
        RECT 205.055 1702.380 206.075 1702.710 ;
        RECT 201.995 1702.200 202.965 1702.330 ;
        RECT 202.165 1702.030 202.965 1702.200 ;
        RECT 201.995 1702.000 202.965 1702.030 ;
        RECT 203.565 1702.210 204.885 1702.330 ;
        RECT 203.565 1702.200 205.685 1702.210 ;
        RECT 203.565 1702.030 204.715 1702.200 ;
        RECT 204.885 1702.040 205.685 1702.200 ;
        RECT 203.565 1702.000 204.885 1702.030 ;
        RECT 201.995 1701.740 202.165 1702.000 ;
      LAYER li1 ;
        RECT 202.335 1701.660 204.545 1701.830 ;
      LAYER li1 ;
        RECT 204.715 1701.740 204.885 1702.000 ;
        RECT 205.905 1701.870 206.075 1702.380 ;
      LAYER li1 ;
        RECT 202.815 1701.575 203.695 1701.660 ;
      LAYER li1 ;
        RECT 201.995 1701.490 202.165 1701.570 ;
        RECT 201.995 1701.280 202.645 1701.490 ;
        RECT 202.165 1701.160 202.645 1701.280 ;
        RECT 201.995 1700.820 202.165 1701.110 ;
      LAYER li1 ;
        RECT 202.815 1700.990 202.985 1701.575 ;
        RECT 202.335 1700.820 202.985 1700.990 ;
      LAYER li1 ;
        RECT 201.995 1700.360 202.645 1700.650 ;
        RECT 202.165 1700.320 202.645 1700.360 ;
        RECT 201.995 1699.900 202.165 1700.190 ;
      LAYER li1 ;
        RECT 202.815 1700.150 202.985 1700.820 ;
        RECT 202.335 1699.980 202.985 1700.150 ;
      LAYER li1 ;
        RECT 202.165 1699.730 202.645 1699.810 ;
        RECT 201.995 1699.480 202.645 1699.730 ;
        RECT 201.995 1699.440 202.165 1699.480 ;
      LAYER li1 ;
        RECT 202.815 1699.310 202.985 1699.980 ;
      LAYER li1 ;
        RECT 201.995 1698.980 202.165 1699.270 ;
      LAYER li1 ;
        RECT 202.335 1699.140 202.985 1699.310 ;
      LAYER li1 ;
        RECT 202.165 1698.810 202.645 1698.970 ;
        RECT 203.155 1698.880 203.325 1701.330 ;
      LAYER li1 ;
        RECT 203.525 1700.990 203.695 1701.575 ;
      LAYER li1 ;
        RECT 204.715 1701.490 204.885 1701.570 ;
        RECT 205.055 1701.540 206.075 1701.870 ;
      LAYER li1 ;
        RECT 206.245 1701.565 206.445 1703.155 ;
      LAYER li1 ;
        RECT 206.710 1703.120 208.330 1703.180 ;
        RECT 206.710 1702.950 207.435 1703.120 ;
        RECT 207.605 1702.950 208.330 1703.120 ;
        RECT 206.710 1702.890 208.330 1702.950 ;
        RECT 208.990 1703.120 210.325 1703.180 ;
        RECT 208.990 1702.950 210.155 1703.120 ;
        RECT 208.990 1702.890 210.325 1702.950 ;
        RECT 207.435 1702.805 207.605 1702.890 ;
        RECT 210.155 1702.805 210.325 1702.890 ;
        RECT 206.615 1702.460 207.265 1702.630 ;
        RECT 206.615 1701.790 206.785 1702.460 ;
        RECT 206.955 1701.960 207.435 1702.290 ;
        RECT 206.615 1701.620 207.260 1701.790 ;
        RECT 203.915 1701.370 204.885 1701.490 ;
        RECT 205.905 1701.385 206.075 1701.540 ;
        RECT 206.615 1701.385 206.785 1701.620 ;
        RECT 203.915 1701.280 205.685 1701.370 ;
        RECT 203.915 1701.160 204.715 1701.280 ;
        RECT 204.885 1701.200 205.685 1701.280 ;
        RECT 205.905 1701.210 206.785 1701.385 ;
      LAYER li1 ;
        RECT 203.525 1700.820 204.545 1700.990 ;
      LAYER li1 ;
        RECT 204.715 1700.820 204.885 1701.110 ;
      LAYER li1 ;
        RECT 203.525 1700.150 203.695 1700.820 ;
        RECT 205.055 1700.780 206.075 1700.950 ;
      LAYER li1 ;
        RECT 203.915 1700.610 204.885 1700.650 ;
        RECT 203.915 1700.360 205.685 1700.610 ;
        RECT 203.915 1700.320 204.715 1700.360 ;
        RECT 204.885 1700.280 205.685 1700.360 ;
      LAYER li1 ;
        RECT 203.525 1699.980 204.545 1700.150 ;
        RECT 203.525 1699.310 203.695 1699.980 ;
      LAYER li1 ;
        RECT 204.715 1699.900 204.885 1700.190 ;
      LAYER li1 ;
        RECT 205.905 1700.110 206.075 1700.780 ;
        RECT 205.055 1699.940 206.075 1700.110 ;
      LAYER li1 ;
        RECT 203.915 1699.730 204.715 1699.810 ;
        RECT 204.885 1699.730 205.685 1699.770 ;
        RECT 203.915 1699.480 205.685 1699.730 ;
        RECT 204.715 1699.440 205.685 1699.480 ;
      LAYER li1 ;
        RECT 203.525 1699.140 204.545 1699.310 ;
        RECT 205.905 1699.270 206.075 1699.940 ;
      LAYER li1 ;
        RECT 204.715 1698.980 204.885 1699.270 ;
      LAYER li1 ;
        RECT 205.055 1699.100 206.075 1699.270 ;
      LAYER li1 ;
        RECT 201.995 1698.640 202.645 1698.810 ;
        RECT 202.815 1698.705 203.695 1698.880 ;
        RECT 203.915 1698.810 204.715 1698.890 ;
        RECT 204.885 1698.810 205.685 1698.930 ;
        RECT 203.915 1698.720 205.685 1698.810 ;
        RECT 201.995 1698.520 202.165 1698.640 ;
        RECT 202.815 1698.470 202.985 1698.705 ;
        RECT 203.525 1698.550 203.695 1698.705 ;
        RECT 204.715 1698.600 205.685 1698.720 ;
        RECT 201.995 1698.130 202.165 1698.350 ;
        RECT 202.340 1698.300 202.985 1698.470 ;
        RECT 201.995 1698.060 202.645 1698.130 ;
        RECT 202.165 1697.890 202.645 1698.060 ;
        RECT 201.995 1697.800 202.645 1697.890 ;
        RECT 201.995 1697.600 202.165 1697.800 ;
        RECT 202.815 1697.630 202.985 1698.300 ;
        RECT 202.335 1697.460 202.985 1697.630 ;
        RECT 201.995 1697.200 202.165 1697.430 ;
      LAYER li1 ;
        RECT 203.155 1697.425 203.355 1698.525 ;
      LAYER li1 ;
        RECT 203.525 1698.220 204.545 1698.550 ;
        RECT 204.715 1698.520 204.885 1698.600 ;
      LAYER li1 ;
        RECT 205.905 1698.515 206.075 1699.100 ;
      LAYER li1 ;
        RECT 206.275 1698.760 206.445 1701.210 ;
        RECT 206.955 1701.120 207.435 1701.450 ;
      LAYER li1 ;
        RECT 206.615 1700.780 207.265 1700.950 ;
        RECT 206.615 1700.110 206.785 1700.780 ;
      LAYER li1 ;
        RECT 206.955 1700.280 207.435 1700.610 ;
      LAYER li1 ;
        RECT 206.615 1699.940 207.265 1700.110 ;
        RECT 206.615 1699.270 206.785 1699.940 ;
      LAYER li1 ;
        RECT 206.955 1699.440 207.435 1699.770 ;
      LAYER li1 ;
        RECT 206.615 1699.100 207.265 1699.270 ;
        RECT 206.615 1698.515 206.785 1699.100 ;
      LAYER li1 ;
        RECT 206.955 1698.600 207.435 1698.930 ;
      LAYER li1 ;
        RECT 205.905 1698.430 206.785 1698.515 ;
      LAYER li1 ;
        RECT 203.525 1697.710 203.695 1698.220 ;
        RECT 204.715 1698.090 204.885 1698.350 ;
      LAYER li1 ;
        RECT 205.055 1698.260 207.265 1698.430 ;
      LAYER li1 ;
        RECT 204.715 1698.060 206.035 1698.090 ;
        RECT 203.915 1697.890 204.715 1698.050 ;
        RECT 204.885 1697.890 206.035 1698.060 ;
        RECT 203.915 1697.880 206.035 1697.890 ;
        RECT 204.715 1697.760 206.035 1697.880 ;
        RECT 206.635 1697.760 207.435 1698.090 ;
        RECT 203.525 1697.380 204.545 1697.710 ;
        RECT 204.715 1697.600 204.885 1697.760 ;
        RECT 204.715 1697.200 204.885 1697.430 ;
        RECT 207.435 1697.200 207.605 1697.285 ;
        RECT 210.155 1697.200 210.325 1697.285 ;
        RECT 201.995 1697.140 202.890 1697.200 ;
        RECT 202.165 1696.970 202.890 1697.140 ;
        RECT 201.995 1696.910 202.890 1696.970 ;
        RECT 203.550 1697.140 206.050 1697.200 ;
        RECT 203.550 1696.970 204.715 1697.140 ;
        RECT 204.885 1696.970 206.050 1697.140 ;
        RECT 203.550 1696.910 206.050 1696.970 ;
        RECT 206.710 1697.140 208.330 1697.200 ;
        RECT 206.710 1696.970 207.435 1697.140 ;
        RECT 207.605 1696.970 208.330 1697.140 ;
        RECT 206.710 1696.910 208.330 1696.970 ;
        RECT 208.990 1697.140 210.325 1697.200 ;
        RECT 208.990 1696.970 210.155 1697.140 ;
        RECT 208.990 1696.910 210.325 1696.970 ;
        RECT 201.995 1696.680 202.165 1696.910 ;
        RECT 204.715 1696.680 204.885 1696.910 ;
        RECT 207.435 1696.825 207.605 1696.910 ;
        RECT 210.155 1696.825 210.325 1696.910 ;
        RECT 201.995 1696.350 202.165 1696.510 ;
        RECT 204.715 1696.350 204.885 1696.510 ;
        RECT 205.055 1696.400 206.075 1696.730 ;
        RECT 201.995 1696.220 202.965 1696.350 ;
        RECT 202.165 1696.050 202.965 1696.220 ;
        RECT 201.995 1696.020 202.965 1696.050 ;
        RECT 203.565 1696.230 204.885 1696.350 ;
        RECT 203.565 1696.220 205.685 1696.230 ;
        RECT 203.565 1696.050 204.715 1696.220 ;
        RECT 204.885 1696.060 205.685 1696.220 ;
        RECT 203.565 1696.020 204.885 1696.050 ;
        RECT 201.995 1695.760 202.165 1696.020 ;
        RECT 204.715 1695.760 204.885 1696.020 ;
        RECT 205.905 1695.890 206.075 1696.400 ;
        RECT 201.995 1695.510 202.165 1695.590 ;
        RECT 204.715 1695.510 204.885 1695.590 ;
        RECT 205.055 1695.560 206.075 1695.890 ;
        RECT 201.995 1695.300 202.645 1695.510 ;
        RECT 203.915 1695.390 204.885 1695.510 ;
        RECT 205.905 1695.405 206.075 1695.560 ;
        RECT 206.615 1696.480 207.265 1696.650 ;
        RECT 206.615 1695.810 206.785 1696.480 ;
        RECT 206.955 1695.980 207.435 1696.310 ;
        RECT 206.615 1695.640 207.260 1695.810 ;
        RECT 206.615 1695.405 206.785 1695.640 ;
        RECT 202.165 1695.180 202.645 1695.300 ;
        RECT 201.995 1694.840 202.165 1695.130 ;
        RECT 201.995 1694.380 202.645 1694.670 ;
        RECT 202.165 1694.340 202.645 1694.380 ;
        RECT 201.995 1693.920 202.165 1694.210 ;
        RECT 202.165 1693.750 202.645 1693.830 ;
        RECT 201.995 1693.500 202.645 1693.750 ;
        RECT 201.995 1693.460 202.165 1693.500 ;
        RECT 201.995 1693.000 202.165 1693.290 ;
        RECT 202.165 1692.830 202.645 1692.990 ;
        RECT 203.155 1692.900 203.325 1695.350 ;
        RECT 203.915 1695.300 205.685 1695.390 ;
        RECT 203.915 1695.180 204.715 1695.300 ;
        RECT 204.885 1695.220 205.685 1695.300 ;
        RECT 205.905 1695.230 206.785 1695.405 ;
        RECT 204.715 1694.840 204.885 1695.130 ;
      LAYER li1 ;
        RECT 205.055 1694.800 206.075 1694.970 ;
      LAYER li1 ;
        RECT 203.915 1694.630 204.885 1694.670 ;
        RECT 203.915 1694.380 205.685 1694.630 ;
        RECT 203.915 1694.340 204.715 1694.380 ;
        RECT 204.885 1694.300 205.685 1694.380 ;
        RECT 204.715 1693.920 204.885 1694.210 ;
      LAYER li1 ;
        RECT 205.905 1694.130 206.075 1694.800 ;
        RECT 205.055 1693.960 206.075 1694.130 ;
      LAYER li1 ;
        RECT 203.915 1693.750 204.715 1693.830 ;
        RECT 204.885 1693.750 205.685 1693.790 ;
        RECT 203.915 1693.500 205.685 1693.750 ;
        RECT 204.715 1693.460 205.685 1693.500 ;
      LAYER li1 ;
        RECT 205.905 1693.290 206.075 1693.960 ;
      LAYER li1 ;
        RECT 204.715 1693.000 204.885 1693.290 ;
      LAYER li1 ;
        RECT 205.055 1693.120 206.075 1693.290 ;
      LAYER li1 ;
        RECT 201.995 1692.660 202.645 1692.830 ;
        RECT 202.815 1692.725 203.695 1692.900 ;
        RECT 203.915 1692.830 204.715 1692.910 ;
        RECT 204.885 1692.830 205.685 1692.950 ;
        RECT 203.915 1692.740 205.685 1692.830 ;
        RECT 201.995 1692.540 202.165 1692.660 ;
        RECT 202.815 1692.490 202.985 1692.725 ;
        RECT 203.525 1692.570 203.695 1692.725 ;
        RECT 204.715 1692.620 205.685 1692.740 ;
        RECT 201.995 1692.150 202.165 1692.370 ;
        RECT 202.340 1692.320 202.985 1692.490 ;
        RECT 201.995 1692.080 202.645 1692.150 ;
        RECT 202.165 1691.910 202.645 1692.080 ;
        RECT 201.995 1691.820 202.645 1691.910 ;
        RECT 201.995 1691.620 202.165 1691.820 ;
        RECT 202.815 1691.650 202.985 1692.320 ;
        RECT 202.335 1691.480 202.985 1691.650 ;
        RECT 201.995 1691.220 202.165 1691.450 ;
      LAYER li1 ;
        RECT 203.155 1691.445 203.355 1692.545 ;
      LAYER li1 ;
        RECT 203.525 1692.240 204.545 1692.570 ;
        RECT 204.715 1692.540 204.885 1692.620 ;
      LAYER li1 ;
        RECT 205.905 1692.535 206.075 1693.120 ;
      LAYER li1 ;
        RECT 206.275 1692.780 206.445 1695.230 ;
        RECT 206.955 1695.140 207.435 1695.470 ;
      LAYER li1 ;
        RECT 206.615 1694.800 207.265 1694.970 ;
        RECT 206.615 1694.130 206.785 1694.800 ;
      LAYER li1 ;
        RECT 206.955 1694.300 207.435 1694.630 ;
      LAYER li1 ;
        RECT 206.615 1693.960 207.265 1694.130 ;
        RECT 206.615 1693.290 206.785 1693.960 ;
      LAYER li1 ;
        RECT 206.955 1693.460 207.435 1693.790 ;
      LAYER li1 ;
        RECT 206.615 1693.120 207.265 1693.290 ;
        RECT 206.615 1692.535 206.785 1693.120 ;
      LAYER li1 ;
        RECT 206.955 1692.620 207.435 1692.950 ;
      LAYER li1 ;
        RECT 205.905 1692.450 206.785 1692.535 ;
      LAYER li1 ;
        RECT 203.525 1691.730 203.695 1692.240 ;
        RECT 204.715 1692.110 204.885 1692.370 ;
      LAYER li1 ;
        RECT 205.055 1692.280 207.265 1692.450 ;
      LAYER li1 ;
        RECT 204.715 1692.080 206.035 1692.110 ;
        RECT 203.915 1691.910 204.715 1692.070 ;
        RECT 204.885 1691.910 206.035 1692.080 ;
        RECT 203.915 1691.900 206.035 1691.910 ;
        RECT 204.715 1691.780 206.035 1691.900 ;
        RECT 206.635 1691.780 207.435 1692.110 ;
        RECT 203.525 1691.400 204.545 1691.730 ;
        RECT 204.715 1691.620 204.885 1691.780 ;
        RECT 204.715 1691.220 204.885 1691.450 ;
        RECT 207.435 1691.220 207.605 1691.305 ;
        RECT 210.155 1691.220 210.325 1691.305 ;
        RECT 201.995 1691.160 202.890 1691.220 ;
        RECT 202.165 1690.990 202.890 1691.160 ;
        RECT 201.995 1690.930 202.890 1690.990 ;
        RECT 203.550 1691.160 206.050 1691.220 ;
        RECT 203.550 1690.990 204.715 1691.160 ;
        RECT 204.885 1690.990 206.050 1691.160 ;
        RECT 203.550 1690.930 206.050 1690.990 ;
        RECT 206.710 1691.160 208.330 1691.220 ;
        RECT 206.710 1690.990 207.435 1691.160 ;
        RECT 207.605 1690.990 208.330 1691.160 ;
        RECT 206.710 1690.930 208.330 1690.990 ;
        RECT 208.990 1691.160 210.325 1691.220 ;
        RECT 208.990 1690.990 210.155 1691.160 ;
        RECT 208.990 1690.930 210.325 1690.990 ;
        RECT 201.995 1690.700 202.165 1690.930 ;
        RECT 204.715 1690.700 204.885 1690.930 ;
        RECT 207.435 1690.845 207.605 1690.930 ;
        RECT 210.155 1690.845 210.325 1690.930 ;
        RECT 201.995 1690.370 202.165 1690.530 ;
        RECT 204.715 1690.370 204.885 1690.530 ;
        RECT 205.055 1690.420 206.075 1690.750 ;
        RECT 201.995 1690.240 202.965 1690.370 ;
        RECT 202.165 1690.070 202.965 1690.240 ;
        RECT 201.995 1690.040 202.965 1690.070 ;
        RECT 203.565 1690.250 204.885 1690.370 ;
        RECT 203.565 1690.240 205.685 1690.250 ;
        RECT 203.565 1690.070 204.715 1690.240 ;
        RECT 204.885 1690.080 205.685 1690.240 ;
        RECT 203.565 1690.040 204.885 1690.070 ;
        RECT 201.995 1689.780 202.165 1690.040 ;
        RECT 204.715 1689.780 204.885 1690.040 ;
        RECT 205.905 1689.910 206.075 1690.420 ;
        RECT 201.995 1689.530 202.165 1689.610 ;
        RECT 204.715 1689.530 204.885 1689.610 ;
        RECT 205.055 1689.580 206.075 1689.910 ;
        RECT 201.995 1689.320 202.645 1689.530 ;
        RECT 203.915 1689.410 204.885 1689.530 ;
        RECT 205.905 1689.425 206.075 1689.580 ;
        RECT 206.615 1690.500 207.265 1690.670 ;
        RECT 206.615 1689.830 206.785 1690.500 ;
        RECT 206.955 1690.000 207.435 1690.330 ;
        RECT 206.615 1689.660 207.260 1689.830 ;
        RECT 206.615 1689.425 206.785 1689.660 ;
        RECT 202.165 1689.200 202.645 1689.320 ;
        RECT 201.995 1688.860 202.165 1689.150 ;
        RECT 201.995 1688.400 202.645 1688.690 ;
        RECT 202.165 1688.360 202.645 1688.400 ;
        RECT 201.995 1687.940 202.165 1688.230 ;
        RECT 202.165 1687.770 202.645 1687.850 ;
        RECT 201.995 1687.520 202.645 1687.770 ;
        RECT 201.995 1687.480 202.165 1687.520 ;
        RECT 201.995 1687.020 202.165 1687.310 ;
        RECT 202.165 1686.850 202.645 1687.010 ;
        RECT 203.155 1686.920 203.325 1689.370 ;
        RECT 203.915 1689.320 205.685 1689.410 ;
        RECT 203.915 1689.200 204.715 1689.320 ;
        RECT 204.885 1689.240 205.685 1689.320 ;
        RECT 205.905 1689.250 206.785 1689.425 ;
        RECT 204.715 1688.860 204.885 1689.150 ;
      LAYER li1 ;
        RECT 205.055 1688.820 206.075 1688.990 ;
      LAYER li1 ;
        RECT 203.915 1688.650 204.885 1688.690 ;
        RECT 203.915 1688.400 205.685 1688.650 ;
        RECT 203.915 1688.360 204.715 1688.400 ;
        RECT 204.885 1688.320 205.685 1688.400 ;
        RECT 204.715 1687.940 204.885 1688.230 ;
      LAYER li1 ;
        RECT 205.905 1688.150 206.075 1688.820 ;
        RECT 205.055 1687.980 206.075 1688.150 ;
      LAYER li1 ;
        RECT 203.915 1687.770 204.715 1687.850 ;
        RECT 204.885 1687.770 205.685 1687.810 ;
        RECT 203.915 1687.520 205.685 1687.770 ;
        RECT 204.715 1687.480 205.685 1687.520 ;
      LAYER li1 ;
        RECT 205.905 1687.310 206.075 1687.980 ;
      LAYER li1 ;
        RECT 204.715 1687.020 204.885 1687.310 ;
      LAYER li1 ;
        RECT 205.055 1687.140 206.075 1687.310 ;
      LAYER li1 ;
        RECT 201.995 1686.680 202.645 1686.850 ;
        RECT 202.815 1686.745 203.695 1686.920 ;
        RECT 203.915 1686.850 204.715 1686.930 ;
        RECT 204.885 1686.850 205.685 1686.970 ;
        RECT 203.915 1686.760 205.685 1686.850 ;
        RECT 201.995 1686.560 202.165 1686.680 ;
        RECT 202.815 1686.510 202.985 1686.745 ;
        RECT 203.525 1686.590 203.695 1686.745 ;
        RECT 204.715 1686.640 205.685 1686.760 ;
        RECT 201.995 1686.170 202.165 1686.390 ;
        RECT 202.340 1686.340 202.985 1686.510 ;
        RECT 201.995 1686.100 202.645 1686.170 ;
        RECT 202.165 1685.930 202.645 1686.100 ;
        RECT 201.995 1685.840 202.645 1685.930 ;
        RECT 201.995 1685.640 202.165 1685.840 ;
        RECT 202.815 1685.670 202.985 1686.340 ;
        RECT 202.335 1685.500 202.985 1685.670 ;
        RECT 201.995 1685.240 202.165 1685.470 ;
      LAYER li1 ;
        RECT 203.155 1685.465 203.355 1686.565 ;
      LAYER li1 ;
        RECT 203.525 1686.260 204.545 1686.590 ;
        RECT 204.715 1686.560 204.885 1686.640 ;
      LAYER li1 ;
        RECT 205.905 1686.555 206.075 1687.140 ;
      LAYER li1 ;
        RECT 206.275 1686.800 206.445 1689.250 ;
        RECT 206.955 1689.160 207.435 1689.490 ;
      LAYER li1 ;
        RECT 206.615 1688.820 207.265 1688.990 ;
        RECT 206.615 1688.150 206.785 1688.820 ;
      LAYER li1 ;
        RECT 206.955 1688.320 207.435 1688.650 ;
      LAYER li1 ;
        RECT 206.615 1687.980 207.265 1688.150 ;
        RECT 206.615 1687.310 206.785 1687.980 ;
      LAYER li1 ;
        RECT 206.955 1687.480 207.435 1687.810 ;
      LAYER li1 ;
        RECT 206.615 1687.140 207.265 1687.310 ;
        RECT 206.615 1686.555 206.785 1687.140 ;
      LAYER li1 ;
        RECT 206.955 1686.640 207.435 1686.970 ;
      LAYER li1 ;
        RECT 205.905 1686.470 206.785 1686.555 ;
      LAYER li1 ;
        RECT 203.525 1685.750 203.695 1686.260 ;
        RECT 204.715 1686.130 204.885 1686.390 ;
      LAYER li1 ;
        RECT 205.055 1686.300 207.265 1686.470 ;
      LAYER li1 ;
        RECT 204.715 1686.100 206.035 1686.130 ;
        RECT 203.915 1685.930 204.715 1686.090 ;
        RECT 204.885 1685.930 206.035 1686.100 ;
        RECT 203.915 1685.920 206.035 1685.930 ;
        RECT 204.715 1685.800 206.035 1685.920 ;
        RECT 206.635 1685.800 207.435 1686.130 ;
        RECT 203.525 1685.420 204.545 1685.750 ;
        RECT 204.715 1685.640 204.885 1685.800 ;
        RECT 204.715 1685.240 204.885 1685.470 ;
        RECT 207.435 1685.240 207.605 1685.325 ;
        RECT 210.155 1685.240 210.325 1685.325 ;
        RECT 201.995 1685.180 202.890 1685.240 ;
        RECT 202.165 1685.010 202.890 1685.180 ;
        RECT 201.995 1684.950 202.890 1685.010 ;
        RECT 203.550 1685.180 206.050 1685.240 ;
        RECT 203.550 1685.010 204.715 1685.180 ;
        RECT 204.885 1685.010 206.050 1685.180 ;
        RECT 203.550 1684.950 206.050 1685.010 ;
        RECT 206.710 1685.180 208.330 1685.240 ;
        RECT 206.710 1685.010 207.435 1685.180 ;
        RECT 207.605 1685.010 208.330 1685.180 ;
        RECT 206.710 1684.950 208.330 1685.010 ;
        RECT 208.990 1685.180 210.325 1685.240 ;
        RECT 208.990 1685.010 210.155 1685.180 ;
        RECT 208.990 1684.950 210.325 1685.010 ;
        RECT 201.995 1684.720 202.165 1684.950 ;
        RECT 204.715 1684.720 204.885 1684.950 ;
        RECT 207.435 1684.865 207.605 1684.950 ;
        RECT 210.155 1684.865 210.325 1684.950 ;
        RECT 201.995 1684.390 202.165 1684.550 ;
        RECT 204.715 1684.390 204.885 1684.550 ;
        RECT 205.055 1684.440 206.075 1684.770 ;
        RECT 201.995 1684.260 202.965 1684.390 ;
        RECT 202.165 1684.090 202.965 1684.260 ;
        RECT 201.995 1684.060 202.965 1684.090 ;
        RECT 203.565 1684.270 204.885 1684.390 ;
        RECT 203.565 1684.260 205.685 1684.270 ;
        RECT 203.565 1684.090 204.715 1684.260 ;
        RECT 204.885 1684.100 205.685 1684.260 ;
        RECT 203.565 1684.060 204.885 1684.090 ;
        RECT 201.995 1683.800 202.165 1684.060 ;
        RECT 204.715 1683.800 204.885 1684.060 ;
        RECT 205.905 1683.930 206.075 1684.440 ;
        RECT 201.995 1683.550 202.165 1683.630 ;
        RECT 204.715 1683.550 204.885 1683.630 ;
        RECT 205.055 1683.600 206.075 1683.930 ;
        RECT 201.995 1683.340 202.645 1683.550 ;
        RECT 203.915 1683.430 204.885 1683.550 ;
        RECT 205.905 1683.445 206.075 1683.600 ;
        RECT 206.615 1684.520 207.265 1684.690 ;
        RECT 206.615 1683.850 206.785 1684.520 ;
        RECT 206.955 1684.020 207.435 1684.350 ;
        RECT 206.615 1683.680 207.260 1683.850 ;
        RECT 206.615 1683.445 206.785 1683.680 ;
        RECT 202.165 1683.220 202.645 1683.340 ;
        RECT 201.995 1682.880 202.165 1683.170 ;
        RECT 201.995 1682.420 202.645 1682.710 ;
        RECT 202.165 1682.380 202.645 1682.420 ;
        RECT 201.995 1681.960 202.165 1682.250 ;
        RECT 202.165 1681.790 202.645 1681.870 ;
        RECT 201.995 1681.540 202.645 1681.790 ;
        RECT 201.995 1681.500 202.165 1681.540 ;
        RECT 201.995 1681.040 202.165 1681.330 ;
        RECT 202.165 1680.870 202.645 1681.030 ;
        RECT 203.155 1680.940 203.325 1683.390 ;
        RECT 203.915 1683.340 205.685 1683.430 ;
        RECT 203.915 1683.220 204.715 1683.340 ;
        RECT 204.885 1683.260 205.685 1683.340 ;
        RECT 205.905 1683.270 206.785 1683.445 ;
        RECT 204.715 1682.880 204.885 1683.170 ;
      LAYER li1 ;
        RECT 205.055 1682.840 206.075 1683.010 ;
      LAYER li1 ;
        RECT 203.915 1682.670 204.885 1682.710 ;
        RECT 203.915 1682.420 205.685 1682.670 ;
        RECT 203.915 1682.380 204.715 1682.420 ;
        RECT 204.885 1682.340 205.685 1682.420 ;
        RECT 204.715 1681.960 204.885 1682.250 ;
      LAYER li1 ;
        RECT 205.905 1682.170 206.075 1682.840 ;
        RECT 205.055 1682.000 206.075 1682.170 ;
      LAYER li1 ;
        RECT 203.915 1681.790 204.715 1681.870 ;
        RECT 204.885 1681.790 205.685 1681.830 ;
        RECT 203.915 1681.540 205.685 1681.790 ;
        RECT 204.715 1681.500 205.685 1681.540 ;
      LAYER li1 ;
        RECT 205.905 1681.330 206.075 1682.000 ;
      LAYER li1 ;
        RECT 204.715 1681.040 204.885 1681.330 ;
      LAYER li1 ;
        RECT 205.055 1681.160 206.075 1681.330 ;
      LAYER li1 ;
        RECT 201.995 1680.700 202.645 1680.870 ;
        RECT 202.815 1680.765 203.695 1680.940 ;
        RECT 203.915 1680.870 204.715 1680.950 ;
        RECT 204.885 1680.870 205.685 1680.990 ;
        RECT 203.915 1680.780 205.685 1680.870 ;
        RECT 201.995 1680.580 202.165 1680.700 ;
        RECT 202.815 1680.530 202.985 1680.765 ;
        RECT 203.525 1680.610 203.695 1680.765 ;
        RECT 204.715 1680.660 205.685 1680.780 ;
        RECT 201.995 1680.190 202.165 1680.410 ;
        RECT 202.340 1680.360 202.985 1680.530 ;
        RECT 201.995 1680.120 202.645 1680.190 ;
        RECT 202.165 1679.950 202.645 1680.120 ;
        RECT 201.995 1679.860 202.645 1679.950 ;
        RECT 201.995 1679.660 202.165 1679.860 ;
        RECT 202.815 1679.690 202.985 1680.360 ;
        RECT 202.335 1679.520 202.985 1679.690 ;
        RECT 201.995 1679.260 202.165 1679.490 ;
      LAYER li1 ;
        RECT 203.155 1679.485 203.355 1680.585 ;
      LAYER li1 ;
        RECT 203.525 1680.280 204.545 1680.610 ;
        RECT 204.715 1680.580 204.885 1680.660 ;
      LAYER li1 ;
        RECT 205.905 1680.575 206.075 1681.160 ;
      LAYER li1 ;
        RECT 206.275 1680.820 206.445 1683.270 ;
        RECT 206.955 1683.180 207.435 1683.510 ;
      LAYER li1 ;
        RECT 206.615 1682.840 207.265 1683.010 ;
        RECT 206.615 1682.170 206.785 1682.840 ;
      LAYER li1 ;
        RECT 206.955 1682.340 207.435 1682.670 ;
      LAYER li1 ;
        RECT 206.615 1682.000 207.265 1682.170 ;
        RECT 206.615 1681.330 206.785 1682.000 ;
      LAYER li1 ;
        RECT 206.955 1681.500 207.435 1681.830 ;
      LAYER li1 ;
        RECT 206.615 1681.160 207.265 1681.330 ;
        RECT 206.615 1680.575 206.785 1681.160 ;
      LAYER li1 ;
        RECT 206.955 1680.660 207.435 1680.990 ;
      LAYER li1 ;
        RECT 205.905 1680.490 206.785 1680.575 ;
      LAYER li1 ;
        RECT 203.525 1679.770 203.695 1680.280 ;
        RECT 204.715 1680.150 204.885 1680.410 ;
      LAYER li1 ;
        RECT 205.055 1680.320 207.265 1680.490 ;
      LAYER li1 ;
        RECT 204.715 1680.120 206.035 1680.150 ;
        RECT 203.915 1679.950 204.715 1680.110 ;
        RECT 204.885 1679.950 206.035 1680.120 ;
        RECT 203.915 1679.940 206.035 1679.950 ;
        RECT 204.715 1679.820 206.035 1679.940 ;
        RECT 206.635 1679.820 207.435 1680.150 ;
        RECT 203.525 1679.440 204.545 1679.770 ;
        RECT 204.715 1679.660 204.885 1679.820 ;
        RECT 204.715 1679.260 204.885 1679.490 ;
        RECT 207.435 1679.260 207.605 1679.345 ;
        RECT 210.155 1679.260 210.325 1679.345 ;
        RECT 201.995 1679.200 202.890 1679.260 ;
        RECT 202.165 1679.030 202.890 1679.200 ;
        RECT 201.995 1678.970 202.890 1679.030 ;
        RECT 203.550 1679.200 206.050 1679.260 ;
        RECT 203.550 1679.030 204.715 1679.200 ;
        RECT 204.885 1679.030 206.050 1679.200 ;
        RECT 203.550 1678.970 206.050 1679.030 ;
        RECT 206.710 1679.200 208.330 1679.260 ;
        RECT 206.710 1679.030 207.435 1679.200 ;
        RECT 207.605 1679.030 208.330 1679.200 ;
        RECT 206.710 1678.970 208.330 1679.030 ;
        RECT 208.990 1679.200 210.325 1679.260 ;
        RECT 208.990 1679.030 210.155 1679.200 ;
        RECT 208.990 1678.970 210.325 1679.030 ;
        RECT 201.995 1678.740 202.165 1678.970 ;
        RECT 204.715 1678.740 204.885 1678.970 ;
        RECT 207.435 1678.885 207.605 1678.970 ;
        RECT 210.155 1678.885 210.325 1678.970 ;
        RECT 201.995 1678.410 202.165 1678.570 ;
        RECT 204.715 1678.410 204.885 1678.570 ;
        RECT 205.055 1678.460 206.075 1678.790 ;
        RECT 201.995 1678.280 202.965 1678.410 ;
        RECT 202.165 1678.110 202.965 1678.280 ;
        RECT 201.995 1678.080 202.965 1678.110 ;
        RECT 203.565 1678.290 204.885 1678.410 ;
        RECT 203.565 1678.280 205.685 1678.290 ;
        RECT 203.565 1678.110 204.715 1678.280 ;
        RECT 204.885 1678.120 205.685 1678.280 ;
        RECT 203.565 1678.080 204.885 1678.110 ;
        RECT 201.995 1677.820 202.165 1678.080 ;
        RECT 204.715 1677.820 204.885 1678.080 ;
        RECT 205.905 1677.950 206.075 1678.460 ;
        RECT 201.995 1677.570 202.165 1677.650 ;
        RECT 204.715 1677.570 204.885 1677.650 ;
        RECT 205.055 1677.620 206.075 1677.950 ;
        RECT 201.995 1677.360 202.645 1677.570 ;
        RECT 203.915 1677.450 204.885 1677.570 ;
        RECT 205.905 1677.465 206.075 1677.620 ;
        RECT 206.615 1678.540 207.265 1678.710 ;
        RECT 206.615 1677.870 206.785 1678.540 ;
        RECT 206.955 1678.040 207.435 1678.370 ;
        RECT 206.615 1677.700 207.260 1677.870 ;
        RECT 206.615 1677.465 206.785 1677.700 ;
        RECT 202.165 1677.240 202.645 1677.360 ;
        RECT 201.995 1676.900 202.165 1677.190 ;
        RECT 201.995 1676.440 202.645 1676.730 ;
        RECT 202.165 1676.400 202.645 1676.440 ;
        RECT 201.995 1675.980 202.165 1676.270 ;
        RECT 202.165 1675.810 202.645 1675.890 ;
        RECT 201.995 1675.560 202.645 1675.810 ;
        RECT 201.995 1675.520 202.165 1675.560 ;
        RECT 201.995 1675.060 202.165 1675.350 ;
        RECT 202.165 1674.890 202.645 1675.050 ;
        RECT 203.155 1674.960 203.325 1677.410 ;
        RECT 203.915 1677.360 205.685 1677.450 ;
        RECT 203.915 1677.240 204.715 1677.360 ;
        RECT 204.885 1677.280 205.685 1677.360 ;
        RECT 205.905 1677.290 206.785 1677.465 ;
        RECT 204.715 1676.900 204.885 1677.190 ;
      LAYER li1 ;
        RECT 205.055 1676.860 206.075 1677.030 ;
      LAYER li1 ;
        RECT 203.915 1676.690 204.885 1676.730 ;
        RECT 203.915 1676.440 205.685 1676.690 ;
        RECT 203.915 1676.400 204.715 1676.440 ;
        RECT 204.885 1676.360 205.685 1676.440 ;
        RECT 204.715 1675.980 204.885 1676.270 ;
      LAYER li1 ;
        RECT 205.905 1676.190 206.075 1676.860 ;
        RECT 205.055 1676.020 206.075 1676.190 ;
      LAYER li1 ;
        RECT 203.915 1675.810 204.715 1675.890 ;
        RECT 204.885 1675.810 205.685 1675.850 ;
        RECT 203.915 1675.560 205.685 1675.810 ;
        RECT 204.715 1675.520 205.685 1675.560 ;
      LAYER li1 ;
        RECT 205.905 1675.350 206.075 1676.020 ;
      LAYER li1 ;
        RECT 204.715 1675.060 204.885 1675.350 ;
      LAYER li1 ;
        RECT 205.055 1675.180 206.075 1675.350 ;
      LAYER li1 ;
        RECT 201.995 1674.720 202.645 1674.890 ;
        RECT 202.815 1674.785 203.695 1674.960 ;
        RECT 203.915 1674.890 204.715 1674.970 ;
        RECT 204.885 1674.890 205.685 1675.010 ;
        RECT 203.915 1674.800 205.685 1674.890 ;
        RECT 201.995 1674.600 202.165 1674.720 ;
        RECT 202.815 1674.550 202.985 1674.785 ;
        RECT 203.525 1674.630 203.695 1674.785 ;
        RECT 204.715 1674.680 205.685 1674.800 ;
        RECT 201.995 1674.210 202.165 1674.430 ;
        RECT 202.340 1674.380 202.985 1674.550 ;
        RECT 201.995 1674.140 202.645 1674.210 ;
        RECT 202.165 1673.970 202.645 1674.140 ;
        RECT 201.995 1673.880 202.645 1673.970 ;
        RECT 201.995 1673.680 202.165 1673.880 ;
        RECT 202.815 1673.710 202.985 1674.380 ;
        RECT 202.335 1673.540 202.985 1673.710 ;
        RECT 201.995 1673.280 202.165 1673.510 ;
      LAYER li1 ;
        RECT 203.155 1673.505 203.355 1674.605 ;
      LAYER li1 ;
        RECT 203.525 1674.300 204.545 1674.630 ;
        RECT 204.715 1674.600 204.885 1674.680 ;
      LAYER li1 ;
        RECT 205.905 1674.595 206.075 1675.180 ;
      LAYER li1 ;
        RECT 206.275 1674.840 206.445 1677.290 ;
        RECT 206.955 1677.200 207.435 1677.530 ;
      LAYER li1 ;
        RECT 206.615 1676.860 207.265 1677.030 ;
        RECT 206.615 1676.190 206.785 1676.860 ;
      LAYER li1 ;
        RECT 206.955 1676.360 207.435 1676.690 ;
      LAYER li1 ;
        RECT 206.615 1676.020 207.265 1676.190 ;
        RECT 206.615 1675.350 206.785 1676.020 ;
      LAYER li1 ;
        RECT 206.955 1675.520 207.435 1675.850 ;
      LAYER li1 ;
        RECT 206.615 1675.180 207.265 1675.350 ;
        RECT 206.615 1674.595 206.785 1675.180 ;
      LAYER li1 ;
        RECT 206.955 1674.680 207.435 1675.010 ;
      LAYER li1 ;
        RECT 205.905 1674.510 206.785 1674.595 ;
      LAYER li1 ;
        RECT 203.525 1673.790 203.695 1674.300 ;
        RECT 204.715 1674.170 204.885 1674.430 ;
      LAYER li1 ;
        RECT 205.055 1674.340 207.265 1674.510 ;
      LAYER li1 ;
        RECT 204.715 1674.140 206.035 1674.170 ;
        RECT 203.915 1673.970 204.715 1674.130 ;
        RECT 204.885 1673.970 206.035 1674.140 ;
        RECT 203.915 1673.960 206.035 1673.970 ;
        RECT 204.715 1673.840 206.035 1673.960 ;
        RECT 206.635 1673.840 207.435 1674.170 ;
        RECT 203.525 1673.460 204.545 1673.790 ;
        RECT 204.715 1673.680 204.885 1673.840 ;
        RECT 204.715 1673.280 204.885 1673.510 ;
        RECT 207.435 1673.280 207.605 1673.365 ;
        RECT 210.155 1673.280 210.325 1673.365 ;
        RECT 201.995 1673.220 202.890 1673.280 ;
        RECT 202.165 1673.050 202.890 1673.220 ;
        RECT 201.995 1672.990 202.890 1673.050 ;
        RECT 203.550 1673.220 206.050 1673.280 ;
        RECT 203.550 1673.050 204.715 1673.220 ;
        RECT 204.885 1673.050 206.050 1673.220 ;
        RECT 203.550 1672.990 206.050 1673.050 ;
        RECT 206.710 1673.220 208.330 1673.280 ;
        RECT 206.710 1673.050 207.435 1673.220 ;
        RECT 207.605 1673.050 208.330 1673.220 ;
        RECT 206.710 1672.990 208.330 1673.050 ;
        RECT 208.990 1673.220 210.325 1673.280 ;
        RECT 208.990 1673.050 210.155 1673.220 ;
        RECT 208.990 1672.990 210.325 1673.050 ;
        RECT 201.995 1672.905 202.165 1672.990 ;
        RECT 204.715 1672.905 204.885 1672.990 ;
        RECT 207.435 1672.905 207.605 1672.990 ;
        RECT 210.155 1672.905 210.325 1672.990 ;
        RECT 669.000 219.760 669.145 219.930 ;
        RECT 669.315 219.760 669.460 219.930 ;
        RECT 674.980 219.760 675.125 219.930 ;
        RECT 675.295 219.760 675.440 219.930 ;
        RECT 680.960 219.760 681.105 219.930 ;
        RECT 681.275 219.760 681.420 219.930 ;
        RECT 686.940 219.760 687.085 219.930 ;
        RECT 687.255 219.760 687.400 219.930 ;
        RECT 692.920 219.760 693.065 219.930 ;
        RECT 693.235 219.760 693.380 219.930 ;
        RECT 698.900 219.760 699.045 219.930 ;
        RECT 699.215 219.760 699.360 219.930 ;
        RECT 704.880 219.760 705.025 219.930 ;
        RECT 705.195 219.760 705.340 219.930 ;
        RECT 710.860 219.760 711.005 219.930 ;
        RECT 711.175 219.760 711.320 219.930 ;
        RECT 716.840 219.760 716.985 219.930 ;
        RECT 717.155 219.760 717.300 219.930 ;
        RECT 722.820 219.760 722.965 219.930 ;
        RECT 723.135 219.760 723.280 219.930 ;
        RECT 728.800 219.760 728.945 219.930 ;
        RECT 729.115 219.760 729.260 219.930 ;
        RECT 734.780 219.760 734.925 219.930 ;
        RECT 735.095 219.760 735.240 219.930 ;
        RECT 740.760 219.760 740.905 219.930 ;
        RECT 741.075 219.760 741.220 219.930 ;
        RECT 746.740 219.760 746.885 219.930 ;
        RECT 747.055 219.760 747.200 219.930 ;
        RECT 752.720 219.760 752.865 219.930 ;
        RECT 753.035 219.760 753.180 219.930 ;
        RECT 758.700 219.760 758.845 219.930 ;
        RECT 759.015 219.760 759.160 219.930 ;
        RECT 764.680 219.760 764.825 219.930 ;
        RECT 764.995 219.760 765.140 219.930 ;
        RECT 770.660 219.760 770.805 219.930 ;
        RECT 770.975 219.760 771.120 219.930 ;
        RECT 776.640 219.760 776.785 219.930 ;
        RECT 776.955 219.760 777.100 219.930 ;
        RECT 782.620 219.760 782.765 219.930 ;
        RECT 782.935 219.760 783.080 219.930 ;
        RECT 788.600 219.760 788.745 219.930 ;
        RECT 788.915 219.760 789.060 219.930 ;
        RECT 794.580 219.760 794.725 219.930 ;
        RECT 794.895 219.760 795.040 219.930 ;
        RECT 2146.000 219.760 2146.145 219.930 ;
        RECT 2146.315 219.760 2146.460 219.930 ;
        RECT 2151.980 219.760 2152.125 219.930 ;
        RECT 2152.295 219.760 2152.440 219.930 ;
        RECT 2157.960 219.760 2158.105 219.930 ;
        RECT 2158.275 219.760 2158.420 219.930 ;
        RECT 2163.940 219.760 2164.085 219.930 ;
        RECT 2164.255 219.760 2164.400 219.930 ;
        RECT 2169.920 219.760 2170.065 219.930 ;
        RECT 2170.235 219.760 2170.380 219.930 ;
        RECT 2175.900 219.760 2176.045 219.930 ;
        RECT 2176.215 219.760 2176.360 219.930 ;
        RECT 2181.880 219.760 2182.025 219.930 ;
        RECT 2182.195 219.760 2182.340 219.930 ;
        RECT 2187.860 219.760 2188.005 219.930 ;
        RECT 2188.175 219.760 2188.320 219.930 ;
        RECT 2193.840 219.760 2193.985 219.930 ;
        RECT 2194.155 219.760 2194.300 219.930 ;
        RECT 2199.820 219.760 2199.965 219.930 ;
        RECT 2200.135 219.760 2200.280 219.930 ;
        RECT 2205.800 219.760 2205.945 219.930 ;
        RECT 2206.115 219.760 2206.260 219.930 ;
        RECT 2211.780 219.760 2211.925 219.930 ;
        RECT 2212.095 219.760 2212.240 219.930 ;
        RECT 2217.760 219.760 2217.905 219.930 ;
        RECT 2218.075 219.760 2218.220 219.930 ;
        RECT 2223.740 219.760 2223.885 219.930 ;
        RECT 2224.055 219.760 2224.200 219.930 ;
        RECT 2229.720 219.760 2229.865 219.930 ;
        RECT 2230.035 219.760 2230.180 219.930 ;
        RECT 2235.700 219.760 2235.845 219.930 ;
        RECT 2236.015 219.760 2236.160 219.930 ;
        RECT 2241.680 219.760 2241.825 219.930 ;
        RECT 2241.995 219.760 2242.140 219.930 ;
        RECT 2247.660 219.760 2247.805 219.930 ;
        RECT 2247.975 219.760 2248.120 219.930 ;
        RECT 2253.640 219.760 2253.785 219.930 ;
        RECT 2253.955 219.760 2254.100 219.930 ;
        RECT 2259.620 219.760 2259.765 219.930 ;
        RECT 2259.935 219.760 2260.080 219.930 ;
        RECT 2265.600 219.760 2265.745 219.930 ;
        RECT 2265.915 219.760 2266.060 219.930 ;
        RECT 2271.580 219.760 2271.725 219.930 ;
        RECT 2271.895 219.760 2272.040 219.930 ;
        RECT 669.085 218.595 669.375 219.760 ;
        RECT 675.065 218.595 675.355 219.760 ;
        RECT 681.045 218.595 681.335 219.760 ;
        RECT 687.025 218.595 687.315 219.760 ;
        RECT 693.005 218.595 693.295 219.760 ;
        RECT 698.985 218.595 699.275 219.760 ;
        RECT 704.965 218.595 705.255 219.760 ;
        RECT 710.945 218.595 711.235 219.760 ;
        RECT 716.925 218.595 717.215 219.760 ;
        RECT 722.905 218.595 723.195 219.760 ;
        RECT 728.885 218.595 729.175 219.760 ;
        RECT 734.865 218.595 735.155 219.760 ;
        RECT 740.845 218.595 741.135 219.760 ;
        RECT 746.825 218.595 747.115 219.760 ;
        RECT 752.805 218.595 753.095 219.760 ;
        RECT 758.785 218.595 759.075 219.760 ;
        RECT 764.765 218.595 765.055 219.760 ;
        RECT 770.745 218.595 771.035 219.760 ;
        RECT 776.725 218.595 777.015 219.760 ;
        RECT 782.705 218.595 782.995 219.760 ;
        RECT 788.685 218.595 788.975 219.760 ;
        RECT 794.665 218.595 794.955 219.760 ;
        RECT 2146.085 218.595 2146.375 219.760 ;
        RECT 2152.065 218.595 2152.355 219.760 ;
        RECT 2158.045 218.595 2158.335 219.760 ;
        RECT 2164.025 218.595 2164.315 219.760 ;
        RECT 2170.005 218.595 2170.295 219.760 ;
        RECT 2175.985 218.595 2176.275 219.760 ;
        RECT 2181.965 218.595 2182.255 219.760 ;
        RECT 2187.945 218.595 2188.235 219.760 ;
        RECT 2193.925 218.595 2194.215 219.760 ;
        RECT 2199.905 218.595 2200.195 219.760 ;
        RECT 2205.885 218.595 2206.175 219.760 ;
        RECT 2211.865 218.595 2212.155 219.760 ;
        RECT 2217.845 218.595 2218.135 219.760 ;
        RECT 2223.825 218.595 2224.115 219.760 ;
        RECT 2229.805 218.595 2230.095 219.760 ;
        RECT 2235.785 218.595 2236.075 219.760 ;
        RECT 2241.765 218.595 2242.055 219.760 ;
        RECT 2247.745 218.595 2248.035 219.760 ;
        RECT 2253.725 218.595 2254.015 219.760 ;
        RECT 2259.705 218.595 2259.995 219.760 ;
        RECT 2265.685 218.595 2265.975 219.760 ;
        RECT 2271.665 218.595 2271.955 219.760 ;
        RECT 669.085 217.210 669.375 217.935 ;
      LAYER li1 ;
        RECT 671.130 217.755 671.470 218.585 ;
        RECT 669.545 217.210 674.890 217.755 ;
      LAYER li1 ;
        RECT 675.065 217.210 675.355 217.935 ;
        RECT 681.045 217.210 681.335 217.935 ;
        RECT 687.025 217.210 687.315 217.935 ;
        RECT 693.005 217.210 693.295 217.935 ;
        RECT 698.985 217.210 699.275 217.935 ;
        RECT 704.965 217.210 705.255 217.935 ;
        RECT 710.945 217.210 711.235 217.935 ;
        RECT 716.925 217.210 717.215 217.935 ;
        RECT 722.905 217.210 723.195 217.935 ;
        RECT 728.885 217.210 729.175 217.935 ;
        RECT 734.865 217.210 735.155 217.935 ;
        RECT 740.845 217.210 741.135 217.935 ;
        RECT 746.825 217.210 747.115 217.935 ;
        RECT 752.805 217.210 753.095 217.935 ;
        RECT 758.785 217.210 759.075 217.935 ;
        RECT 764.765 217.210 765.055 217.935 ;
        RECT 770.745 217.210 771.035 217.935 ;
        RECT 776.725 217.210 777.015 217.935 ;
        RECT 782.705 217.210 782.995 217.935 ;
        RECT 788.685 217.210 788.975 217.935 ;
        RECT 794.665 217.210 794.955 217.935 ;
        RECT 2146.085 217.210 2146.375 217.935 ;
        RECT 2152.065 217.210 2152.355 217.935 ;
        RECT 2158.045 217.210 2158.335 217.935 ;
        RECT 2164.025 217.210 2164.315 217.935 ;
        RECT 2170.005 217.210 2170.295 217.935 ;
        RECT 2175.985 217.210 2176.275 217.935 ;
        RECT 2181.965 217.210 2182.255 217.935 ;
        RECT 2187.945 217.210 2188.235 217.935 ;
        RECT 2193.925 217.210 2194.215 217.935 ;
        RECT 2199.905 217.210 2200.195 217.935 ;
        RECT 2205.885 217.210 2206.175 217.935 ;
        RECT 2211.865 217.210 2212.155 217.935 ;
        RECT 2217.845 217.210 2218.135 217.935 ;
        RECT 2223.825 217.210 2224.115 217.935 ;
        RECT 2229.805 217.210 2230.095 217.935 ;
        RECT 2235.785 217.210 2236.075 217.935 ;
      LAYER li1 ;
        RECT 2237.830 217.755 2238.170 218.585 ;
        RECT 2236.245 217.210 2241.590 217.755 ;
      LAYER li1 ;
        RECT 2241.765 217.210 2242.055 217.935 ;
      LAYER li1 ;
        RECT 2243.810 217.755 2244.150 218.585 ;
        RECT 2242.225 217.210 2247.570 217.755 ;
      LAYER li1 ;
        RECT 2247.745 217.210 2248.035 217.935 ;
      LAYER li1 ;
        RECT 2249.790 217.755 2250.130 218.585 ;
        RECT 2248.205 217.210 2253.550 217.755 ;
      LAYER li1 ;
        RECT 2253.725 217.210 2254.015 217.935 ;
      LAYER li1 ;
        RECT 2255.770 217.755 2256.110 218.585 ;
        RECT 2254.185 217.210 2259.530 217.755 ;
      LAYER li1 ;
        RECT 2259.705 217.210 2259.995 217.935 ;
      LAYER li1 ;
        RECT 2261.750 217.755 2262.090 218.585 ;
        RECT 2260.165 217.210 2265.510 217.755 ;
      LAYER li1 ;
        RECT 2265.685 217.210 2265.975 217.935 ;
      LAYER li1 ;
        RECT 2267.730 217.755 2268.070 218.585 ;
        RECT 2266.145 217.210 2271.490 217.755 ;
      LAYER li1 ;
        RECT 2271.665 217.210 2271.955 217.935 ;
        RECT 669.000 217.040 669.145 217.210 ;
        RECT 669.315 217.040 669.605 217.210 ;
        RECT 669.775 217.040 670.065 217.210 ;
        RECT 670.235 217.040 670.525 217.210 ;
        RECT 670.695 217.040 670.985 217.210 ;
        RECT 671.155 217.040 671.445 217.210 ;
        RECT 671.615 217.040 671.905 217.210 ;
        RECT 672.075 217.040 672.365 217.210 ;
        RECT 672.535 217.040 672.825 217.210 ;
        RECT 672.995 217.040 673.285 217.210 ;
        RECT 673.455 217.040 673.745 217.210 ;
        RECT 673.915 217.040 674.205 217.210 ;
        RECT 674.375 217.040 674.665 217.210 ;
        RECT 674.835 217.040 675.125 217.210 ;
        RECT 675.295 217.040 675.440 217.210 ;
        RECT 680.960 217.040 681.105 217.210 ;
        RECT 681.275 217.040 681.420 217.210 ;
        RECT 686.940 217.040 687.085 217.210 ;
        RECT 687.255 217.040 687.400 217.210 ;
        RECT 692.920 217.040 693.065 217.210 ;
        RECT 693.235 217.040 693.380 217.210 ;
        RECT 698.900 217.040 699.045 217.210 ;
        RECT 699.215 217.040 699.360 217.210 ;
        RECT 704.880 217.040 705.025 217.210 ;
        RECT 705.195 217.040 705.340 217.210 ;
        RECT 710.860 217.040 711.005 217.210 ;
        RECT 711.175 217.040 711.320 217.210 ;
        RECT 716.840 217.040 716.985 217.210 ;
        RECT 717.155 217.040 717.300 217.210 ;
        RECT 722.820 217.040 722.965 217.210 ;
        RECT 723.135 217.040 723.280 217.210 ;
        RECT 728.800 217.040 728.945 217.210 ;
        RECT 729.115 217.040 729.260 217.210 ;
        RECT 734.780 217.040 734.925 217.210 ;
        RECT 735.095 217.040 735.240 217.210 ;
        RECT 740.760 217.040 740.905 217.210 ;
        RECT 741.075 217.040 741.220 217.210 ;
        RECT 746.740 217.040 746.885 217.210 ;
        RECT 747.055 217.040 747.200 217.210 ;
        RECT 752.720 217.040 752.865 217.210 ;
        RECT 753.035 217.040 753.180 217.210 ;
        RECT 758.700 217.040 758.845 217.210 ;
        RECT 759.015 217.040 759.160 217.210 ;
        RECT 764.680 217.040 764.825 217.210 ;
        RECT 764.995 217.040 765.140 217.210 ;
        RECT 770.660 217.040 770.805 217.210 ;
        RECT 770.975 217.040 771.120 217.210 ;
        RECT 776.640 217.040 776.785 217.210 ;
        RECT 776.955 217.040 777.100 217.210 ;
        RECT 782.620 217.040 782.765 217.210 ;
        RECT 782.935 217.040 783.080 217.210 ;
        RECT 788.600 217.040 788.745 217.210 ;
        RECT 788.915 217.040 789.060 217.210 ;
        RECT 794.580 217.040 794.725 217.210 ;
        RECT 794.895 217.040 795.040 217.210 ;
        RECT 2146.000 217.040 2146.145 217.210 ;
        RECT 2146.315 217.040 2146.460 217.210 ;
        RECT 2151.980 217.040 2152.125 217.210 ;
        RECT 2152.295 217.040 2152.440 217.210 ;
        RECT 2157.960 217.040 2158.105 217.210 ;
        RECT 2158.275 217.040 2158.420 217.210 ;
        RECT 2163.940 217.040 2164.085 217.210 ;
        RECT 2164.255 217.040 2164.400 217.210 ;
        RECT 2169.920 217.040 2170.065 217.210 ;
        RECT 2170.235 217.040 2170.380 217.210 ;
        RECT 2175.900 217.040 2176.045 217.210 ;
        RECT 2176.215 217.040 2176.360 217.210 ;
        RECT 2181.880 217.040 2182.025 217.210 ;
        RECT 2182.195 217.040 2182.340 217.210 ;
        RECT 2187.860 217.040 2188.005 217.210 ;
        RECT 2188.175 217.040 2188.320 217.210 ;
        RECT 2193.840 217.040 2193.985 217.210 ;
        RECT 2194.155 217.040 2194.300 217.210 ;
        RECT 2199.820 217.040 2199.965 217.210 ;
        RECT 2200.135 217.040 2200.280 217.210 ;
        RECT 2205.800 217.040 2205.945 217.210 ;
        RECT 2206.115 217.040 2206.260 217.210 ;
        RECT 2211.780 217.040 2211.925 217.210 ;
        RECT 2212.095 217.040 2212.240 217.210 ;
        RECT 2217.760 217.040 2217.905 217.210 ;
        RECT 2218.075 217.040 2218.220 217.210 ;
        RECT 2223.740 217.040 2223.885 217.210 ;
        RECT 2224.055 217.040 2224.200 217.210 ;
        RECT 2229.720 217.040 2229.865 217.210 ;
        RECT 2230.035 217.040 2230.180 217.210 ;
        RECT 2235.700 217.040 2235.845 217.210 ;
        RECT 2236.015 217.040 2236.305 217.210 ;
        RECT 2236.475 217.040 2236.765 217.210 ;
        RECT 2236.935 217.040 2237.225 217.210 ;
        RECT 2237.395 217.040 2237.685 217.210 ;
        RECT 2237.855 217.040 2238.145 217.210 ;
        RECT 2238.315 217.040 2238.605 217.210 ;
        RECT 2238.775 217.040 2239.065 217.210 ;
        RECT 2239.235 217.040 2239.525 217.210 ;
        RECT 2239.695 217.040 2239.985 217.210 ;
        RECT 2240.155 217.040 2240.445 217.210 ;
        RECT 2240.615 217.040 2240.905 217.210 ;
        RECT 2241.075 217.040 2241.365 217.210 ;
        RECT 2241.535 217.040 2241.825 217.210 ;
        RECT 2241.995 217.040 2242.285 217.210 ;
        RECT 2242.455 217.040 2242.745 217.210 ;
        RECT 2242.915 217.040 2243.205 217.210 ;
        RECT 2243.375 217.040 2243.665 217.210 ;
        RECT 2243.835 217.040 2244.125 217.210 ;
        RECT 2244.295 217.040 2244.585 217.210 ;
        RECT 2244.755 217.040 2245.045 217.210 ;
        RECT 2245.215 217.040 2245.505 217.210 ;
        RECT 2245.675 217.040 2245.965 217.210 ;
        RECT 2246.135 217.040 2246.425 217.210 ;
        RECT 2246.595 217.040 2246.885 217.210 ;
        RECT 2247.055 217.040 2247.345 217.210 ;
        RECT 2247.515 217.040 2247.805 217.210 ;
        RECT 2247.975 217.040 2248.265 217.210 ;
        RECT 2248.435 217.040 2248.725 217.210 ;
        RECT 2248.895 217.040 2249.185 217.210 ;
        RECT 2249.355 217.040 2249.645 217.210 ;
        RECT 2249.815 217.040 2250.105 217.210 ;
        RECT 2250.275 217.040 2250.565 217.210 ;
        RECT 2250.735 217.040 2251.025 217.210 ;
        RECT 2251.195 217.040 2251.485 217.210 ;
        RECT 2251.655 217.040 2251.945 217.210 ;
        RECT 2252.115 217.040 2252.405 217.210 ;
        RECT 2252.575 217.040 2252.865 217.210 ;
        RECT 2253.035 217.040 2253.325 217.210 ;
        RECT 2253.495 217.040 2253.785 217.210 ;
        RECT 2253.955 217.040 2254.245 217.210 ;
        RECT 2254.415 217.040 2254.705 217.210 ;
        RECT 2254.875 217.040 2255.165 217.210 ;
        RECT 2255.335 217.040 2255.625 217.210 ;
        RECT 2255.795 217.040 2256.085 217.210 ;
        RECT 2256.255 217.040 2256.545 217.210 ;
        RECT 2256.715 217.040 2257.005 217.210 ;
        RECT 2257.175 217.040 2257.465 217.210 ;
        RECT 2257.635 217.040 2257.925 217.210 ;
        RECT 2258.095 217.040 2258.385 217.210 ;
        RECT 2258.555 217.040 2258.845 217.210 ;
        RECT 2259.015 217.040 2259.305 217.210 ;
        RECT 2259.475 217.040 2259.765 217.210 ;
        RECT 2259.935 217.040 2260.225 217.210 ;
        RECT 2260.395 217.040 2260.685 217.210 ;
        RECT 2260.855 217.040 2261.145 217.210 ;
        RECT 2261.315 217.040 2261.605 217.210 ;
        RECT 2261.775 217.040 2262.065 217.210 ;
        RECT 2262.235 217.040 2262.525 217.210 ;
        RECT 2262.695 217.040 2262.985 217.210 ;
        RECT 2263.155 217.040 2263.445 217.210 ;
        RECT 2263.615 217.040 2263.905 217.210 ;
        RECT 2264.075 217.040 2264.365 217.210 ;
        RECT 2264.535 217.040 2264.825 217.210 ;
        RECT 2264.995 217.040 2265.285 217.210 ;
        RECT 2265.455 217.040 2265.745 217.210 ;
        RECT 2265.915 217.040 2266.205 217.210 ;
        RECT 2266.375 217.040 2266.665 217.210 ;
        RECT 2266.835 217.040 2267.125 217.210 ;
        RECT 2267.295 217.040 2267.585 217.210 ;
        RECT 2267.755 217.040 2268.045 217.210 ;
        RECT 2268.215 217.040 2268.505 217.210 ;
        RECT 2268.675 217.040 2268.965 217.210 ;
        RECT 2269.135 217.040 2269.425 217.210 ;
        RECT 2269.595 217.040 2269.885 217.210 ;
        RECT 2270.055 217.040 2270.345 217.210 ;
        RECT 2270.515 217.040 2270.805 217.210 ;
        RECT 2270.975 217.040 2271.265 217.210 ;
        RECT 2271.435 217.040 2271.725 217.210 ;
        RECT 2271.895 217.040 2272.040 217.210 ;
        RECT 669.085 216.315 669.375 217.040 ;
        RECT 669.935 216.240 670.265 217.040 ;
      LAYER li1 ;
        RECT 670.435 216.390 670.605 216.870 ;
      LAYER li1 ;
        RECT 670.775 216.560 671.105 217.040 ;
      LAYER li1 ;
        RECT 671.275 216.390 671.445 216.870 ;
      LAYER li1 ;
        RECT 671.615 216.560 671.945 217.040 ;
      LAYER li1 ;
        RECT 672.115 216.390 672.285 216.870 ;
      LAYER li1 ;
        RECT 672.455 216.560 672.785 217.040 ;
      LAYER li1 ;
        RECT 672.955 216.390 673.125 216.870 ;
      LAYER li1 ;
        RECT 673.295 216.560 673.625 217.040 ;
        RECT 673.795 216.390 673.965 216.865 ;
        RECT 674.135 216.560 674.465 217.040 ;
        RECT 674.635 216.390 674.805 216.870 ;
      LAYER li1 ;
        RECT 670.435 216.220 673.125 216.390 ;
      LAYER li1 ;
        RECT 673.385 216.220 674.805 216.390 ;
        RECT 675.065 216.315 675.355 217.040 ;
        RECT 675.915 216.240 676.245 217.040 ;
      LAYER li1 ;
        RECT 676.415 216.390 676.585 216.870 ;
      LAYER li1 ;
        RECT 676.755 216.560 677.085 217.040 ;
      LAYER li1 ;
        RECT 677.255 216.390 677.425 216.870 ;
      LAYER li1 ;
        RECT 677.595 216.560 677.925 217.040 ;
      LAYER li1 ;
        RECT 678.095 216.390 678.265 216.870 ;
      LAYER li1 ;
        RECT 678.435 216.560 678.765 217.040 ;
      LAYER li1 ;
        RECT 678.935 216.390 679.105 216.870 ;
      LAYER li1 ;
        RECT 679.275 216.560 679.605 217.040 ;
        RECT 679.775 216.390 679.945 216.865 ;
        RECT 680.115 216.560 680.445 217.040 ;
        RECT 680.615 216.390 680.785 216.870 ;
      LAYER li1 ;
        RECT 676.415 216.220 679.105 216.390 ;
      LAYER li1 ;
        RECT 679.365 216.220 680.785 216.390 ;
        RECT 681.045 216.315 681.335 217.040 ;
        RECT 681.895 216.240 682.225 217.040 ;
      LAYER li1 ;
        RECT 682.395 216.390 682.565 216.870 ;
      LAYER li1 ;
        RECT 682.735 216.560 683.065 217.040 ;
      LAYER li1 ;
        RECT 683.235 216.390 683.405 216.870 ;
      LAYER li1 ;
        RECT 683.575 216.560 683.905 217.040 ;
      LAYER li1 ;
        RECT 684.075 216.390 684.245 216.870 ;
      LAYER li1 ;
        RECT 684.415 216.560 684.745 217.040 ;
      LAYER li1 ;
        RECT 684.915 216.390 685.085 216.870 ;
      LAYER li1 ;
        RECT 685.255 216.560 685.585 217.040 ;
        RECT 685.755 216.390 685.925 216.865 ;
        RECT 686.095 216.560 686.425 217.040 ;
        RECT 686.595 216.390 686.765 216.870 ;
      LAYER li1 ;
        RECT 682.395 216.220 685.085 216.390 ;
      LAYER li1 ;
        RECT 685.345 216.220 686.765 216.390 ;
        RECT 687.025 216.315 687.315 217.040 ;
        RECT 687.875 216.240 688.205 217.040 ;
      LAYER li1 ;
        RECT 688.375 216.390 688.545 216.870 ;
      LAYER li1 ;
        RECT 688.715 216.560 689.045 217.040 ;
      LAYER li1 ;
        RECT 689.215 216.390 689.385 216.870 ;
      LAYER li1 ;
        RECT 689.555 216.560 689.885 217.040 ;
      LAYER li1 ;
        RECT 690.055 216.390 690.225 216.870 ;
      LAYER li1 ;
        RECT 690.395 216.560 690.725 217.040 ;
      LAYER li1 ;
        RECT 690.895 216.390 691.065 216.870 ;
      LAYER li1 ;
        RECT 691.235 216.560 691.565 217.040 ;
        RECT 691.735 216.390 691.905 216.865 ;
        RECT 692.075 216.560 692.405 217.040 ;
        RECT 692.575 216.390 692.745 216.870 ;
      LAYER li1 ;
        RECT 688.375 216.220 691.065 216.390 ;
      LAYER li1 ;
        RECT 691.325 216.220 692.745 216.390 ;
        RECT 693.005 216.315 693.295 217.040 ;
        RECT 693.855 216.240 694.185 217.040 ;
      LAYER li1 ;
        RECT 694.355 216.390 694.525 216.870 ;
      LAYER li1 ;
        RECT 694.695 216.560 695.025 217.040 ;
      LAYER li1 ;
        RECT 695.195 216.390 695.365 216.870 ;
      LAYER li1 ;
        RECT 695.535 216.560 695.865 217.040 ;
      LAYER li1 ;
        RECT 696.035 216.390 696.205 216.870 ;
      LAYER li1 ;
        RECT 696.375 216.560 696.705 217.040 ;
      LAYER li1 ;
        RECT 696.875 216.390 697.045 216.870 ;
      LAYER li1 ;
        RECT 697.215 216.560 697.545 217.040 ;
        RECT 697.715 216.390 697.885 216.865 ;
        RECT 698.055 216.560 698.385 217.040 ;
        RECT 698.555 216.390 698.725 216.870 ;
      LAYER li1 ;
        RECT 694.355 216.220 697.045 216.390 ;
      LAYER li1 ;
        RECT 697.305 216.220 698.725 216.390 ;
        RECT 698.985 216.315 699.275 217.040 ;
        RECT 699.835 216.240 700.165 217.040 ;
      LAYER li1 ;
        RECT 700.335 216.390 700.505 216.870 ;
      LAYER li1 ;
        RECT 700.675 216.560 701.005 217.040 ;
      LAYER li1 ;
        RECT 701.175 216.390 701.345 216.870 ;
      LAYER li1 ;
        RECT 701.515 216.560 701.845 217.040 ;
      LAYER li1 ;
        RECT 702.015 216.390 702.185 216.870 ;
      LAYER li1 ;
        RECT 702.355 216.560 702.685 217.040 ;
      LAYER li1 ;
        RECT 702.855 216.390 703.025 216.870 ;
      LAYER li1 ;
        RECT 703.195 216.560 703.525 217.040 ;
        RECT 703.695 216.390 703.865 216.865 ;
        RECT 704.035 216.560 704.365 217.040 ;
        RECT 704.535 216.390 704.705 216.870 ;
      LAYER li1 ;
        RECT 700.335 216.220 703.025 216.390 ;
      LAYER li1 ;
        RECT 703.285 216.220 704.705 216.390 ;
        RECT 704.965 216.315 705.255 217.040 ;
        RECT 705.815 216.240 706.145 217.040 ;
      LAYER li1 ;
        RECT 706.315 216.390 706.485 216.870 ;
      LAYER li1 ;
        RECT 706.655 216.560 706.985 217.040 ;
      LAYER li1 ;
        RECT 707.155 216.390 707.325 216.870 ;
      LAYER li1 ;
        RECT 707.495 216.560 707.825 217.040 ;
      LAYER li1 ;
        RECT 707.995 216.390 708.165 216.870 ;
      LAYER li1 ;
        RECT 708.335 216.560 708.665 217.040 ;
      LAYER li1 ;
        RECT 708.835 216.390 709.005 216.870 ;
      LAYER li1 ;
        RECT 709.175 216.560 709.505 217.040 ;
        RECT 709.675 216.390 709.845 216.865 ;
        RECT 710.015 216.560 710.345 217.040 ;
        RECT 710.515 216.390 710.685 216.870 ;
      LAYER li1 ;
        RECT 706.315 216.220 709.005 216.390 ;
      LAYER li1 ;
        RECT 709.265 216.220 710.685 216.390 ;
        RECT 710.945 216.315 711.235 217.040 ;
        RECT 711.795 216.240 712.125 217.040 ;
      LAYER li1 ;
        RECT 712.295 216.390 712.465 216.870 ;
      LAYER li1 ;
        RECT 712.635 216.560 712.965 217.040 ;
      LAYER li1 ;
        RECT 713.135 216.390 713.305 216.870 ;
      LAYER li1 ;
        RECT 713.475 216.560 713.805 217.040 ;
      LAYER li1 ;
        RECT 713.975 216.390 714.145 216.870 ;
      LAYER li1 ;
        RECT 714.315 216.560 714.645 217.040 ;
      LAYER li1 ;
        RECT 714.815 216.390 714.985 216.870 ;
      LAYER li1 ;
        RECT 715.155 216.560 715.485 217.040 ;
        RECT 715.655 216.390 715.825 216.865 ;
        RECT 715.995 216.560 716.325 217.040 ;
        RECT 716.495 216.390 716.665 216.870 ;
      LAYER li1 ;
        RECT 712.295 216.220 714.985 216.390 ;
      LAYER li1 ;
        RECT 715.245 216.220 716.665 216.390 ;
        RECT 716.925 216.315 717.215 217.040 ;
        RECT 717.775 216.240 718.105 217.040 ;
      LAYER li1 ;
        RECT 718.275 216.390 718.445 216.870 ;
      LAYER li1 ;
        RECT 718.615 216.560 718.945 217.040 ;
      LAYER li1 ;
        RECT 719.115 216.390 719.285 216.870 ;
      LAYER li1 ;
        RECT 719.455 216.560 719.785 217.040 ;
      LAYER li1 ;
        RECT 719.955 216.390 720.125 216.870 ;
      LAYER li1 ;
        RECT 720.295 216.560 720.625 217.040 ;
      LAYER li1 ;
        RECT 720.795 216.390 720.965 216.870 ;
      LAYER li1 ;
        RECT 721.135 216.560 721.465 217.040 ;
        RECT 721.635 216.390 721.805 216.865 ;
        RECT 721.975 216.560 722.305 217.040 ;
        RECT 722.475 216.390 722.645 216.870 ;
      LAYER li1 ;
        RECT 718.275 216.220 720.965 216.390 ;
      LAYER li1 ;
        RECT 721.225 216.220 722.645 216.390 ;
        RECT 722.905 216.315 723.195 217.040 ;
        RECT 723.755 216.240 724.085 217.040 ;
      LAYER li1 ;
        RECT 724.255 216.390 724.425 216.870 ;
      LAYER li1 ;
        RECT 724.595 216.560 724.925 217.040 ;
      LAYER li1 ;
        RECT 725.095 216.390 725.265 216.870 ;
      LAYER li1 ;
        RECT 725.435 216.560 725.765 217.040 ;
      LAYER li1 ;
        RECT 725.935 216.390 726.105 216.870 ;
      LAYER li1 ;
        RECT 726.275 216.560 726.605 217.040 ;
      LAYER li1 ;
        RECT 726.775 216.390 726.945 216.870 ;
      LAYER li1 ;
        RECT 727.115 216.560 727.445 217.040 ;
        RECT 727.615 216.390 727.785 216.865 ;
        RECT 727.955 216.560 728.285 217.040 ;
        RECT 728.455 216.390 728.625 216.870 ;
      LAYER li1 ;
        RECT 724.255 216.220 726.945 216.390 ;
      LAYER li1 ;
        RECT 727.205 216.220 728.625 216.390 ;
        RECT 728.885 216.315 729.175 217.040 ;
        RECT 729.735 216.240 730.065 217.040 ;
      LAYER li1 ;
        RECT 730.235 216.390 730.405 216.870 ;
      LAYER li1 ;
        RECT 730.575 216.560 730.905 217.040 ;
      LAYER li1 ;
        RECT 731.075 216.390 731.245 216.870 ;
      LAYER li1 ;
        RECT 731.415 216.560 731.745 217.040 ;
      LAYER li1 ;
        RECT 731.915 216.390 732.085 216.870 ;
      LAYER li1 ;
        RECT 732.255 216.560 732.585 217.040 ;
      LAYER li1 ;
        RECT 732.755 216.390 732.925 216.870 ;
      LAYER li1 ;
        RECT 733.095 216.560 733.425 217.040 ;
        RECT 733.595 216.390 733.765 216.865 ;
        RECT 733.935 216.560 734.265 217.040 ;
        RECT 734.435 216.390 734.605 216.870 ;
      LAYER li1 ;
        RECT 730.235 216.220 732.925 216.390 ;
      LAYER li1 ;
        RECT 733.185 216.220 734.605 216.390 ;
        RECT 734.865 216.315 735.155 217.040 ;
        RECT 735.715 216.240 736.045 217.040 ;
      LAYER li1 ;
        RECT 736.215 216.390 736.385 216.870 ;
      LAYER li1 ;
        RECT 736.555 216.560 736.885 217.040 ;
      LAYER li1 ;
        RECT 737.055 216.390 737.225 216.870 ;
      LAYER li1 ;
        RECT 737.395 216.560 737.725 217.040 ;
      LAYER li1 ;
        RECT 737.895 216.390 738.065 216.870 ;
      LAYER li1 ;
        RECT 738.235 216.560 738.565 217.040 ;
      LAYER li1 ;
        RECT 738.735 216.390 738.905 216.870 ;
      LAYER li1 ;
        RECT 739.075 216.560 739.405 217.040 ;
        RECT 739.575 216.390 739.745 216.865 ;
        RECT 739.915 216.560 740.245 217.040 ;
        RECT 740.415 216.390 740.585 216.870 ;
      LAYER li1 ;
        RECT 736.215 216.220 738.905 216.390 ;
      LAYER li1 ;
        RECT 739.165 216.220 740.585 216.390 ;
        RECT 740.845 216.315 741.135 217.040 ;
        RECT 741.695 216.240 742.025 217.040 ;
      LAYER li1 ;
        RECT 742.195 216.390 742.365 216.870 ;
      LAYER li1 ;
        RECT 742.535 216.560 742.865 217.040 ;
      LAYER li1 ;
        RECT 743.035 216.390 743.205 216.870 ;
      LAYER li1 ;
        RECT 743.375 216.560 743.705 217.040 ;
      LAYER li1 ;
        RECT 743.875 216.390 744.045 216.870 ;
      LAYER li1 ;
        RECT 744.215 216.560 744.545 217.040 ;
      LAYER li1 ;
        RECT 744.715 216.390 744.885 216.870 ;
      LAYER li1 ;
        RECT 745.055 216.560 745.385 217.040 ;
        RECT 745.555 216.390 745.725 216.865 ;
        RECT 745.895 216.560 746.225 217.040 ;
        RECT 746.395 216.390 746.565 216.870 ;
      LAYER li1 ;
        RECT 742.195 216.220 744.885 216.390 ;
      LAYER li1 ;
        RECT 745.145 216.220 746.565 216.390 ;
        RECT 746.825 216.315 747.115 217.040 ;
        RECT 747.675 216.240 748.005 217.040 ;
      LAYER li1 ;
        RECT 748.175 216.390 748.345 216.870 ;
      LAYER li1 ;
        RECT 748.515 216.560 748.845 217.040 ;
      LAYER li1 ;
        RECT 749.015 216.390 749.185 216.870 ;
      LAYER li1 ;
        RECT 749.355 216.560 749.685 217.040 ;
      LAYER li1 ;
        RECT 749.855 216.390 750.025 216.870 ;
      LAYER li1 ;
        RECT 750.195 216.560 750.525 217.040 ;
      LAYER li1 ;
        RECT 750.695 216.390 750.865 216.870 ;
      LAYER li1 ;
        RECT 751.035 216.560 751.365 217.040 ;
        RECT 751.535 216.390 751.705 216.865 ;
        RECT 751.875 216.560 752.205 217.040 ;
        RECT 752.375 216.390 752.545 216.870 ;
      LAYER li1 ;
        RECT 748.175 216.220 750.865 216.390 ;
      LAYER li1 ;
        RECT 751.125 216.220 752.545 216.390 ;
        RECT 752.805 216.315 753.095 217.040 ;
        RECT 753.655 216.240 753.985 217.040 ;
      LAYER li1 ;
        RECT 754.155 216.390 754.325 216.870 ;
      LAYER li1 ;
        RECT 754.495 216.560 754.825 217.040 ;
      LAYER li1 ;
        RECT 754.995 216.390 755.165 216.870 ;
      LAYER li1 ;
        RECT 755.335 216.560 755.665 217.040 ;
      LAYER li1 ;
        RECT 755.835 216.390 756.005 216.870 ;
      LAYER li1 ;
        RECT 756.175 216.560 756.505 217.040 ;
      LAYER li1 ;
        RECT 756.675 216.390 756.845 216.870 ;
      LAYER li1 ;
        RECT 757.015 216.560 757.345 217.040 ;
        RECT 757.515 216.390 757.685 216.865 ;
        RECT 757.855 216.560 758.185 217.040 ;
        RECT 758.355 216.390 758.525 216.870 ;
      LAYER li1 ;
        RECT 754.155 216.220 756.845 216.390 ;
      LAYER li1 ;
        RECT 757.105 216.220 758.525 216.390 ;
        RECT 758.785 216.315 759.075 217.040 ;
        RECT 759.635 216.240 759.965 217.040 ;
        RECT 760.475 216.560 760.805 217.040 ;
        RECT 761.315 216.560 761.645 217.040 ;
        RECT 762.155 216.560 762.485 217.040 ;
        RECT 762.995 216.560 763.325 217.040 ;
        RECT 763.495 216.390 763.665 216.865 ;
        RECT 763.835 216.560 764.165 217.040 ;
        RECT 764.335 216.390 764.505 216.870 ;
        RECT 763.085 216.220 764.505 216.390 ;
        RECT 764.765 216.315 765.055 217.040 ;
        RECT 765.615 216.240 765.945 217.040 ;
        RECT 766.455 216.560 766.785 217.040 ;
        RECT 767.295 216.560 767.625 217.040 ;
        RECT 768.135 216.560 768.465 217.040 ;
        RECT 768.975 216.560 769.305 217.040 ;
        RECT 769.475 216.390 769.645 216.865 ;
        RECT 769.815 216.560 770.145 217.040 ;
        RECT 770.315 216.390 770.485 216.870 ;
        RECT 769.065 216.220 770.485 216.390 ;
        RECT 770.745 216.315 771.035 217.040 ;
        RECT 771.595 216.240 771.925 217.040 ;
        RECT 772.435 216.560 772.765 217.040 ;
        RECT 773.275 216.560 773.605 217.040 ;
        RECT 774.115 216.560 774.445 217.040 ;
        RECT 774.955 216.560 775.285 217.040 ;
        RECT 775.455 216.390 775.625 216.865 ;
        RECT 775.795 216.560 776.125 217.040 ;
        RECT 776.295 216.390 776.465 216.870 ;
        RECT 775.045 216.220 776.465 216.390 ;
        RECT 776.725 216.315 777.015 217.040 ;
        RECT 777.575 216.240 777.905 217.040 ;
        RECT 778.415 216.560 778.745 217.040 ;
        RECT 779.255 216.560 779.585 217.040 ;
        RECT 780.095 216.560 780.425 217.040 ;
        RECT 780.935 216.560 781.265 217.040 ;
        RECT 781.435 216.390 781.605 216.865 ;
        RECT 781.775 216.560 782.105 217.040 ;
        RECT 782.275 216.390 782.445 216.870 ;
        RECT 781.025 216.220 782.445 216.390 ;
        RECT 782.705 216.315 782.995 217.040 ;
        RECT 783.555 216.240 783.885 217.040 ;
        RECT 784.395 216.560 784.725 217.040 ;
        RECT 785.235 216.560 785.565 217.040 ;
        RECT 786.075 216.560 786.405 217.040 ;
        RECT 786.915 216.560 787.245 217.040 ;
        RECT 787.415 216.390 787.585 216.865 ;
        RECT 787.755 216.560 788.085 217.040 ;
        RECT 788.255 216.390 788.425 216.870 ;
        RECT 787.005 216.220 788.425 216.390 ;
        RECT 788.685 216.315 788.975 217.040 ;
        RECT 789.535 216.240 789.865 217.040 ;
        RECT 790.375 216.560 790.705 217.040 ;
        RECT 791.215 216.560 791.545 217.040 ;
        RECT 792.055 216.560 792.385 217.040 ;
        RECT 792.895 216.560 793.225 217.040 ;
        RECT 793.395 216.390 793.565 216.865 ;
        RECT 793.735 216.560 794.065 217.040 ;
        RECT 794.235 216.390 794.405 216.870 ;
        RECT 792.985 216.220 794.405 216.390 ;
        RECT 794.665 216.315 794.955 217.040 ;
        RECT 2146.085 216.315 2146.375 217.040 ;
        RECT 2146.935 216.240 2147.265 217.040 ;
      LAYER li1 ;
        RECT 2147.435 216.390 2147.605 216.870 ;
      LAYER li1 ;
        RECT 2147.775 216.560 2148.105 217.040 ;
      LAYER li1 ;
        RECT 2148.275 216.390 2148.445 216.870 ;
      LAYER li1 ;
        RECT 2148.615 216.560 2148.945 217.040 ;
      LAYER li1 ;
        RECT 2149.115 216.390 2149.285 216.870 ;
      LAYER li1 ;
        RECT 2149.455 216.560 2149.785 217.040 ;
      LAYER li1 ;
        RECT 2149.955 216.390 2150.125 216.870 ;
      LAYER li1 ;
        RECT 2150.295 216.560 2150.625 217.040 ;
        RECT 2150.795 216.390 2150.965 216.865 ;
        RECT 2151.135 216.560 2151.465 217.040 ;
        RECT 2151.635 216.390 2151.805 216.870 ;
      LAYER li1 ;
        RECT 2147.435 216.220 2150.125 216.390 ;
      LAYER li1 ;
        RECT 2150.385 216.220 2151.805 216.390 ;
        RECT 2152.065 216.315 2152.355 217.040 ;
        RECT 2152.915 216.240 2153.245 217.040 ;
      LAYER li1 ;
        RECT 2153.415 216.390 2153.585 216.870 ;
      LAYER li1 ;
        RECT 2153.755 216.560 2154.085 217.040 ;
      LAYER li1 ;
        RECT 2154.255 216.390 2154.425 216.870 ;
      LAYER li1 ;
        RECT 2154.595 216.560 2154.925 217.040 ;
      LAYER li1 ;
        RECT 2155.095 216.390 2155.265 216.870 ;
      LAYER li1 ;
        RECT 2155.435 216.560 2155.765 217.040 ;
      LAYER li1 ;
        RECT 2155.935 216.390 2156.105 216.870 ;
      LAYER li1 ;
        RECT 2156.275 216.560 2156.605 217.040 ;
        RECT 2156.775 216.390 2156.945 216.865 ;
        RECT 2157.115 216.560 2157.445 217.040 ;
        RECT 2157.615 216.390 2157.785 216.870 ;
      LAYER li1 ;
        RECT 2153.415 216.220 2156.105 216.390 ;
      LAYER li1 ;
        RECT 2156.365 216.220 2157.785 216.390 ;
        RECT 2158.045 216.315 2158.335 217.040 ;
        RECT 2158.895 216.240 2159.225 217.040 ;
      LAYER li1 ;
        RECT 2159.395 216.390 2159.565 216.870 ;
      LAYER li1 ;
        RECT 2159.735 216.560 2160.065 217.040 ;
      LAYER li1 ;
        RECT 2160.235 216.390 2160.405 216.870 ;
      LAYER li1 ;
        RECT 2160.575 216.560 2160.905 217.040 ;
      LAYER li1 ;
        RECT 2161.075 216.390 2161.245 216.870 ;
      LAYER li1 ;
        RECT 2161.415 216.560 2161.745 217.040 ;
      LAYER li1 ;
        RECT 2161.915 216.390 2162.085 216.870 ;
      LAYER li1 ;
        RECT 2162.255 216.560 2162.585 217.040 ;
        RECT 2162.755 216.390 2162.925 216.865 ;
        RECT 2163.095 216.560 2163.425 217.040 ;
        RECT 2163.595 216.390 2163.765 216.870 ;
      LAYER li1 ;
        RECT 2159.395 216.220 2162.085 216.390 ;
      LAYER li1 ;
        RECT 2162.345 216.220 2163.765 216.390 ;
        RECT 2164.025 216.315 2164.315 217.040 ;
        RECT 2164.875 216.240 2165.205 217.040 ;
      LAYER li1 ;
        RECT 2165.375 216.390 2165.545 216.870 ;
      LAYER li1 ;
        RECT 2165.715 216.560 2166.045 217.040 ;
      LAYER li1 ;
        RECT 2166.215 216.390 2166.385 216.870 ;
      LAYER li1 ;
        RECT 2166.555 216.560 2166.885 217.040 ;
      LAYER li1 ;
        RECT 2167.055 216.390 2167.225 216.870 ;
      LAYER li1 ;
        RECT 2167.395 216.560 2167.725 217.040 ;
      LAYER li1 ;
        RECT 2167.895 216.390 2168.065 216.870 ;
      LAYER li1 ;
        RECT 2168.235 216.560 2168.565 217.040 ;
        RECT 2168.735 216.390 2168.905 216.865 ;
        RECT 2169.075 216.560 2169.405 217.040 ;
        RECT 2169.575 216.390 2169.745 216.870 ;
      LAYER li1 ;
        RECT 2165.375 216.220 2168.065 216.390 ;
      LAYER li1 ;
        RECT 2168.325 216.220 2169.745 216.390 ;
        RECT 2170.005 216.315 2170.295 217.040 ;
        RECT 2170.855 216.240 2171.185 217.040 ;
      LAYER li1 ;
        RECT 2171.355 216.390 2171.525 216.870 ;
      LAYER li1 ;
        RECT 2171.695 216.560 2172.025 217.040 ;
      LAYER li1 ;
        RECT 2172.195 216.390 2172.365 216.870 ;
      LAYER li1 ;
        RECT 2172.535 216.560 2172.865 217.040 ;
      LAYER li1 ;
        RECT 2173.035 216.390 2173.205 216.870 ;
      LAYER li1 ;
        RECT 2173.375 216.560 2173.705 217.040 ;
      LAYER li1 ;
        RECT 2173.875 216.390 2174.045 216.870 ;
      LAYER li1 ;
        RECT 2174.215 216.560 2174.545 217.040 ;
        RECT 2174.715 216.390 2174.885 216.865 ;
        RECT 2175.055 216.560 2175.385 217.040 ;
        RECT 2175.555 216.390 2175.725 216.870 ;
      LAYER li1 ;
        RECT 2171.355 216.220 2174.045 216.390 ;
      LAYER li1 ;
        RECT 2174.305 216.220 2175.725 216.390 ;
        RECT 2175.985 216.315 2176.275 217.040 ;
        RECT 2176.835 216.240 2177.165 217.040 ;
      LAYER li1 ;
        RECT 2177.335 216.390 2177.505 216.870 ;
      LAYER li1 ;
        RECT 2177.675 216.560 2178.005 217.040 ;
      LAYER li1 ;
        RECT 2178.175 216.390 2178.345 216.870 ;
      LAYER li1 ;
        RECT 2178.515 216.560 2178.845 217.040 ;
      LAYER li1 ;
        RECT 2179.015 216.390 2179.185 216.870 ;
      LAYER li1 ;
        RECT 2179.355 216.560 2179.685 217.040 ;
      LAYER li1 ;
        RECT 2179.855 216.390 2180.025 216.870 ;
      LAYER li1 ;
        RECT 2180.195 216.560 2180.525 217.040 ;
        RECT 2180.695 216.390 2180.865 216.865 ;
        RECT 2181.035 216.560 2181.365 217.040 ;
        RECT 2181.535 216.390 2181.705 216.870 ;
      LAYER li1 ;
        RECT 2177.335 216.220 2180.025 216.390 ;
      LAYER li1 ;
        RECT 2180.285 216.220 2181.705 216.390 ;
        RECT 2181.965 216.315 2182.255 217.040 ;
        RECT 2182.815 216.240 2183.145 217.040 ;
      LAYER li1 ;
        RECT 2183.315 216.390 2183.485 216.870 ;
      LAYER li1 ;
        RECT 2183.655 216.560 2183.985 217.040 ;
      LAYER li1 ;
        RECT 2184.155 216.390 2184.325 216.870 ;
      LAYER li1 ;
        RECT 2184.495 216.560 2184.825 217.040 ;
      LAYER li1 ;
        RECT 2184.995 216.390 2185.165 216.870 ;
      LAYER li1 ;
        RECT 2185.335 216.560 2185.665 217.040 ;
      LAYER li1 ;
        RECT 2185.835 216.390 2186.005 216.870 ;
      LAYER li1 ;
        RECT 2186.175 216.560 2186.505 217.040 ;
        RECT 2186.675 216.390 2186.845 216.865 ;
        RECT 2187.015 216.560 2187.345 217.040 ;
        RECT 2187.515 216.390 2187.685 216.870 ;
      LAYER li1 ;
        RECT 2183.315 216.220 2186.005 216.390 ;
      LAYER li1 ;
        RECT 2186.265 216.220 2187.685 216.390 ;
        RECT 2187.945 216.315 2188.235 217.040 ;
        RECT 2188.795 216.240 2189.125 217.040 ;
      LAYER li1 ;
        RECT 2189.295 216.390 2189.465 216.870 ;
      LAYER li1 ;
        RECT 2189.635 216.560 2189.965 217.040 ;
      LAYER li1 ;
        RECT 2190.135 216.390 2190.305 216.870 ;
      LAYER li1 ;
        RECT 2190.475 216.560 2190.805 217.040 ;
      LAYER li1 ;
        RECT 2190.975 216.390 2191.145 216.870 ;
      LAYER li1 ;
        RECT 2191.315 216.560 2191.645 217.040 ;
      LAYER li1 ;
        RECT 2191.815 216.390 2191.985 216.870 ;
      LAYER li1 ;
        RECT 2192.155 216.560 2192.485 217.040 ;
        RECT 2192.655 216.390 2192.825 216.865 ;
        RECT 2192.995 216.560 2193.325 217.040 ;
        RECT 2193.495 216.390 2193.665 216.870 ;
      LAYER li1 ;
        RECT 2189.295 216.220 2191.985 216.390 ;
      LAYER li1 ;
        RECT 2192.245 216.220 2193.665 216.390 ;
        RECT 2193.925 216.315 2194.215 217.040 ;
        RECT 2194.775 216.240 2195.105 217.040 ;
      LAYER li1 ;
        RECT 2195.275 216.390 2195.445 216.870 ;
      LAYER li1 ;
        RECT 2195.615 216.560 2195.945 217.040 ;
      LAYER li1 ;
        RECT 2196.115 216.390 2196.285 216.870 ;
      LAYER li1 ;
        RECT 2196.455 216.560 2196.785 217.040 ;
      LAYER li1 ;
        RECT 2196.955 216.390 2197.125 216.870 ;
      LAYER li1 ;
        RECT 2197.295 216.560 2197.625 217.040 ;
      LAYER li1 ;
        RECT 2197.795 216.390 2197.965 216.870 ;
      LAYER li1 ;
        RECT 2198.135 216.560 2198.465 217.040 ;
        RECT 2198.635 216.390 2198.805 216.865 ;
        RECT 2198.975 216.560 2199.305 217.040 ;
        RECT 2199.475 216.390 2199.645 216.870 ;
      LAYER li1 ;
        RECT 2195.275 216.220 2197.965 216.390 ;
      LAYER li1 ;
        RECT 2198.225 216.220 2199.645 216.390 ;
        RECT 2199.905 216.315 2200.195 217.040 ;
        RECT 2200.755 216.240 2201.085 217.040 ;
      LAYER li1 ;
        RECT 2201.255 216.390 2201.425 216.870 ;
      LAYER li1 ;
        RECT 2201.595 216.560 2201.925 217.040 ;
      LAYER li1 ;
        RECT 2202.095 216.390 2202.265 216.870 ;
      LAYER li1 ;
        RECT 2202.435 216.560 2202.765 217.040 ;
      LAYER li1 ;
        RECT 2202.935 216.390 2203.105 216.870 ;
      LAYER li1 ;
        RECT 2203.275 216.560 2203.605 217.040 ;
      LAYER li1 ;
        RECT 2203.775 216.390 2203.945 216.870 ;
      LAYER li1 ;
        RECT 2204.115 216.560 2204.445 217.040 ;
        RECT 2204.615 216.390 2204.785 216.865 ;
        RECT 2204.955 216.560 2205.285 217.040 ;
        RECT 2205.455 216.390 2205.625 216.870 ;
      LAYER li1 ;
        RECT 2201.255 216.220 2203.945 216.390 ;
      LAYER li1 ;
        RECT 2204.205 216.220 2205.625 216.390 ;
        RECT 2205.885 216.315 2206.175 217.040 ;
        RECT 2206.735 216.240 2207.065 217.040 ;
      LAYER li1 ;
        RECT 2207.235 216.390 2207.405 216.870 ;
      LAYER li1 ;
        RECT 2207.575 216.560 2207.905 217.040 ;
      LAYER li1 ;
        RECT 2208.075 216.390 2208.245 216.870 ;
      LAYER li1 ;
        RECT 2208.415 216.560 2208.745 217.040 ;
      LAYER li1 ;
        RECT 2208.915 216.390 2209.085 216.870 ;
      LAYER li1 ;
        RECT 2209.255 216.560 2209.585 217.040 ;
      LAYER li1 ;
        RECT 2209.755 216.390 2209.925 216.870 ;
      LAYER li1 ;
        RECT 2210.095 216.560 2210.425 217.040 ;
        RECT 2210.595 216.390 2210.765 216.865 ;
        RECT 2210.935 216.560 2211.265 217.040 ;
        RECT 2211.435 216.390 2211.605 216.870 ;
      LAYER li1 ;
        RECT 2207.235 216.220 2209.925 216.390 ;
      LAYER li1 ;
        RECT 2210.185 216.220 2211.605 216.390 ;
        RECT 2211.865 216.315 2212.155 217.040 ;
        RECT 2212.715 216.240 2213.045 217.040 ;
      LAYER li1 ;
        RECT 2213.215 216.390 2213.385 216.870 ;
      LAYER li1 ;
        RECT 2213.555 216.560 2213.885 217.040 ;
      LAYER li1 ;
        RECT 2214.055 216.390 2214.225 216.870 ;
      LAYER li1 ;
        RECT 2214.395 216.560 2214.725 217.040 ;
      LAYER li1 ;
        RECT 2214.895 216.390 2215.065 216.870 ;
      LAYER li1 ;
        RECT 2215.235 216.560 2215.565 217.040 ;
      LAYER li1 ;
        RECT 2215.735 216.390 2215.905 216.870 ;
      LAYER li1 ;
        RECT 2216.075 216.560 2216.405 217.040 ;
        RECT 2216.575 216.390 2216.745 216.865 ;
        RECT 2216.915 216.560 2217.245 217.040 ;
        RECT 2217.415 216.390 2217.585 216.870 ;
      LAYER li1 ;
        RECT 2213.215 216.220 2215.905 216.390 ;
      LAYER li1 ;
        RECT 2216.165 216.220 2217.585 216.390 ;
        RECT 2217.845 216.315 2218.135 217.040 ;
        RECT 2218.695 216.240 2219.025 217.040 ;
      LAYER li1 ;
        RECT 2219.195 216.390 2219.365 216.870 ;
      LAYER li1 ;
        RECT 2219.535 216.560 2219.865 217.040 ;
      LAYER li1 ;
        RECT 2220.035 216.390 2220.205 216.870 ;
      LAYER li1 ;
        RECT 2220.375 216.560 2220.705 217.040 ;
      LAYER li1 ;
        RECT 2220.875 216.390 2221.045 216.870 ;
      LAYER li1 ;
        RECT 2221.215 216.560 2221.545 217.040 ;
      LAYER li1 ;
        RECT 2221.715 216.390 2221.885 216.870 ;
      LAYER li1 ;
        RECT 2222.055 216.560 2222.385 217.040 ;
        RECT 2222.555 216.390 2222.725 216.865 ;
        RECT 2222.895 216.560 2223.225 217.040 ;
        RECT 2223.395 216.390 2223.565 216.870 ;
      LAYER li1 ;
        RECT 2219.195 216.220 2221.885 216.390 ;
      LAYER li1 ;
        RECT 2222.145 216.220 2223.565 216.390 ;
        RECT 2223.825 216.315 2224.115 217.040 ;
        RECT 2224.675 216.240 2225.005 217.040 ;
      LAYER li1 ;
        RECT 2225.175 216.390 2225.345 216.870 ;
      LAYER li1 ;
        RECT 2225.515 216.560 2225.845 217.040 ;
      LAYER li1 ;
        RECT 2226.015 216.390 2226.185 216.870 ;
      LAYER li1 ;
        RECT 2226.355 216.560 2226.685 217.040 ;
      LAYER li1 ;
        RECT 2226.855 216.390 2227.025 216.870 ;
      LAYER li1 ;
        RECT 2227.195 216.560 2227.525 217.040 ;
      LAYER li1 ;
        RECT 2227.695 216.390 2227.865 216.870 ;
      LAYER li1 ;
        RECT 2228.035 216.560 2228.365 217.040 ;
        RECT 2228.535 216.390 2228.705 216.865 ;
        RECT 2228.875 216.560 2229.205 217.040 ;
        RECT 2229.375 216.390 2229.545 216.870 ;
      LAYER li1 ;
        RECT 2225.175 216.220 2227.865 216.390 ;
      LAYER li1 ;
        RECT 2228.125 216.220 2229.545 216.390 ;
        RECT 2229.805 216.315 2230.095 217.040 ;
        RECT 2230.655 216.240 2230.985 217.040 ;
      LAYER li1 ;
        RECT 2231.155 216.390 2231.325 216.870 ;
      LAYER li1 ;
        RECT 2231.495 216.560 2231.825 217.040 ;
      LAYER li1 ;
        RECT 2231.995 216.390 2232.165 216.870 ;
      LAYER li1 ;
        RECT 2232.335 216.560 2232.665 217.040 ;
      LAYER li1 ;
        RECT 2232.835 216.390 2233.005 216.870 ;
      LAYER li1 ;
        RECT 2233.175 216.560 2233.505 217.040 ;
      LAYER li1 ;
        RECT 2233.675 216.390 2233.845 216.870 ;
      LAYER li1 ;
        RECT 2234.015 216.560 2234.345 217.040 ;
        RECT 2234.515 216.390 2234.685 216.865 ;
        RECT 2234.855 216.560 2235.185 217.040 ;
        RECT 2235.355 216.390 2235.525 216.870 ;
      LAYER li1 ;
        RECT 2231.155 216.220 2233.845 216.390 ;
      LAYER li1 ;
        RECT 2234.105 216.220 2235.525 216.390 ;
        RECT 2235.785 216.315 2236.075 217.040 ;
        RECT 2236.635 216.240 2236.965 217.040 ;
      LAYER li1 ;
        RECT 2237.135 216.390 2237.305 216.870 ;
      LAYER li1 ;
        RECT 2237.475 216.560 2237.805 217.040 ;
      LAYER li1 ;
        RECT 2237.975 216.390 2238.145 216.870 ;
      LAYER li1 ;
        RECT 2238.315 216.560 2238.645 217.040 ;
      LAYER li1 ;
        RECT 2238.815 216.390 2238.985 216.870 ;
      LAYER li1 ;
        RECT 2239.155 216.560 2239.485 217.040 ;
      LAYER li1 ;
        RECT 2239.655 216.390 2239.825 216.870 ;
      LAYER li1 ;
        RECT 2239.995 216.560 2240.325 217.040 ;
        RECT 2240.495 216.390 2240.665 216.865 ;
        RECT 2240.835 216.560 2241.165 217.040 ;
        RECT 2241.335 216.390 2241.505 216.870 ;
      LAYER li1 ;
        RECT 2237.135 216.220 2239.825 216.390 ;
      LAYER li1 ;
        RECT 2240.085 216.220 2241.505 216.390 ;
        RECT 2241.765 216.315 2242.055 217.040 ;
        RECT 2242.615 216.240 2242.945 217.040 ;
      LAYER li1 ;
        RECT 2243.115 216.390 2243.285 216.870 ;
      LAYER li1 ;
        RECT 2243.455 216.560 2243.785 217.040 ;
      LAYER li1 ;
        RECT 2243.955 216.390 2244.125 216.870 ;
      LAYER li1 ;
        RECT 2244.295 216.560 2244.625 217.040 ;
      LAYER li1 ;
        RECT 2244.795 216.390 2244.965 216.870 ;
      LAYER li1 ;
        RECT 2245.135 216.560 2245.465 217.040 ;
      LAYER li1 ;
        RECT 2245.635 216.390 2245.805 216.870 ;
      LAYER li1 ;
        RECT 2245.975 216.560 2246.305 217.040 ;
        RECT 2246.475 216.390 2246.645 216.865 ;
        RECT 2246.815 216.560 2247.145 217.040 ;
        RECT 2247.315 216.390 2247.485 216.870 ;
      LAYER li1 ;
        RECT 2243.115 216.220 2245.805 216.390 ;
      LAYER li1 ;
        RECT 2246.065 216.220 2247.485 216.390 ;
        RECT 2247.745 216.315 2248.035 217.040 ;
        RECT 2248.595 216.240 2248.925 217.040 ;
      LAYER li1 ;
        RECT 2249.095 216.390 2249.265 216.870 ;
      LAYER li1 ;
        RECT 2249.435 216.560 2249.765 217.040 ;
      LAYER li1 ;
        RECT 2249.935 216.390 2250.105 216.870 ;
      LAYER li1 ;
        RECT 2250.275 216.560 2250.605 217.040 ;
      LAYER li1 ;
        RECT 2250.775 216.390 2250.945 216.870 ;
      LAYER li1 ;
        RECT 2251.115 216.560 2251.445 217.040 ;
      LAYER li1 ;
        RECT 2251.615 216.390 2251.785 216.870 ;
      LAYER li1 ;
        RECT 2251.955 216.560 2252.285 217.040 ;
        RECT 2252.455 216.390 2252.625 216.865 ;
        RECT 2252.795 216.560 2253.125 217.040 ;
        RECT 2253.295 216.390 2253.465 216.870 ;
      LAYER li1 ;
        RECT 2249.095 216.220 2251.785 216.390 ;
      LAYER li1 ;
        RECT 2252.045 216.220 2253.465 216.390 ;
        RECT 2253.725 216.315 2254.015 217.040 ;
        RECT 2254.575 216.240 2254.905 217.040 ;
      LAYER li1 ;
        RECT 2255.075 216.390 2255.245 216.870 ;
      LAYER li1 ;
        RECT 2255.415 216.560 2255.745 217.040 ;
      LAYER li1 ;
        RECT 2255.915 216.390 2256.085 216.870 ;
      LAYER li1 ;
        RECT 2256.255 216.560 2256.585 217.040 ;
      LAYER li1 ;
        RECT 2256.755 216.390 2256.925 216.870 ;
      LAYER li1 ;
        RECT 2257.095 216.560 2257.425 217.040 ;
      LAYER li1 ;
        RECT 2257.595 216.390 2257.765 216.870 ;
      LAYER li1 ;
        RECT 2257.935 216.560 2258.265 217.040 ;
        RECT 2258.435 216.390 2258.605 216.865 ;
        RECT 2258.775 216.560 2259.105 217.040 ;
        RECT 2259.275 216.390 2259.445 216.870 ;
      LAYER li1 ;
        RECT 2255.075 216.220 2257.765 216.390 ;
      LAYER li1 ;
        RECT 2258.025 216.220 2259.445 216.390 ;
        RECT 2259.705 216.315 2259.995 217.040 ;
        RECT 2260.555 216.240 2260.885 217.040 ;
      LAYER li1 ;
        RECT 2261.055 216.390 2261.225 216.870 ;
      LAYER li1 ;
        RECT 2261.395 216.560 2261.725 217.040 ;
      LAYER li1 ;
        RECT 2261.895 216.390 2262.065 216.870 ;
      LAYER li1 ;
        RECT 2262.235 216.560 2262.565 217.040 ;
      LAYER li1 ;
        RECT 2262.735 216.390 2262.905 216.870 ;
      LAYER li1 ;
        RECT 2263.075 216.560 2263.405 217.040 ;
      LAYER li1 ;
        RECT 2263.575 216.390 2263.745 216.870 ;
      LAYER li1 ;
        RECT 2263.915 216.560 2264.245 217.040 ;
        RECT 2264.415 216.390 2264.585 216.865 ;
        RECT 2264.755 216.560 2265.085 217.040 ;
        RECT 2265.255 216.390 2265.425 216.870 ;
      LAYER li1 ;
        RECT 2261.055 216.220 2263.745 216.390 ;
      LAYER li1 ;
        RECT 2264.005 216.220 2265.425 216.390 ;
        RECT 2265.685 216.315 2265.975 217.040 ;
        RECT 2266.535 216.240 2266.865 217.040 ;
      LAYER li1 ;
        RECT 2267.035 216.390 2267.205 216.870 ;
      LAYER li1 ;
        RECT 2267.375 216.560 2267.705 217.040 ;
      LAYER li1 ;
        RECT 2267.875 216.390 2268.045 216.870 ;
      LAYER li1 ;
        RECT 2268.215 216.560 2268.545 217.040 ;
      LAYER li1 ;
        RECT 2268.715 216.390 2268.885 216.870 ;
      LAYER li1 ;
        RECT 2269.055 216.560 2269.385 217.040 ;
      LAYER li1 ;
        RECT 2269.555 216.390 2269.725 216.870 ;
      LAYER li1 ;
        RECT 2269.895 216.560 2270.225 217.040 ;
        RECT 2270.395 216.390 2270.565 216.865 ;
        RECT 2270.735 216.560 2271.065 217.040 ;
        RECT 2271.235 216.390 2271.405 216.870 ;
      LAYER li1 ;
        RECT 2267.035 216.220 2269.725 216.390 ;
      LAYER li1 ;
        RECT 2269.985 216.220 2271.405 216.390 ;
        RECT 2271.665 216.315 2271.955 217.040 ;
      LAYER li1 ;
        RECT 670.435 215.680 670.690 216.220 ;
      LAYER li1 ;
        RECT 673.385 216.050 673.560 216.220 ;
        RECT 670.935 215.880 673.560 216.050 ;
        RECT 673.385 215.680 673.560 215.880 ;
      LAYER li1 ;
        RECT 673.740 215.850 675.330 216.050 ;
        RECT 676.415 215.680 676.670 216.220 ;
      LAYER li1 ;
        RECT 679.365 216.050 679.540 216.220 ;
        RECT 676.915 215.880 679.540 216.050 ;
        RECT 679.365 215.680 679.540 215.880 ;
      LAYER li1 ;
        RECT 679.720 215.850 681.310 216.050 ;
        RECT 682.395 215.680 682.650 216.220 ;
      LAYER li1 ;
        RECT 685.345 216.050 685.520 216.220 ;
        RECT 682.895 215.880 685.520 216.050 ;
        RECT 685.345 215.680 685.520 215.880 ;
      LAYER li1 ;
        RECT 685.700 215.850 687.290 216.050 ;
        RECT 688.375 215.680 688.630 216.220 ;
      LAYER li1 ;
        RECT 691.325 216.050 691.500 216.220 ;
        RECT 688.875 215.880 691.500 216.050 ;
        RECT 691.325 215.680 691.500 215.880 ;
      LAYER li1 ;
        RECT 691.680 215.850 693.270 216.050 ;
        RECT 694.355 215.680 694.610 216.220 ;
      LAYER li1 ;
        RECT 697.305 216.050 697.480 216.220 ;
        RECT 694.855 215.880 697.480 216.050 ;
        RECT 697.305 215.680 697.480 215.880 ;
      LAYER li1 ;
        RECT 697.660 215.850 699.250 216.050 ;
        RECT 700.335 215.680 700.590 216.220 ;
      LAYER li1 ;
        RECT 703.285 216.050 703.460 216.220 ;
        RECT 700.835 215.880 703.460 216.050 ;
        RECT 703.285 215.680 703.460 215.880 ;
      LAYER li1 ;
        RECT 703.640 215.850 705.230 216.050 ;
        RECT 706.315 215.680 706.570 216.220 ;
      LAYER li1 ;
        RECT 709.265 216.050 709.440 216.220 ;
        RECT 706.815 215.880 709.440 216.050 ;
        RECT 709.265 215.680 709.440 215.880 ;
      LAYER li1 ;
        RECT 709.620 215.850 711.210 216.050 ;
        RECT 712.295 215.680 712.550 216.220 ;
      LAYER li1 ;
        RECT 715.245 216.050 715.420 216.220 ;
        RECT 712.795 215.880 715.420 216.050 ;
        RECT 715.245 215.680 715.420 215.880 ;
      LAYER li1 ;
        RECT 715.600 215.850 717.190 216.050 ;
        RECT 718.275 215.680 718.530 216.220 ;
      LAYER li1 ;
        RECT 721.225 216.050 721.400 216.220 ;
        RECT 718.775 215.880 721.400 216.050 ;
        RECT 721.225 215.680 721.400 215.880 ;
      LAYER li1 ;
        RECT 721.580 215.850 723.170 216.050 ;
        RECT 724.255 215.680 724.510 216.220 ;
      LAYER li1 ;
        RECT 727.205 216.050 727.380 216.220 ;
        RECT 724.755 215.880 727.380 216.050 ;
        RECT 727.205 215.680 727.380 215.880 ;
      LAYER li1 ;
        RECT 727.560 215.850 729.150 216.050 ;
        RECT 730.235 215.680 730.490 216.220 ;
      LAYER li1 ;
        RECT 733.185 216.050 733.360 216.220 ;
        RECT 730.735 215.880 733.360 216.050 ;
        RECT 733.185 215.680 733.360 215.880 ;
      LAYER li1 ;
        RECT 733.540 215.850 735.130 216.050 ;
        RECT 736.215 215.680 736.470 216.220 ;
      LAYER li1 ;
        RECT 739.165 216.050 739.340 216.220 ;
        RECT 736.715 215.880 739.340 216.050 ;
        RECT 739.165 215.680 739.340 215.880 ;
      LAYER li1 ;
        RECT 739.520 215.850 741.110 216.050 ;
        RECT 742.195 215.680 742.450 216.220 ;
      LAYER li1 ;
        RECT 745.145 216.050 745.320 216.220 ;
        RECT 742.695 215.880 745.320 216.050 ;
        RECT 745.145 215.680 745.320 215.880 ;
      LAYER li1 ;
        RECT 745.500 215.850 747.090 216.050 ;
        RECT 748.175 215.680 748.430 216.220 ;
      LAYER li1 ;
        RECT 751.125 216.050 751.300 216.220 ;
        RECT 748.675 215.880 751.300 216.050 ;
        RECT 751.125 215.680 751.300 215.880 ;
      LAYER li1 ;
        RECT 751.480 215.850 753.070 216.050 ;
        RECT 754.155 215.680 754.410 216.220 ;
      LAYER li1 ;
        RECT 757.105 216.050 757.280 216.220 ;
        RECT 763.085 216.050 763.260 216.220 ;
        RECT 769.065 216.050 769.240 216.220 ;
        RECT 775.045 216.050 775.220 216.220 ;
        RECT 781.025 216.050 781.200 216.220 ;
        RECT 787.005 216.050 787.180 216.220 ;
        RECT 792.985 216.050 793.160 216.220 ;
        RECT 754.655 215.880 757.280 216.050 ;
        RECT 757.105 215.680 757.280 215.880 ;
      LAYER li1 ;
        RECT 757.460 215.850 759.050 216.050 ;
      LAYER li1 ;
        RECT 760.635 215.880 763.260 216.050 ;
        RECT 763.085 215.680 763.260 215.880 ;
      LAYER li1 ;
        RECT 763.440 215.850 765.030 216.050 ;
      LAYER li1 ;
        RECT 766.615 215.880 769.240 216.050 ;
        RECT 769.065 215.680 769.240 215.880 ;
      LAYER li1 ;
        RECT 769.420 215.850 771.010 216.050 ;
      LAYER li1 ;
        RECT 772.595 215.880 775.220 216.050 ;
        RECT 775.045 215.680 775.220 215.880 ;
      LAYER li1 ;
        RECT 775.400 215.850 776.990 216.050 ;
      LAYER li1 ;
        RECT 778.575 215.880 781.200 216.050 ;
        RECT 781.025 215.680 781.200 215.880 ;
      LAYER li1 ;
        RECT 781.380 215.850 782.970 216.050 ;
      LAYER li1 ;
        RECT 784.555 215.880 787.180 216.050 ;
        RECT 787.005 215.680 787.180 215.880 ;
      LAYER li1 ;
        RECT 787.360 215.850 788.950 216.050 ;
      LAYER li1 ;
        RECT 790.535 215.880 793.160 216.050 ;
        RECT 792.985 215.680 793.160 215.880 ;
      LAYER li1 ;
        RECT 793.340 215.850 794.930 216.050 ;
        RECT 2147.435 215.680 2147.690 216.220 ;
      LAYER li1 ;
        RECT 2150.385 216.050 2150.560 216.220 ;
        RECT 2147.935 215.880 2150.560 216.050 ;
        RECT 2150.385 215.680 2150.560 215.880 ;
      LAYER li1 ;
        RECT 2153.415 215.680 2153.670 216.220 ;
      LAYER li1 ;
        RECT 2156.365 216.050 2156.540 216.220 ;
        RECT 2153.915 215.880 2156.540 216.050 ;
        RECT 2156.365 215.680 2156.540 215.880 ;
      LAYER li1 ;
        RECT 2159.395 215.680 2159.650 216.220 ;
      LAYER li1 ;
        RECT 2162.345 216.050 2162.520 216.220 ;
        RECT 2159.895 215.880 2162.520 216.050 ;
        RECT 2162.345 215.680 2162.520 215.880 ;
      LAYER li1 ;
        RECT 2165.375 215.680 2165.630 216.220 ;
      LAYER li1 ;
        RECT 2168.325 216.050 2168.500 216.220 ;
        RECT 2165.875 215.880 2168.500 216.050 ;
        RECT 2168.325 215.680 2168.500 215.880 ;
      LAYER li1 ;
        RECT 2171.355 215.680 2171.610 216.220 ;
      LAYER li1 ;
        RECT 2174.305 216.050 2174.480 216.220 ;
        RECT 2171.855 215.880 2174.480 216.050 ;
        RECT 2174.305 215.680 2174.480 215.880 ;
      LAYER li1 ;
        RECT 2177.335 215.680 2177.590 216.220 ;
      LAYER li1 ;
        RECT 2180.285 216.050 2180.460 216.220 ;
        RECT 2177.835 215.880 2180.460 216.050 ;
        RECT 2180.285 215.680 2180.460 215.880 ;
      LAYER li1 ;
        RECT 2183.315 215.680 2183.570 216.220 ;
      LAYER li1 ;
        RECT 2186.265 216.050 2186.440 216.220 ;
        RECT 2183.815 215.880 2186.440 216.050 ;
        RECT 2186.265 215.680 2186.440 215.880 ;
      LAYER li1 ;
        RECT 2189.295 215.680 2189.550 216.220 ;
      LAYER li1 ;
        RECT 2192.245 216.050 2192.420 216.220 ;
        RECT 2189.795 215.880 2192.420 216.050 ;
        RECT 2192.245 215.680 2192.420 215.880 ;
      LAYER li1 ;
        RECT 2195.275 215.680 2195.530 216.220 ;
      LAYER li1 ;
        RECT 2198.225 216.050 2198.400 216.220 ;
        RECT 2195.775 215.880 2198.400 216.050 ;
        RECT 2198.225 215.680 2198.400 215.880 ;
      LAYER li1 ;
        RECT 2201.255 215.680 2201.510 216.220 ;
      LAYER li1 ;
        RECT 2204.205 216.050 2204.380 216.220 ;
        RECT 2201.755 215.880 2204.380 216.050 ;
        RECT 2204.205 215.680 2204.380 215.880 ;
      LAYER li1 ;
        RECT 2207.235 215.680 2207.490 216.220 ;
      LAYER li1 ;
        RECT 2210.185 216.050 2210.360 216.220 ;
        RECT 2207.735 215.880 2210.360 216.050 ;
        RECT 2210.185 215.680 2210.360 215.880 ;
      LAYER li1 ;
        RECT 2213.215 215.680 2213.470 216.220 ;
      LAYER li1 ;
        RECT 2216.165 216.050 2216.340 216.220 ;
        RECT 2213.715 215.880 2216.340 216.050 ;
        RECT 2216.165 215.680 2216.340 215.880 ;
      LAYER li1 ;
        RECT 2219.195 215.680 2219.450 216.220 ;
      LAYER li1 ;
        RECT 2222.145 216.050 2222.320 216.220 ;
        RECT 2219.695 215.880 2222.320 216.050 ;
        RECT 2222.145 215.680 2222.320 215.880 ;
      LAYER li1 ;
        RECT 2225.175 215.680 2225.430 216.220 ;
      LAYER li1 ;
        RECT 2228.125 216.050 2228.300 216.220 ;
        RECT 2225.675 215.880 2228.300 216.050 ;
        RECT 2228.125 215.680 2228.300 215.880 ;
      LAYER li1 ;
        RECT 2231.155 215.680 2231.410 216.220 ;
      LAYER li1 ;
        RECT 2234.105 216.050 2234.280 216.220 ;
        RECT 2231.655 215.880 2234.280 216.050 ;
        RECT 2234.105 215.680 2234.280 215.880 ;
      LAYER li1 ;
        RECT 2237.135 215.680 2237.390 216.220 ;
      LAYER li1 ;
        RECT 2240.085 216.050 2240.260 216.220 ;
        RECT 2237.635 215.880 2240.260 216.050 ;
        RECT 2240.085 215.680 2240.260 215.880 ;
      LAYER li1 ;
        RECT 2243.115 215.680 2243.370 216.220 ;
      LAYER li1 ;
        RECT 2246.065 216.050 2246.240 216.220 ;
        RECT 2243.615 215.880 2246.240 216.050 ;
        RECT 2246.065 215.680 2246.240 215.880 ;
      LAYER li1 ;
        RECT 2249.095 215.680 2249.350 216.220 ;
      LAYER li1 ;
        RECT 2252.045 216.050 2252.220 216.220 ;
        RECT 2249.595 215.880 2252.220 216.050 ;
        RECT 2252.045 215.680 2252.220 215.880 ;
      LAYER li1 ;
        RECT 2255.075 215.680 2255.330 216.220 ;
      LAYER li1 ;
        RECT 2258.025 216.050 2258.200 216.220 ;
        RECT 2255.575 215.880 2258.200 216.050 ;
        RECT 2258.025 215.680 2258.200 215.880 ;
      LAYER li1 ;
        RECT 2261.055 215.680 2261.310 216.220 ;
      LAYER li1 ;
        RECT 2264.005 216.050 2264.180 216.220 ;
        RECT 2261.555 215.880 2264.180 216.050 ;
        RECT 2264.005 215.680 2264.180 215.880 ;
      LAYER li1 ;
        RECT 2267.035 215.680 2267.290 216.220 ;
      LAYER li1 ;
        RECT 2269.985 216.050 2270.160 216.220 ;
        RECT 2267.535 215.880 2270.160 216.050 ;
        RECT 2269.985 215.680 2270.160 215.880 ;
        RECT 669.085 214.490 669.375 215.655 ;
        RECT 669.935 214.490 670.265 215.640 ;
      LAYER li1 ;
        RECT 670.435 215.510 673.125 215.680 ;
      LAYER li1 ;
        RECT 673.385 215.510 674.885 215.680 ;
      LAYER li1 ;
        RECT 670.435 214.660 670.605 215.510 ;
      LAYER li1 ;
        RECT 670.775 214.490 671.105 215.290 ;
      LAYER li1 ;
        RECT 671.275 214.660 671.445 215.510 ;
      LAYER li1 ;
        RECT 671.615 214.490 671.945 215.290 ;
      LAYER li1 ;
        RECT 672.115 214.660 672.285 215.510 ;
      LAYER li1 ;
        RECT 672.455 214.490 672.785 215.290 ;
      LAYER li1 ;
        RECT 672.955 214.660 673.125 215.510 ;
      LAYER li1 ;
        RECT 673.375 214.490 673.545 215.290 ;
        RECT 673.715 214.660 674.045 215.510 ;
        RECT 674.215 214.490 674.385 215.290 ;
        RECT 674.555 214.660 674.885 215.510 ;
        RECT 675.065 214.490 675.355 215.655 ;
        RECT 675.915 214.490 676.245 215.640 ;
      LAYER li1 ;
        RECT 676.415 215.510 679.105 215.680 ;
      LAYER li1 ;
        RECT 679.365 215.510 680.865 215.680 ;
      LAYER li1 ;
        RECT 676.415 214.660 676.585 215.510 ;
      LAYER li1 ;
        RECT 676.755 214.490 677.085 215.290 ;
      LAYER li1 ;
        RECT 677.255 214.660 677.425 215.510 ;
      LAYER li1 ;
        RECT 677.595 214.490 677.925 215.290 ;
      LAYER li1 ;
        RECT 678.095 214.660 678.265 215.510 ;
      LAYER li1 ;
        RECT 678.435 214.490 678.765 215.290 ;
      LAYER li1 ;
        RECT 678.935 214.660 679.105 215.510 ;
      LAYER li1 ;
        RECT 679.355 214.490 679.525 215.290 ;
        RECT 679.695 214.660 680.025 215.510 ;
        RECT 680.195 214.490 680.365 215.290 ;
        RECT 680.535 214.660 680.865 215.510 ;
        RECT 681.045 214.490 681.335 215.655 ;
        RECT 681.895 214.490 682.225 215.640 ;
      LAYER li1 ;
        RECT 682.395 215.510 685.085 215.680 ;
      LAYER li1 ;
        RECT 685.345 215.510 686.845 215.680 ;
      LAYER li1 ;
        RECT 682.395 214.660 682.565 215.510 ;
      LAYER li1 ;
        RECT 682.735 214.490 683.065 215.290 ;
      LAYER li1 ;
        RECT 683.235 214.660 683.405 215.510 ;
      LAYER li1 ;
        RECT 683.575 214.490 683.905 215.290 ;
      LAYER li1 ;
        RECT 684.075 214.660 684.245 215.510 ;
      LAYER li1 ;
        RECT 684.415 214.490 684.745 215.290 ;
      LAYER li1 ;
        RECT 684.915 214.660 685.085 215.510 ;
      LAYER li1 ;
        RECT 685.335 214.490 685.505 215.290 ;
        RECT 685.675 214.660 686.005 215.510 ;
        RECT 686.175 214.490 686.345 215.290 ;
        RECT 686.515 214.660 686.845 215.510 ;
        RECT 687.025 214.490 687.315 215.655 ;
        RECT 687.875 214.490 688.205 215.640 ;
      LAYER li1 ;
        RECT 688.375 215.510 691.065 215.680 ;
      LAYER li1 ;
        RECT 691.325 215.510 692.825 215.680 ;
      LAYER li1 ;
        RECT 688.375 214.660 688.545 215.510 ;
      LAYER li1 ;
        RECT 688.715 214.490 689.045 215.290 ;
      LAYER li1 ;
        RECT 689.215 214.660 689.385 215.510 ;
      LAYER li1 ;
        RECT 689.555 214.490 689.885 215.290 ;
      LAYER li1 ;
        RECT 690.055 214.660 690.225 215.510 ;
      LAYER li1 ;
        RECT 690.395 214.490 690.725 215.290 ;
      LAYER li1 ;
        RECT 690.895 214.660 691.065 215.510 ;
      LAYER li1 ;
        RECT 691.315 214.490 691.485 215.290 ;
        RECT 691.655 214.660 691.985 215.510 ;
        RECT 692.155 214.490 692.325 215.290 ;
        RECT 692.495 214.660 692.825 215.510 ;
        RECT 693.005 214.490 693.295 215.655 ;
        RECT 693.855 214.490 694.185 215.640 ;
      LAYER li1 ;
        RECT 694.355 215.510 697.045 215.680 ;
      LAYER li1 ;
        RECT 697.305 215.510 698.805 215.680 ;
      LAYER li1 ;
        RECT 694.355 214.660 694.525 215.510 ;
      LAYER li1 ;
        RECT 694.695 214.490 695.025 215.290 ;
      LAYER li1 ;
        RECT 695.195 214.660 695.365 215.510 ;
      LAYER li1 ;
        RECT 695.535 214.490 695.865 215.290 ;
      LAYER li1 ;
        RECT 696.035 214.660 696.205 215.510 ;
      LAYER li1 ;
        RECT 696.375 214.490 696.705 215.290 ;
      LAYER li1 ;
        RECT 696.875 214.660 697.045 215.510 ;
      LAYER li1 ;
        RECT 697.295 214.490 697.465 215.290 ;
        RECT 697.635 214.660 697.965 215.510 ;
        RECT 698.135 214.490 698.305 215.290 ;
        RECT 698.475 214.660 698.805 215.510 ;
        RECT 698.985 214.490 699.275 215.655 ;
        RECT 699.835 214.490 700.165 215.640 ;
      LAYER li1 ;
        RECT 700.335 215.510 703.025 215.680 ;
      LAYER li1 ;
        RECT 703.285 215.510 704.785 215.680 ;
      LAYER li1 ;
        RECT 700.335 214.660 700.505 215.510 ;
      LAYER li1 ;
        RECT 700.675 214.490 701.005 215.290 ;
      LAYER li1 ;
        RECT 701.175 214.660 701.345 215.510 ;
      LAYER li1 ;
        RECT 701.515 214.490 701.845 215.290 ;
      LAYER li1 ;
        RECT 702.015 214.660 702.185 215.510 ;
      LAYER li1 ;
        RECT 702.355 214.490 702.685 215.290 ;
      LAYER li1 ;
        RECT 702.855 214.660 703.025 215.510 ;
      LAYER li1 ;
        RECT 703.275 214.490 703.445 215.290 ;
        RECT 703.615 214.660 703.945 215.510 ;
        RECT 704.115 214.490 704.285 215.290 ;
        RECT 704.455 214.660 704.785 215.510 ;
        RECT 704.965 214.490 705.255 215.655 ;
        RECT 705.815 214.490 706.145 215.640 ;
      LAYER li1 ;
        RECT 706.315 215.510 709.005 215.680 ;
      LAYER li1 ;
        RECT 709.265 215.510 710.765 215.680 ;
      LAYER li1 ;
        RECT 706.315 214.660 706.485 215.510 ;
      LAYER li1 ;
        RECT 706.655 214.490 706.985 215.290 ;
      LAYER li1 ;
        RECT 707.155 214.660 707.325 215.510 ;
      LAYER li1 ;
        RECT 707.495 214.490 707.825 215.290 ;
      LAYER li1 ;
        RECT 707.995 214.660 708.165 215.510 ;
      LAYER li1 ;
        RECT 708.335 214.490 708.665 215.290 ;
      LAYER li1 ;
        RECT 708.835 214.660 709.005 215.510 ;
      LAYER li1 ;
        RECT 709.255 214.490 709.425 215.290 ;
        RECT 709.595 214.660 709.925 215.510 ;
        RECT 710.095 214.490 710.265 215.290 ;
        RECT 710.435 214.660 710.765 215.510 ;
        RECT 710.945 214.490 711.235 215.655 ;
        RECT 711.795 214.490 712.125 215.640 ;
      LAYER li1 ;
        RECT 712.295 215.510 714.985 215.680 ;
      LAYER li1 ;
        RECT 715.245 215.510 716.745 215.680 ;
      LAYER li1 ;
        RECT 712.295 214.660 712.465 215.510 ;
      LAYER li1 ;
        RECT 712.635 214.490 712.965 215.290 ;
      LAYER li1 ;
        RECT 713.135 214.660 713.305 215.510 ;
      LAYER li1 ;
        RECT 713.475 214.490 713.805 215.290 ;
      LAYER li1 ;
        RECT 713.975 214.660 714.145 215.510 ;
      LAYER li1 ;
        RECT 714.315 214.490 714.645 215.290 ;
      LAYER li1 ;
        RECT 714.815 214.660 714.985 215.510 ;
      LAYER li1 ;
        RECT 715.235 214.490 715.405 215.290 ;
        RECT 715.575 214.660 715.905 215.510 ;
        RECT 716.075 214.490 716.245 215.290 ;
        RECT 716.415 214.660 716.745 215.510 ;
        RECT 716.925 214.490 717.215 215.655 ;
        RECT 717.775 214.490 718.105 215.640 ;
      LAYER li1 ;
        RECT 718.275 215.510 720.965 215.680 ;
      LAYER li1 ;
        RECT 721.225 215.510 722.725 215.680 ;
      LAYER li1 ;
        RECT 718.275 214.660 718.445 215.510 ;
      LAYER li1 ;
        RECT 718.615 214.490 718.945 215.290 ;
      LAYER li1 ;
        RECT 719.115 214.660 719.285 215.510 ;
      LAYER li1 ;
        RECT 719.455 214.490 719.785 215.290 ;
      LAYER li1 ;
        RECT 719.955 214.660 720.125 215.510 ;
      LAYER li1 ;
        RECT 720.295 214.490 720.625 215.290 ;
      LAYER li1 ;
        RECT 720.795 214.660 720.965 215.510 ;
      LAYER li1 ;
        RECT 721.215 214.490 721.385 215.290 ;
        RECT 721.555 214.660 721.885 215.510 ;
        RECT 722.055 214.490 722.225 215.290 ;
        RECT 722.395 214.660 722.725 215.510 ;
        RECT 722.905 214.490 723.195 215.655 ;
        RECT 723.755 214.490 724.085 215.640 ;
      LAYER li1 ;
        RECT 724.255 215.510 726.945 215.680 ;
      LAYER li1 ;
        RECT 727.205 215.510 728.705 215.680 ;
      LAYER li1 ;
        RECT 724.255 214.660 724.425 215.510 ;
      LAYER li1 ;
        RECT 724.595 214.490 724.925 215.290 ;
      LAYER li1 ;
        RECT 725.095 214.660 725.265 215.510 ;
      LAYER li1 ;
        RECT 725.435 214.490 725.765 215.290 ;
      LAYER li1 ;
        RECT 725.935 214.660 726.105 215.510 ;
      LAYER li1 ;
        RECT 726.275 214.490 726.605 215.290 ;
      LAYER li1 ;
        RECT 726.775 214.660 726.945 215.510 ;
      LAYER li1 ;
        RECT 727.195 214.490 727.365 215.290 ;
        RECT 727.535 214.660 727.865 215.510 ;
        RECT 728.035 214.490 728.205 215.290 ;
        RECT 728.375 214.660 728.705 215.510 ;
        RECT 728.885 214.490 729.175 215.655 ;
        RECT 729.735 214.490 730.065 215.640 ;
      LAYER li1 ;
        RECT 730.235 215.510 732.925 215.680 ;
      LAYER li1 ;
        RECT 733.185 215.510 734.685 215.680 ;
      LAYER li1 ;
        RECT 730.235 214.660 730.405 215.510 ;
      LAYER li1 ;
        RECT 730.575 214.490 730.905 215.290 ;
      LAYER li1 ;
        RECT 731.075 214.660 731.245 215.510 ;
      LAYER li1 ;
        RECT 731.415 214.490 731.745 215.290 ;
      LAYER li1 ;
        RECT 731.915 214.660 732.085 215.510 ;
      LAYER li1 ;
        RECT 732.255 214.490 732.585 215.290 ;
      LAYER li1 ;
        RECT 732.755 214.660 732.925 215.510 ;
      LAYER li1 ;
        RECT 733.175 214.490 733.345 215.290 ;
        RECT 733.515 214.660 733.845 215.510 ;
        RECT 734.015 214.490 734.185 215.290 ;
        RECT 734.355 214.660 734.685 215.510 ;
        RECT 734.865 214.490 735.155 215.655 ;
        RECT 735.715 214.490 736.045 215.640 ;
      LAYER li1 ;
        RECT 736.215 215.510 738.905 215.680 ;
      LAYER li1 ;
        RECT 739.165 215.510 740.665 215.680 ;
      LAYER li1 ;
        RECT 736.215 214.660 736.385 215.510 ;
      LAYER li1 ;
        RECT 736.555 214.490 736.885 215.290 ;
      LAYER li1 ;
        RECT 737.055 214.660 737.225 215.510 ;
      LAYER li1 ;
        RECT 737.395 214.490 737.725 215.290 ;
      LAYER li1 ;
        RECT 737.895 214.660 738.065 215.510 ;
      LAYER li1 ;
        RECT 738.235 214.490 738.565 215.290 ;
      LAYER li1 ;
        RECT 738.735 214.660 738.905 215.510 ;
      LAYER li1 ;
        RECT 739.155 214.490 739.325 215.290 ;
        RECT 739.495 214.660 739.825 215.510 ;
        RECT 739.995 214.490 740.165 215.290 ;
        RECT 740.335 214.660 740.665 215.510 ;
        RECT 740.845 214.490 741.135 215.655 ;
        RECT 741.695 214.490 742.025 215.640 ;
      LAYER li1 ;
        RECT 742.195 215.510 744.885 215.680 ;
      LAYER li1 ;
        RECT 745.145 215.510 746.645 215.680 ;
      LAYER li1 ;
        RECT 742.195 214.660 742.365 215.510 ;
      LAYER li1 ;
        RECT 742.535 214.490 742.865 215.290 ;
      LAYER li1 ;
        RECT 743.035 214.660 743.205 215.510 ;
      LAYER li1 ;
        RECT 743.375 214.490 743.705 215.290 ;
      LAYER li1 ;
        RECT 743.875 214.660 744.045 215.510 ;
      LAYER li1 ;
        RECT 744.215 214.490 744.545 215.290 ;
      LAYER li1 ;
        RECT 744.715 214.660 744.885 215.510 ;
      LAYER li1 ;
        RECT 745.135 214.490 745.305 215.290 ;
        RECT 745.475 214.660 745.805 215.510 ;
        RECT 745.975 214.490 746.145 215.290 ;
        RECT 746.315 214.660 746.645 215.510 ;
        RECT 746.825 214.490 747.115 215.655 ;
        RECT 747.675 214.490 748.005 215.640 ;
      LAYER li1 ;
        RECT 748.175 215.510 750.865 215.680 ;
      LAYER li1 ;
        RECT 751.125 215.510 752.625 215.680 ;
      LAYER li1 ;
        RECT 748.175 214.660 748.345 215.510 ;
      LAYER li1 ;
        RECT 748.515 214.490 748.845 215.290 ;
      LAYER li1 ;
        RECT 749.015 214.660 749.185 215.510 ;
      LAYER li1 ;
        RECT 749.355 214.490 749.685 215.290 ;
      LAYER li1 ;
        RECT 749.855 214.660 750.025 215.510 ;
      LAYER li1 ;
        RECT 750.195 214.490 750.525 215.290 ;
      LAYER li1 ;
        RECT 750.695 214.660 750.865 215.510 ;
      LAYER li1 ;
        RECT 751.115 214.490 751.285 215.290 ;
        RECT 751.455 214.660 751.785 215.510 ;
        RECT 751.955 214.490 752.125 215.290 ;
        RECT 752.295 214.660 752.625 215.510 ;
        RECT 752.805 214.490 753.095 215.655 ;
        RECT 753.655 214.490 753.985 215.640 ;
      LAYER li1 ;
        RECT 754.155 215.510 756.845 215.680 ;
      LAYER li1 ;
        RECT 757.105 215.510 758.605 215.680 ;
      LAYER li1 ;
        RECT 754.155 214.660 754.325 215.510 ;
      LAYER li1 ;
        RECT 754.495 214.490 754.825 215.290 ;
      LAYER li1 ;
        RECT 754.995 214.660 755.165 215.510 ;
      LAYER li1 ;
        RECT 755.335 214.490 755.665 215.290 ;
      LAYER li1 ;
        RECT 755.835 214.660 756.005 215.510 ;
      LAYER li1 ;
        RECT 756.175 214.490 756.505 215.290 ;
      LAYER li1 ;
        RECT 756.675 214.660 756.845 215.510 ;
      LAYER li1 ;
        RECT 757.095 214.490 757.265 215.290 ;
        RECT 757.435 214.660 757.765 215.510 ;
        RECT 757.935 214.490 758.105 215.290 ;
        RECT 758.275 214.660 758.605 215.510 ;
        RECT 758.785 214.490 759.075 215.655 ;
        RECT 759.635 214.490 759.965 215.640 ;
        RECT 763.085 215.510 764.585 215.680 ;
        RECT 760.475 214.490 760.805 215.290 ;
        RECT 761.315 214.490 761.645 215.290 ;
        RECT 762.155 214.490 762.485 215.290 ;
        RECT 763.075 214.490 763.245 215.290 ;
        RECT 763.415 214.660 763.745 215.510 ;
        RECT 763.915 214.490 764.085 215.290 ;
        RECT 764.255 214.660 764.585 215.510 ;
        RECT 764.765 214.490 765.055 215.655 ;
        RECT 765.615 214.490 765.945 215.640 ;
        RECT 769.065 215.510 770.565 215.680 ;
        RECT 766.455 214.490 766.785 215.290 ;
        RECT 767.295 214.490 767.625 215.290 ;
        RECT 768.135 214.490 768.465 215.290 ;
        RECT 769.055 214.490 769.225 215.290 ;
        RECT 769.395 214.660 769.725 215.510 ;
        RECT 769.895 214.490 770.065 215.290 ;
        RECT 770.235 214.660 770.565 215.510 ;
        RECT 770.745 214.490 771.035 215.655 ;
        RECT 771.595 214.490 771.925 215.640 ;
        RECT 775.045 215.510 776.545 215.680 ;
        RECT 772.435 214.490 772.765 215.290 ;
        RECT 773.275 214.490 773.605 215.290 ;
        RECT 774.115 214.490 774.445 215.290 ;
        RECT 775.035 214.490 775.205 215.290 ;
        RECT 775.375 214.660 775.705 215.510 ;
        RECT 775.875 214.490 776.045 215.290 ;
        RECT 776.215 214.660 776.545 215.510 ;
        RECT 776.725 214.490 777.015 215.655 ;
        RECT 777.575 214.490 777.905 215.640 ;
        RECT 781.025 215.510 782.525 215.680 ;
        RECT 778.415 214.490 778.745 215.290 ;
        RECT 779.255 214.490 779.585 215.290 ;
        RECT 780.095 214.490 780.425 215.290 ;
        RECT 781.015 214.490 781.185 215.290 ;
        RECT 781.355 214.660 781.685 215.510 ;
        RECT 781.855 214.490 782.025 215.290 ;
        RECT 782.195 214.660 782.525 215.510 ;
        RECT 782.705 214.490 782.995 215.655 ;
        RECT 783.555 214.490 783.885 215.640 ;
        RECT 787.005 215.510 788.505 215.680 ;
        RECT 784.395 214.490 784.725 215.290 ;
        RECT 785.235 214.490 785.565 215.290 ;
        RECT 786.075 214.490 786.405 215.290 ;
        RECT 786.995 214.490 787.165 215.290 ;
        RECT 787.335 214.660 787.665 215.510 ;
        RECT 787.835 214.490 788.005 215.290 ;
        RECT 788.175 214.660 788.505 215.510 ;
        RECT 788.685 214.490 788.975 215.655 ;
        RECT 789.535 214.490 789.865 215.640 ;
        RECT 792.985 215.510 794.485 215.680 ;
        RECT 790.375 214.490 790.705 215.290 ;
        RECT 791.215 214.490 791.545 215.290 ;
        RECT 792.055 214.490 792.385 215.290 ;
        RECT 792.975 214.490 793.145 215.290 ;
        RECT 793.315 214.660 793.645 215.510 ;
        RECT 793.815 214.490 793.985 215.290 ;
        RECT 794.155 214.660 794.485 215.510 ;
        RECT 794.665 214.490 794.955 215.655 ;
        RECT 2146.085 214.490 2146.375 215.655 ;
        RECT 2146.935 214.490 2147.265 215.640 ;
      LAYER li1 ;
        RECT 2147.435 215.510 2150.125 215.680 ;
      LAYER li1 ;
        RECT 2150.385 215.510 2151.885 215.680 ;
      LAYER li1 ;
        RECT 2147.435 214.660 2147.605 215.510 ;
      LAYER li1 ;
        RECT 2147.775 214.490 2148.105 215.290 ;
      LAYER li1 ;
        RECT 2148.275 214.660 2148.445 215.510 ;
      LAYER li1 ;
        RECT 2148.615 214.490 2148.945 215.290 ;
      LAYER li1 ;
        RECT 2149.115 214.660 2149.285 215.510 ;
      LAYER li1 ;
        RECT 2149.455 214.490 2149.785 215.290 ;
      LAYER li1 ;
        RECT 2149.955 214.660 2150.125 215.510 ;
      LAYER li1 ;
        RECT 2150.375 214.490 2150.545 215.290 ;
        RECT 2150.715 214.660 2151.045 215.510 ;
        RECT 2151.215 214.490 2151.385 215.290 ;
        RECT 2151.555 214.660 2151.885 215.510 ;
        RECT 2152.065 214.490 2152.355 215.655 ;
        RECT 2152.915 214.490 2153.245 215.640 ;
      LAYER li1 ;
        RECT 2153.415 215.510 2156.105 215.680 ;
      LAYER li1 ;
        RECT 2156.365 215.510 2157.865 215.680 ;
      LAYER li1 ;
        RECT 2153.415 214.660 2153.585 215.510 ;
      LAYER li1 ;
        RECT 2153.755 214.490 2154.085 215.290 ;
      LAYER li1 ;
        RECT 2154.255 214.660 2154.425 215.510 ;
      LAYER li1 ;
        RECT 2154.595 214.490 2154.925 215.290 ;
      LAYER li1 ;
        RECT 2155.095 214.660 2155.265 215.510 ;
      LAYER li1 ;
        RECT 2155.435 214.490 2155.765 215.290 ;
      LAYER li1 ;
        RECT 2155.935 214.660 2156.105 215.510 ;
      LAYER li1 ;
        RECT 2156.355 214.490 2156.525 215.290 ;
        RECT 2156.695 214.660 2157.025 215.510 ;
        RECT 2157.195 214.490 2157.365 215.290 ;
        RECT 2157.535 214.660 2157.865 215.510 ;
        RECT 2158.045 214.490 2158.335 215.655 ;
        RECT 2158.895 214.490 2159.225 215.640 ;
      LAYER li1 ;
        RECT 2159.395 215.510 2162.085 215.680 ;
      LAYER li1 ;
        RECT 2162.345 215.510 2163.845 215.680 ;
      LAYER li1 ;
        RECT 2159.395 214.660 2159.565 215.510 ;
      LAYER li1 ;
        RECT 2159.735 214.490 2160.065 215.290 ;
      LAYER li1 ;
        RECT 2160.235 214.660 2160.405 215.510 ;
      LAYER li1 ;
        RECT 2160.575 214.490 2160.905 215.290 ;
      LAYER li1 ;
        RECT 2161.075 214.660 2161.245 215.510 ;
      LAYER li1 ;
        RECT 2161.415 214.490 2161.745 215.290 ;
      LAYER li1 ;
        RECT 2161.915 214.660 2162.085 215.510 ;
      LAYER li1 ;
        RECT 2162.335 214.490 2162.505 215.290 ;
        RECT 2162.675 214.660 2163.005 215.510 ;
        RECT 2163.175 214.490 2163.345 215.290 ;
        RECT 2163.515 214.660 2163.845 215.510 ;
        RECT 2164.025 214.490 2164.315 215.655 ;
        RECT 2164.875 214.490 2165.205 215.640 ;
      LAYER li1 ;
        RECT 2165.375 215.510 2168.065 215.680 ;
      LAYER li1 ;
        RECT 2168.325 215.510 2169.825 215.680 ;
      LAYER li1 ;
        RECT 2165.375 214.660 2165.545 215.510 ;
      LAYER li1 ;
        RECT 2165.715 214.490 2166.045 215.290 ;
      LAYER li1 ;
        RECT 2166.215 214.660 2166.385 215.510 ;
      LAYER li1 ;
        RECT 2166.555 214.490 2166.885 215.290 ;
      LAYER li1 ;
        RECT 2167.055 214.660 2167.225 215.510 ;
      LAYER li1 ;
        RECT 2167.395 214.490 2167.725 215.290 ;
      LAYER li1 ;
        RECT 2167.895 214.660 2168.065 215.510 ;
      LAYER li1 ;
        RECT 2168.315 214.490 2168.485 215.290 ;
        RECT 2168.655 214.660 2168.985 215.510 ;
        RECT 2169.155 214.490 2169.325 215.290 ;
        RECT 2169.495 214.660 2169.825 215.510 ;
        RECT 2170.005 214.490 2170.295 215.655 ;
        RECT 2170.855 214.490 2171.185 215.640 ;
      LAYER li1 ;
        RECT 2171.355 215.510 2174.045 215.680 ;
      LAYER li1 ;
        RECT 2174.305 215.510 2175.805 215.680 ;
      LAYER li1 ;
        RECT 2171.355 214.660 2171.525 215.510 ;
      LAYER li1 ;
        RECT 2171.695 214.490 2172.025 215.290 ;
      LAYER li1 ;
        RECT 2172.195 214.660 2172.365 215.510 ;
      LAYER li1 ;
        RECT 2172.535 214.490 2172.865 215.290 ;
      LAYER li1 ;
        RECT 2173.035 214.660 2173.205 215.510 ;
      LAYER li1 ;
        RECT 2173.375 214.490 2173.705 215.290 ;
      LAYER li1 ;
        RECT 2173.875 214.660 2174.045 215.510 ;
      LAYER li1 ;
        RECT 2174.295 214.490 2174.465 215.290 ;
        RECT 2174.635 214.660 2174.965 215.510 ;
        RECT 2175.135 214.490 2175.305 215.290 ;
        RECT 2175.475 214.660 2175.805 215.510 ;
        RECT 2175.985 214.490 2176.275 215.655 ;
        RECT 2176.835 214.490 2177.165 215.640 ;
      LAYER li1 ;
        RECT 2177.335 215.510 2180.025 215.680 ;
      LAYER li1 ;
        RECT 2180.285 215.510 2181.785 215.680 ;
      LAYER li1 ;
        RECT 2177.335 214.660 2177.505 215.510 ;
      LAYER li1 ;
        RECT 2177.675 214.490 2178.005 215.290 ;
      LAYER li1 ;
        RECT 2178.175 214.660 2178.345 215.510 ;
      LAYER li1 ;
        RECT 2178.515 214.490 2178.845 215.290 ;
      LAYER li1 ;
        RECT 2179.015 214.660 2179.185 215.510 ;
      LAYER li1 ;
        RECT 2179.355 214.490 2179.685 215.290 ;
      LAYER li1 ;
        RECT 2179.855 214.660 2180.025 215.510 ;
      LAYER li1 ;
        RECT 2180.275 214.490 2180.445 215.290 ;
        RECT 2180.615 214.660 2180.945 215.510 ;
        RECT 2181.115 214.490 2181.285 215.290 ;
        RECT 2181.455 214.660 2181.785 215.510 ;
        RECT 2181.965 214.490 2182.255 215.655 ;
        RECT 2182.815 214.490 2183.145 215.640 ;
      LAYER li1 ;
        RECT 2183.315 215.510 2186.005 215.680 ;
      LAYER li1 ;
        RECT 2186.265 215.510 2187.765 215.680 ;
      LAYER li1 ;
        RECT 2183.315 214.660 2183.485 215.510 ;
      LAYER li1 ;
        RECT 2183.655 214.490 2183.985 215.290 ;
      LAYER li1 ;
        RECT 2184.155 214.660 2184.325 215.510 ;
      LAYER li1 ;
        RECT 2184.495 214.490 2184.825 215.290 ;
      LAYER li1 ;
        RECT 2184.995 214.660 2185.165 215.510 ;
      LAYER li1 ;
        RECT 2185.335 214.490 2185.665 215.290 ;
      LAYER li1 ;
        RECT 2185.835 214.660 2186.005 215.510 ;
      LAYER li1 ;
        RECT 2186.255 214.490 2186.425 215.290 ;
        RECT 2186.595 214.660 2186.925 215.510 ;
        RECT 2187.095 214.490 2187.265 215.290 ;
        RECT 2187.435 214.660 2187.765 215.510 ;
        RECT 2187.945 214.490 2188.235 215.655 ;
        RECT 2188.795 214.490 2189.125 215.640 ;
      LAYER li1 ;
        RECT 2189.295 215.510 2191.985 215.680 ;
      LAYER li1 ;
        RECT 2192.245 215.510 2193.745 215.680 ;
      LAYER li1 ;
        RECT 2189.295 214.660 2189.465 215.510 ;
      LAYER li1 ;
        RECT 2189.635 214.490 2189.965 215.290 ;
      LAYER li1 ;
        RECT 2190.135 214.660 2190.305 215.510 ;
      LAYER li1 ;
        RECT 2190.475 214.490 2190.805 215.290 ;
      LAYER li1 ;
        RECT 2190.975 214.660 2191.145 215.510 ;
      LAYER li1 ;
        RECT 2191.315 214.490 2191.645 215.290 ;
      LAYER li1 ;
        RECT 2191.815 214.660 2191.985 215.510 ;
      LAYER li1 ;
        RECT 2192.235 214.490 2192.405 215.290 ;
        RECT 2192.575 214.660 2192.905 215.510 ;
        RECT 2193.075 214.490 2193.245 215.290 ;
        RECT 2193.415 214.660 2193.745 215.510 ;
        RECT 2193.925 214.490 2194.215 215.655 ;
        RECT 2194.775 214.490 2195.105 215.640 ;
      LAYER li1 ;
        RECT 2195.275 215.510 2197.965 215.680 ;
      LAYER li1 ;
        RECT 2198.225 215.510 2199.725 215.680 ;
      LAYER li1 ;
        RECT 2195.275 214.660 2195.445 215.510 ;
      LAYER li1 ;
        RECT 2195.615 214.490 2195.945 215.290 ;
      LAYER li1 ;
        RECT 2196.115 214.660 2196.285 215.510 ;
      LAYER li1 ;
        RECT 2196.455 214.490 2196.785 215.290 ;
      LAYER li1 ;
        RECT 2196.955 214.660 2197.125 215.510 ;
      LAYER li1 ;
        RECT 2197.295 214.490 2197.625 215.290 ;
      LAYER li1 ;
        RECT 2197.795 214.660 2197.965 215.510 ;
      LAYER li1 ;
        RECT 2198.215 214.490 2198.385 215.290 ;
        RECT 2198.555 214.660 2198.885 215.510 ;
        RECT 2199.055 214.490 2199.225 215.290 ;
        RECT 2199.395 214.660 2199.725 215.510 ;
        RECT 2199.905 214.490 2200.195 215.655 ;
        RECT 2200.755 214.490 2201.085 215.640 ;
      LAYER li1 ;
        RECT 2201.255 215.510 2203.945 215.680 ;
      LAYER li1 ;
        RECT 2204.205 215.510 2205.705 215.680 ;
      LAYER li1 ;
        RECT 2201.255 214.660 2201.425 215.510 ;
      LAYER li1 ;
        RECT 2201.595 214.490 2201.925 215.290 ;
      LAYER li1 ;
        RECT 2202.095 214.660 2202.265 215.510 ;
      LAYER li1 ;
        RECT 2202.435 214.490 2202.765 215.290 ;
      LAYER li1 ;
        RECT 2202.935 214.660 2203.105 215.510 ;
      LAYER li1 ;
        RECT 2203.275 214.490 2203.605 215.290 ;
      LAYER li1 ;
        RECT 2203.775 214.660 2203.945 215.510 ;
      LAYER li1 ;
        RECT 2204.195 214.490 2204.365 215.290 ;
        RECT 2204.535 214.660 2204.865 215.510 ;
        RECT 2205.035 214.490 2205.205 215.290 ;
        RECT 2205.375 214.660 2205.705 215.510 ;
        RECT 2205.885 214.490 2206.175 215.655 ;
        RECT 2206.735 214.490 2207.065 215.640 ;
      LAYER li1 ;
        RECT 2207.235 215.510 2209.925 215.680 ;
      LAYER li1 ;
        RECT 2210.185 215.510 2211.685 215.680 ;
      LAYER li1 ;
        RECT 2207.235 214.660 2207.405 215.510 ;
      LAYER li1 ;
        RECT 2207.575 214.490 2207.905 215.290 ;
      LAYER li1 ;
        RECT 2208.075 214.660 2208.245 215.510 ;
      LAYER li1 ;
        RECT 2208.415 214.490 2208.745 215.290 ;
      LAYER li1 ;
        RECT 2208.915 214.660 2209.085 215.510 ;
      LAYER li1 ;
        RECT 2209.255 214.490 2209.585 215.290 ;
      LAYER li1 ;
        RECT 2209.755 214.660 2209.925 215.510 ;
      LAYER li1 ;
        RECT 2210.175 214.490 2210.345 215.290 ;
        RECT 2210.515 214.660 2210.845 215.510 ;
        RECT 2211.015 214.490 2211.185 215.290 ;
        RECT 2211.355 214.660 2211.685 215.510 ;
        RECT 2211.865 214.490 2212.155 215.655 ;
        RECT 2212.715 214.490 2213.045 215.640 ;
      LAYER li1 ;
        RECT 2213.215 215.510 2215.905 215.680 ;
      LAYER li1 ;
        RECT 2216.165 215.510 2217.665 215.680 ;
      LAYER li1 ;
        RECT 2213.215 214.660 2213.385 215.510 ;
      LAYER li1 ;
        RECT 2213.555 214.490 2213.885 215.290 ;
      LAYER li1 ;
        RECT 2214.055 214.660 2214.225 215.510 ;
      LAYER li1 ;
        RECT 2214.395 214.490 2214.725 215.290 ;
      LAYER li1 ;
        RECT 2214.895 214.660 2215.065 215.510 ;
      LAYER li1 ;
        RECT 2215.235 214.490 2215.565 215.290 ;
      LAYER li1 ;
        RECT 2215.735 214.660 2215.905 215.510 ;
      LAYER li1 ;
        RECT 2216.155 214.490 2216.325 215.290 ;
        RECT 2216.495 214.660 2216.825 215.510 ;
        RECT 2216.995 214.490 2217.165 215.290 ;
        RECT 2217.335 214.660 2217.665 215.510 ;
        RECT 2217.845 214.490 2218.135 215.655 ;
        RECT 2218.695 214.490 2219.025 215.640 ;
      LAYER li1 ;
        RECT 2219.195 215.510 2221.885 215.680 ;
      LAYER li1 ;
        RECT 2222.145 215.510 2223.645 215.680 ;
      LAYER li1 ;
        RECT 2219.195 214.660 2219.365 215.510 ;
      LAYER li1 ;
        RECT 2219.535 214.490 2219.865 215.290 ;
      LAYER li1 ;
        RECT 2220.035 214.660 2220.205 215.510 ;
      LAYER li1 ;
        RECT 2220.375 214.490 2220.705 215.290 ;
      LAYER li1 ;
        RECT 2220.875 214.660 2221.045 215.510 ;
      LAYER li1 ;
        RECT 2221.215 214.490 2221.545 215.290 ;
      LAYER li1 ;
        RECT 2221.715 214.660 2221.885 215.510 ;
      LAYER li1 ;
        RECT 2222.135 214.490 2222.305 215.290 ;
        RECT 2222.475 214.660 2222.805 215.510 ;
        RECT 2222.975 214.490 2223.145 215.290 ;
        RECT 2223.315 214.660 2223.645 215.510 ;
        RECT 2223.825 214.490 2224.115 215.655 ;
        RECT 2224.675 214.490 2225.005 215.640 ;
      LAYER li1 ;
        RECT 2225.175 215.510 2227.865 215.680 ;
      LAYER li1 ;
        RECT 2228.125 215.510 2229.625 215.680 ;
      LAYER li1 ;
        RECT 2225.175 214.660 2225.345 215.510 ;
      LAYER li1 ;
        RECT 2225.515 214.490 2225.845 215.290 ;
      LAYER li1 ;
        RECT 2226.015 214.660 2226.185 215.510 ;
      LAYER li1 ;
        RECT 2226.355 214.490 2226.685 215.290 ;
      LAYER li1 ;
        RECT 2226.855 214.660 2227.025 215.510 ;
      LAYER li1 ;
        RECT 2227.195 214.490 2227.525 215.290 ;
      LAYER li1 ;
        RECT 2227.695 214.660 2227.865 215.510 ;
      LAYER li1 ;
        RECT 2228.115 214.490 2228.285 215.290 ;
        RECT 2228.455 214.660 2228.785 215.510 ;
        RECT 2228.955 214.490 2229.125 215.290 ;
        RECT 2229.295 214.660 2229.625 215.510 ;
        RECT 2229.805 214.490 2230.095 215.655 ;
        RECT 2230.655 214.490 2230.985 215.640 ;
      LAYER li1 ;
        RECT 2231.155 215.510 2233.845 215.680 ;
      LAYER li1 ;
        RECT 2234.105 215.510 2235.605 215.680 ;
      LAYER li1 ;
        RECT 2231.155 214.660 2231.325 215.510 ;
      LAYER li1 ;
        RECT 2231.495 214.490 2231.825 215.290 ;
      LAYER li1 ;
        RECT 2231.995 214.660 2232.165 215.510 ;
      LAYER li1 ;
        RECT 2232.335 214.490 2232.665 215.290 ;
      LAYER li1 ;
        RECT 2232.835 214.660 2233.005 215.510 ;
      LAYER li1 ;
        RECT 2233.175 214.490 2233.505 215.290 ;
      LAYER li1 ;
        RECT 2233.675 214.660 2233.845 215.510 ;
      LAYER li1 ;
        RECT 2234.095 214.490 2234.265 215.290 ;
        RECT 2234.435 214.660 2234.765 215.510 ;
        RECT 2234.935 214.490 2235.105 215.290 ;
        RECT 2235.275 214.660 2235.605 215.510 ;
        RECT 2235.785 214.490 2236.075 215.655 ;
        RECT 2236.635 214.490 2236.965 215.640 ;
      LAYER li1 ;
        RECT 2237.135 215.510 2239.825 215.680 ;
      LAYER li1 ;
        RECT 2240.085 215.510 2241.585 215.680 ;
      LAYER li1 ;
        RECT 2237.135 214.660 2237.305 215.510 ;
      LAYER li1 ;
        RECT 2237.475 214.490 2237.805 215.290 ;
      LAYER li1 ;
        RECT 2237.975 214.660 2238.145 215.510 ;
      LAYER li1 ;
        RECT 2238.315 214.490 2238.645 215.290 ;
      LAYER li1 ;
        RECT 2238.815 214.660 2238.985 215.510 ;
      LAYER li1 ;
        RECT 2239.155 214.490 2239.485 215.290 ;
      LAYER li1 ;
        RECT 2239.655 214.660 2239.825 215.510 ;
      LAYER li1 ;
        RECT 2240.075 214.490 2240.245 215.290 ;
        RECT 2240.415 214.660 2240.745 215.510 ;
        RECT 2240.915 214.490 2241.085 215.290 ;
        RECT 2241.255 214.660 2241.585 215.510 ;
        RECT 2241.765 214.490 2242.055 215.655 ;
        RECT 2242.615 214.490 2242.945 215.640 ;
      LAYER li1 ;
        RECT 2243.115 215.510 2245.805 215.680 ;
      LAYER li1 ;
        RECT 2246.065 215.510 2247.565 215.680 ;
      LAYER li1 ;
        RECT 2243.115 214.660 2243.285 215.510 ;
      LAYER li1 ;
        RECT 2243.455 214.490 2243.785 215.290 ;
      LAYER li1 ;
        RECT 2243.955 214.660 2244.125 215.510 ;
      LAYER li1 ;
        RECT 2244.295 214.490 2244.625 215.290 ;
      LAYER li1 ;
        RECT 2244.795 214.660 2244.965 215.510 ;
      LAYER li1 ;
        RECT 2245.135 214.490 2245.465 215.290 ;
      LAYER li1 ;
        RECT 2245.635 214.660 2245.805 215.510 ;
      LAYER li1 ;
        RECT 2246.055 214.490 2246.225 215.290 ;
        RECT 2246.395 214.660 2246.725 215.510 ;
        RECT 2246.895 214.490 2247.065 215.290 ;
        RECT 2247.235 214.660 2247.565 215.510 ;
        RECT 2247.745 214.490 2248.035 215.655 ;
        RECT 2248.595 214.490 2248.925 215.640 ;
      LAYER li1 ;
        RECT 2249.095 215.510 2251.785 215.680 ;
      LAYER li1 ;
        RECT 2252.045 215.510 2253.545 215.680 ;
      LAYER li1 ;
        RECT 2249.095 214.660 2249.265 215.510 ;
      LAYER li1 ;
        RECT 2249.435 214.490 2249.765 215.290 ;
      LAYER li1 ;
        RECT 2249.935 214.660 2250.105 215.510 ;
      LAYER li1 ;
        RECT 2250.275 214.490 2250.605 215.290 ;
      LAYER li1 ;
        RECT 2250.775 214.660 2250.945 215.510 ;
      LAYER li1 ;
        RECT 2251.115 214.490 2251.445 215.290 ;
      LAYER li1 ;
        RECT 2251.615 214.660 2251.785 215.510 ;
      LAYER li1 ;
        RECT 2252.035 214.490 2252.205 215.290 ;
        RECT 2252.375 214.660 2252.705 215.510 ;
        RECT 2252.875 214.490 2253.045 215.290 ;
        RECT 2253.215 214.660 2253.545 215.510 ;
        RECT 2253.725 214.490 2254.015 215.655 ;
        RECT 2254.575 214.490 2254.905 215.640 ;
      LAYER li1 ;
        RECT 2255.075 215.510 2257.765 215.680 ;
      LAYER li1 ;
        RECT 2258.025 215.510 2259.525 215.680 ;
      LAYER li1 ;
        RECT 2255.075 214.660 2255.245 215.510 ;
      LAYER li1 ;
        RECT 2255.415 214.490 2255.745 215.290 ;
      LAYER li1 ;
        RECT 2255.915 214.660 2256.085 215.510 ;
      LAYER li1 ;
        RECT 2256.255 214.490 2256.585 215.290 ;
      LAYER li1 ;
        RECT 2256.755 214.660 2256.925 215.510 ;
      LAYER li1 ;
        RECT 2257.095 214.490 2257.425 215.290 ;
      LAYER li1 ;
        RECT 2257.595 214.660 2257.765 215.510 ;
      LAYER li1 ;
        RECT 2258.015 214.490 2258.185 215.290 ;
        RECT 2258.355 214.660 2258.685 215.510 ;
        RECT 2258.855 214.490 2259.025 215.290 ;
        RECT 2259.195 214.660 2259.525 215.510 ;
        RECT 2259.705 214.490 2259.995 215.655 ;
        RECT 2260.555 214.490 2260.885 215.640 ;
      LAYER li1 ;
        RECT 2261.055 215.510 2263.745 215.680 ;
      LAYER li1 ;
        RECT 2264.005 215.510 2265.505 215.680 ;
      LAYER li1 ;
        RECT 2261.055 214.660 2261.225 215.510 ;
      LAYER li1 ;
        RECT 2261.395 214.490 2261.725 215.290 ;
      LAYER li1 ;
        RECT 2261.895 214.660 2262.065 215.510 ;
      LAYER li1 ;
        RECT 2262.235 214.490 2262.565 215.290 ;
      LAYER li1 ;
        RECT 2262.735 214.660 2262.905 215.510 ;
      LAYER li1 ;
        RECT 2263.075 214.490 2263.405 215.290 ;
      LAYER li1 ;
        RECT 2263.575 214.660 2263.745 215.510 ;
      LAYER li1 ;
        RECT 2263.995 214.490 2264.165 215.290 ;
        RECT 2264.335 214.660 2264.665 215.510 ;
        RECT 2264.835 214.490 2265.005 215.290 ;
        RECT 2265.175 214.660 2265.505 215.510 ;
        RECT 2265.685 214.490 2265.975 215.655 ;
        RECT 2266.535 214.490 2266.865 215.640 ;
      LAYER li1 ;
        RECT 2267.035 215.510 2269.725 215.680 ;
      LAYER li1 ;
        RECT 2269.985 215.510 2271.485 215.680 ;
      LAYER li1 ;
        RECT 2267.035 214.660 2267.205 215.510 ;
      LAYER li1 ;
        RECT 2267.375 214.490 2267.705 215.290 ;
      LAYER li1 ;
        RECT 2267.875 214.660 2268.045 215.510 ;
      LAYER li1 ;
        RECT 2268.215 214.490 2268.545 215.290 ;
      LAYER li1 ;
        RECT 2268.715 214.660 2268.885 215.510 ;
      LAYER li1 ;
        RECT 2269.055 214.490 2269.385 215.290 ;
      LAYER li1 ;
        RECT 2269.555 214.660 2269.725 215.510 ;
      LAYER li1 ;
        RECT 2269.975 214.490 2270.145 215.290 ;
        RECT 2270.315 214.660 2270.645 215.510 ;
        RECT 2270.815 214.490 2270.985 215.290 ;
        RECT 2271.155 214.660 2271.485 215.510 ;
        RECT 2271.665 214.490 2271.955 215.655 ;
        RECT 669.000 214.320 669.145 214.490 ;
        RECT 669.315 214.320 669.605 214.490 ;
        RECT 669.775 214.320 670.065 214.490 ;
        RECT 670.235 214.320 670.525 214.490 ;
        RECT 670.695 214.320 670.985 214.490 ;
        RECT 671.155 214.320 671.445 214.490 ;
        RECT 671.615 214.320 671.905 214.490 ;
        RECT 672.075 214.320 672.365 214.490 ;
        RECT 672.535 214.320 672.825 214.490 ;
        RECT 672.995 214.320 673.285 214.490 ;
        RECT 673.455 214.320 673.745 214.490 ;
        RECT 673.915 214.320 674.205 214.490 ;
        RECT 674.375 214.320 674.665 214.490 ;
        RECT 674.835 214.320 675.125 214.490 ;
        RECT 675.295 214.320 675.585 214.490 ;
        RECT 675.755 214.320 676.045 214.490 ;
        RECT 676.215 214.320 676.505 214.490 ;
        RECT 676.675 214.320 676.965 214.490 ;
        RECT 677.135 214.320 677.425 214.490 ;
        RECT 677.595 214.320 677.885 214.490 ;
        RECT 678.055 214.320 678.345 214.490 ;
        RECT 678.515 214.320 678.805 214.490 ;
        RECT 678.975 214.320 679.265 214.490 ;
        RECT 679.435 214.320 679.725 214.490 ;
        RECT 679.895 214.320 680.185 214.490 ;
        RECT 680.355 214.320 680.645 214.490 ;
        RECT 680.815 214.320 681.105 214.490 ;
        RECT 681.275 214.320 681.565 214.490 ;
        RECT 681.735 214.320 682.025 214.490 ;
        RECT 682.195 214.320 682.485 214.490 ;
        RECT 682.655 214.320 682.945 214.490 ;
        RECT 683.115 214.320 683.405 214.490 ;
        RECT 683.575 214.320 683.865 214.490 ;
        RECT 684.035 214.320 684.325 214.490 ;
        RECT 684.495 214.320 684.785 214.490 ;
        RECT 684.955 214.320 685.245 214.490 ;
        RECT 685.415 214.320 685.705 214.490 ;
        RECT 685.875 214.320 686.165 214.490 ;
        RECT 686.335 214.320 686.625 214.490 ;
        RECT 686.795 214.320 687.085 214.490 ;
        RECT 687.255 214.320 687.545 214.490 ;
        RECT 687.715 214.320 688.005 214.490 ;
        RECT 688.175 214.320 688.465 214.490 ;
        RECT 688.635 214.320 688.925 214.490 ;
        RECT 689.095 214.320 689.385 214.490 ;
        RECT 689.555 214.320 689.845 214.490 ;
        RECT 690.015 214.320 690.305 214.490 ;
        RECT 690.475 214.320 690.765 214.490 ;
        RECT 690.935 214.320 691.225 214.490 ;
        RECT 691.395 214.320 691.685 214.490 ;
        RECT 691.855 214.320 692.145 214.490 ;
        RECT 692.315 214.320 692.605 214.490 ;
        RECT 692.775 214.320 693.065 214.490 ;
        RECT 693.235 214.320 693.525 214.490 ;
        RECT 693.695 214.320 693.985 214.490 ;
        RECT 694.155 214.320 694.445 214.490 ;
        RECT 694.615 214.320 694.905 214.490 ;
        RECT 695.075 214.320 695.365 214.490 ;
        RECT 695.535 214.320 695.825 214.490 ;
        RECT 695.995 214.320 696.285 214.490 ;
        RECT 696.455 214.320 696.745 214.490 ;
        RECT 696.915 214.320 697.205 214.490 ;
        RECT 697.375 214.320 697.665 214.490 ;
        RECT 697.835 214.320 698.125 214.490 ;
        RECT 698.295 214.320 698.585 214.490 ;
        RECT 698.755 214.320 699.045 214.490 ;
        RECT 699.215 214.320 699.505 214.490 ;
        RECT 699.675 214.320 699.965 214.490 ;
        RECT 700.135 214.320 700.425 214.490 ;
        RECT 700.595 214.320 700.885 214.490 ;
        RECT 701.055 214.320 701.345 214.490 ;
        RECT 701.515 214.320 701.805 214.490 ;
        RECT 701.975 214.320 702.265 214.490 ;
        RECT 702.435 214.320 702.725 214.490 ;
        RECT 702.895 214.320 703.185 214.490 ;
        RECT 703.355 214.320 703.645 214.490 ;
        RECT 703.815 214.320 704.105 214.490 ;
        RECT 704.275 214.320 704.565 214.490 ;
        RECT 704.735 214.320 705.025 214.490 ;
        RECT 705.195 214.320 705.485 214.490 ;
        RECT 705.655 214.320 705.945 214.490 ;
        RECT 706.115 214.320 706.405 214.490 ;
        RECT 706.575 214.320 706.865 214.490 ;
        RECT 707.035 214.320 707.325 214.490 ;
        RECT 707.495 214.320 707.785 214.490 ;
        RECT 707.955 214.320 708.245 214.490 ;
        RECT 708.415 214.320 708.705 214.490 ;
        RECT 708.875 214.320 709.165 214.490 ;
        RECT 709.335 214.320 709.625 214.490 ;
        RECT 709.795 214.320 710.085 214.490 ;
        RECT 710.255 214.320 710.545 214.490 ;
        RECT 710.715 214.320 711.005 214.490 ;
        RECT 711.175 214.320 711.465 214.490 ;
        RECT 711.635 214.320 711.925 214.490 ;
        RECT 712.095 214.320 712.385 214.490 ;
        RECT 712.555 214.320 712.845 214.490 ;
        RECT 713.015 214.320 713.305 214.490 ;
        RECT 713.475 214.320 713.765 214.490 ;
        RECT 713.935 214.320 714.225 214.490 ;
        RECT 714.395 214.320 714.685 214.490 ;
        RECT 714.855 214.320 715.145 214.490 ;
        RECT 715.315 214.320 715.605 214.490 ;
        RECT 715.775 214.320 716.065 214.490 ;
        RECT 716.235 214.320 716.525 214.490 ;
        RECT 716.695 214.320 716.985 214.490 ;
        RECT 717.155 214.320 717.445 214.490 ;
        RECT 717.615 214.320 717.905 214.490 ;
        RECT 718.075 214.320 718.365 214.490 ;
        RECT 718.535 214.320 718.825 214.490 ;
        RECT 718.995 214.320 719.285 214.490 ;
        RECT 719.455 214.320 719.745 214.490 ;
        RECT 719.915 214.320 720.205 214.490 ;
        RECT 720.375 214.320 720.665 214.490 ;
        RECT 720.835 214.320 721.125 214.490 ;
        RECT 721.295 214.320 721.585 214.490 ;
        RECT 721.755 214.320 722.045 214.490 ;
        RECT 722.215 214.320 722.505 214.490 ;
        RECT 722.675 214.320 722.965 214.490 ;
        RECT 723.135 214.320 723.425 214.490 ;
        RECT 723.595 214.320 723.885 214.490 ;
        RECT 724.055 214.320 724.345 214.490 ;
        RECT 724.515 214.320 724.805 214.490 ;
        RECT 724.975 214.320 725.265 214.490 ;
        RECT 725.435 214.320 725.725 214.490 ;
        RECT 725.895 214.320 726.185 214.490 ;
        RECT 726.355 214.320 726.645 214.490 ;
        RECT 726.815 214.320 727.105 214.490 ;
        RECT 727.275 214.320 727.565 214.490 ;
        RECT 727.735 214.320 728.025 214.490 ;
        RECT 728.195 214.320 728.485 214.490 ;
        RECT 728.655 214.320 728.945 214.490 ;
        RECT 729.115 214.320 729.405 214.490 ;
        RECT 729.575 214.320 729.865 214.490 ;
        RECT 730.035 214.320 730.325 214.490 ;
        RECT 730.495 214.320 730.785 214.490 ;
        RECT 730.955 214.320 731.245 214.490 ;
        RECT 731.415 214.320 731.705 214.490 ;
        RECT 731.875 214.320 732.165 214.490 ;
        RECT 732.335 214.320 732.625 214.490 ;
        RECT 732.795 214.320 733.085 214.490 ;
        RECT 733.255 214.320 733.545 214.490 ;
        RECT 733.715 214.320 734.005 214.490 ;
        RECT 734.175 214.320 734.465 214.490 ;
        RECT 734.635 214.320 734.925 214.490 ;
        RECT 735.095 214.320 735.385 214.490 ;
        RECT 735.555 214.320 735.845 214.490 ;
        RECT 736.015 214.320 736.305 214.490 ;
        RECT 736.475 214.320 736.765 214.490 ;
        RECT 736.935 214.320 737.225 214.490 ;
        RECT 737.395 214.320 737.685 214.490 ;
        RECT 737.855 214.320 738.145 214.490 ;
        RECT 738.315 214.320 738.605 214.490 ;
        RECT 738.775 214.320 739.065 214.490 ;
        RECT 739.235 214.320 739.525 214.490 ;
        RECT 739.695 214.320 739.985 214.490 ;
        RECT 740.155 214.320 740.445 214.490 ;
        RECT 740.615 214.320 740.905 214.490 ;
        RECT 741.075 214.320 741.365 214.490 ;
        RECT 741.535 214.320 741.825 214.490 ;
        RECT 741.995 214.320 742.285 214.490 ;
        RECT 742.455 214.320 742.745 214.490 ;
        RECT 742.915 214.320 743.205 214.490 ;
        RECT 743.375 214.320 743.665 214.490 ;
        RECT 743.835 214.320 744.125 214.490 ;
        RECT 744.295 214.320 744.585 214.490 ;
        RECT 744.755 214.320 745.045 214.490 ;
        RECT 745.215 214.320 745.505 214.490 ;
        RECT 745.675 214.320 745.965 214.490 ;
        RECT 746.135 214.320 746.425 214.490 ;
        RECT 746.595 214.320 746.885 214.490 ;
        RECT 747.055 214.320 747.345 214.490 ;
        RECT 747.515 214.320 747.805 214.490 ;
        RECT 747.975 214.320 748.265 214.490 ;
        RECT 748.435 214.320 748.725 214.490 ;
        RECT 748.895 214.320 749.185 214.490 ;
        RECT 749.355 214.320 749.645 214.490 ;
        RECT 749.815 214.320 750.105 214.490 ;
        RECT 750.275 214.320 750.565 214.490 ;
        RECT 750.735 214.320 751.025 214.490 ;
        RECT 751.195 214.320 751.485 214.490 ;
        RECT 751.655 214.320 751.945 214.490 ;
        RECT 752.115 214.320 752.405 214.490 ;
        RECT 752.575 214.320 752.865 214.490 ;
        RECT 753.035 214.320 753.325 214.490 ;
        RECT 753.495 214.320 753.785 214.490 ;
        RECT 753.955 214.320 754.245 214.490 ;
        RECT 754.415 214.320 754.705 214.490 ;
        RECT 754.875 214.320 755.165 214.490 ;
        RECT 755.335 214.320 755.625 214.490 ;
        RECT 755.795 214.320 756.085 214.490 ;
        RECT 756.255 214.320 756.545 214.490 ;
        RECT 756.715 214.320 757.005 214.490 ;
        RECT 757.175 214.320 757.465 214.490 ;
        RECT 757.635 214.320 757.925 214.490 ;
        RECT 758.095 214.320 758.385 214.490 ;
        RECT 758.555 214.320 758.845 214.490 ;
        RECT 759.015 214.320 759.305 214.490 ;
        RECT 759.475 214.320 759.765 214.490 ;
        RECT 759.935 214.320 760.225 214.490 ;
        RECT 760.395 214.320 760.685 214.490 ;
        RECT 760.855 214.320 761.145 214.490 ;
        RECT 761.315 214.320 761.605 214.490 ;
        RECT 761.775 214.320 762.065 214.490 ;
        RECT 762.235 214.320 762.525 214.490 ;
        RECT 762.695 214.320 762.985 214.490 ;
        RECT 763.155 214.320 763.445 214.490 ;
        RECT 763.615 214.320 763.905 214.490 ;
        RECT 764.075 214.320 764.365 214.490 ;
        RECT 764.535 214.320 764.825 214.490 ;
        RECT 764.995 214.320 765.285 214.490 ;
        RECT 765.455 214.320 765.745 214.490 ;
        RECT 765.915 214.320 766.205 214.490 ;
        RECT 766.375 214.320 766.665 214.490 ;
        RECT 766.835 214.320 767.125 214.490 ;
        RECT 767.295 214.320 767.585 214.490 ;
        RECT 767.755 214.320 768.045 214.490 ;
        RECT 768.215 214.320 768.505 214.490 ;
        RECT 768.675 214.320 768.965 214.490 ;
        RECT 769.135 214.320 769.425 214.490 ;
        RECT 769.595 214.320 769.885 214.490 ;
        RECT 770.055 214.320 770.345 214.490 ;
        RECT 770.515 214.320 770.805 214.490 ;
        RECT 770.975 214.320 771.265 214.490 ;
        RECT 771.435 214.320 771.725 214.490 ;
        RECT 771.895 214.320 772.185 214.490 ;
        RECT 772.355 214.320 772.645 214.490 ;
        RECT 772.815 214.320 773.105 214.490 ;
        RECT 773.275 214.320 773.565 214.490 ;
        RECT 773.735 214.320 774.025 214.490 ;
        RECT 774.195 214.320 774.485 214.490 ;
        RECT 774.655 214.320 774.945 214.490 ;
        RECT 775.115 214.320 775.405 214.490 ;
        RECT 775.575 214.320 775.865 214.490 ;
        RECT 776.035 214.320 776.325 214.490 ;
        RECT 776.495 214.320 776.785 214.490 ;
        RECT 776.955 214.320 777.245 214.490 ;
        RECT 777.415 214.320 777.705 214.490 ;
        RECT 777.875 214.320 778.165 214.490 ;
        RECT 778.335 214.320 778.625 214.490 ;
        RECT 778.795 214.320 779.085 214.490 ;
        RECT 779.255 214.320 779.545 214.490 ;
        RECT 779.715 214.320 780.005 214.490 ;
        RECT 780.175 214.320 780.465 214.490 ;
        RECT 780.635 214.320 780.925 214.490 ;
        RECT 781.095 214.320 781.385 214.490 ;
        RECT 781.555 214.320 781.845 214.490 ;
        RECT 782.015 214.320 782.305 214.490 ;
        RECT 782.475 214.320 782.765 214.490 ;
        RECT 782.935 214.320 783.225 214.490 ;
        RECT 783.395 214.320 783.685 214.490 ;
        RECT 783.855 214.320 784.145 214.490 ;
        RECT 784.315 214.320 784.605 214.490 ;
        RECT 784.775 214.320 785.065 214.490 ;
        RECT 785.235 214.320 785.525 214.490 ;
        RECT 785.695 214.320 785.985 214.490 ;
        RECT 786.155 214.320 786.445 214.490 ;
        RECT 786.615 214.320 786.905 214.490 ;
        RECT 787.075 214.320 787.365 214.490 ;
        RECT 787.535 214.320 787.825 214.490 ;
        RECT 787.995 214.320 788.285 214.490 ;
        RECT 788.455 214.320 788.745 214.490 ;
        RECT 788.915 214.320 789.205 214.490 ;
        RECT 789.375 214.320 789.665 214.490 ;
        RECT 789.835 214.320 790.125 214.490 ;
        RECT 790.295 214.320 790.585 214.490 ;
        RECT 790.755 214.320 791.045 214.490 ;
        RECT 791.215 214.320 791.505 214.490 ;
        RECT 791.675 214.320 791.965 214.490 ;
        RECT 792.135 214.320 792.425 214.490 ;
        RECT 792.595 214.320 792.885 214.490 ;
        RECT 793.055 214.320 793.345 214.490 ;
        RECT 793.515 214.320 793.805 214.490 ;
        RECT 793.975 214.320 794.265 214.490 ;
        RECT 794.435 214.320 794.725 214.490 ;
        RECT 794.895 214.320 795.040 214.490 ;
        RECT 2146.000 214.320 2146.145 214.490 ;
        RECT 2146.315 214.320 2146.605 214.490 ;
        RECT 2146.775 214.320 2147.065 214.490 ;
        RECT 2147.235 214.320 2147.525 214.490 ;
        RECT 2147.695 214.320 2147.985 214.490 ;
        RECT 2148.155 214.320 2148.445 214.490 ;
        RECT 2148.615 214.320 2148.905 214.490 ;
        RECT 2149.075 214.320 2149.365 214.490 ;
        RECT 2149.535 214.320 2149.825 214.490 ;
        RECT 2149.995 214.320 2150.285 214.490 ;
        RECT 2150.455 214.320 2150.745 214.490 ;
        RECT 2150.915 214.320 2151.205 214.490 ;
        RECT 2151.375 214.320 2151.665 214.490 ;
        RECT 2151.835 214.320 2152.125 214.490 ;
        RECT 2152.295 214.320 2152.585 214.490 ;
        RECT 2152.755 214.320 2153.045 214.490 ;
        RECT 2153.215 214.320 2153.505 214.490 ;
        RECT 2153.675 214.320 2153.965 214.490 ;
        RECT 2154.135 214.320 2154.425 214.490 ;
        RECT 2154.595 214.320 2154.885 214.490 ;
        RECT 2155.055 214.320 2155.345 214.490 ;
        RECT 2155.515 214.320 2155.805 214.490 ;
        RECT 2155.975 214.320 2156.265 214.490 ;
        RECT 2156.435 214.320 2156.725 214.490 ;
        RECT 2156.895 214.320 2157.185 214.490 ;
        RECT 2157.355 214.320 2157.645 214.490 ;
        RECT 2157.815 214.320 2158.105 214.490 ;
        RECT 2158.275 214.320 2158.565 214.490 ;
        RECT 2158.735 214.320 2159.025 214.490 ;
        RECT 2159.195 214.320 2159.485 214.490 ;
        RECT 2159.655 214.320 2159.945 214.490 ;
        RECT 2160.115 214.320 2160.405 214.490 ;
        RECT 2160.575 214.320 2160.865 214.490 ;
        RECT 2161.035 214.320 2161.325 214.490 ;
        RECT 2161.495 214.320 2161.785 214.490 ;
        RECT 2161.955 214.320 2162.245 214.490 ;
        RECT 2162.415 214.320 2162.705 214.490 ;
        RECT 2162.875 214.320 2163.165 214.490 ;
        RECT 2163.335 214.320 2163.625 214.490 ;
        RECT 2163.795 214.320 2164.085 214.490 ;
        RECT 2164.255 214.320 2164.545 214.490 ;
        RECT 2164.715 214.320 2165.005 214.490 ;
        RECT 2165.175 214.320 2165.465 214.490 ;
        RECT 2165.635 214.320 2165.925 214.490 ;
        RECT 2166.095 214.320 2166.385 214.490 ;
        RECT 2166.555 214.320 2166.845 214.490 ;
        RECT 2167.015 214.320 2167.305 214.490 ;
        RECT 2167.475 214.320 2167.765 214.490 ;
        RECT 2167.935 214.320 2168.225 214.490 ;
        RECT 2168.395 214.320 2168.685 214.490 ;
        RECT 2168.855 214.320 2169.145 214.490 ;
        RECT 2169.315 214.320 2169.605 214.490 ;
        RECT 2169.775 214.320 2170.065 214.490 ;
        RECT 2170.235 214.320 2170.525 214.490 ;
        RECT 2170.695 214.320 2170.985 214.490 ;
        RECT 2171.155 214.320 2171.445 214.490 ;
        RECT 2171.615 214.320 2171.905 214.490 ;
        RECT 2172.075 214.320 2172.365 214.490 ;
        RECT 2172.535 214.320 2172.825 214.490 ;
        RECT 2172.995 214.320 2173.285 214.490 ;
        RECT 2173.455 214.320 2173.745 214.490 ;
        RECT 2173.915 214.320 2174.205 214.490 ;
        RECT 2174.375 214.320 2174.665 214.490 ;
        RECT 2174.835 214.320 2175.125 214.490 ;
        RECT 2175.295 214.320 2175.585 214.490 ;
        RECT 2175.755 214.320 2176.045 214.490 ;
        RECT 2176.215 214.320 2176.505 214.490 ;
        RECT 2176.675 214.320 2176.965 214.490 ;
        RECT 2177.135 214.320 2177.425 214.490 ;
        RECT 2177.595 214.320 2177.885 214.490 ;
        RECT 2178.055 214.320 2178.345 214.490 ;
        RECT 2178.515 214.320 2178.805 214.490 ;
        RECT 2178.975 214.320 2179.265 214.490 ;
        RECT 2179.435 214.320 2179.725 214.490 ;
        RECT 2179.895 214.320 2180.185 214.490 ;
        RECT 2180.355 214.320 2180.645 214.490 ;
        RECT 2180.815 214.320 2181.105 214.490 ;
        RECT 2181.275 214.320 2181.565 214.490 ;
        RECT 2181.735 214.320 2182.025 214.490 ;
        RECT 2182.195 214.320 2182.485 214.490 ;
        RECT 2182.655 214.320 2182.945 214.490 ;
        RECT 2183.115 214.320 2183.405 214.490 ;
        RECT 2183.575 214.320 2183.865 214.490 ;
        RECT 2184.035 214.320 2184.325 214.490 ;
        RECT 2184.495 214.320 2184.785 214.490 ;
        RECT 2184.955 214.320 2185.245 214.490 ;
        RECT 2185.415 214.320 2185.705 214.490 ;
        RECT 2185.875 214.320 2186.165 214.490 ;
        RECT 2186.335 214.320 2186.625 214.490 ;
        RECT 2186.795 214.320 2187.085 214.490 ;
        RECT 2187.255 214.320 2187.545 214.490 ;
        RECT 2187.715 214.320 2188.005 214.490 ;
        RECT 2188.175 214.320 2188.465 214.490 ;
        RECT 2188.635 214.320 2188.925 214.490 ;
        RECT 2189.095 214.320 2189.385 214.490 ;
        RECT 2189.555 214.320 2189.845 214.490 ;
        RECT 2190.015 214.320 2190.305 214.490 ;
        RECT 2190.475 214.320 2190.765 214.490 ;
        RECT 2190.935 214.320 2191.225 214.490 ;
        RECT 2191.395 214.320 2191.685 214.490 ;
        RECT 2191.855 214.320 2192.145 214.490 ;
        RECT 2192.315 214.320 2192.605 214.490 ;
        RECT 2192.775 214.320 2193.065 214.490 ;
        RECT 2193.235 214.320 2193.525 214.490 ;
        RECT 2193.695 214.320 2193.985 214.490 ;
        RECT 2194.155 214.320 2194.445 214.490 ;
        RECT 2194.615 214.320 2194.905 214.490 ;
        RECT 2195.075 214.320 2195.365 214.490 ;
        RECT 2195.535 214.320 2195.825 214.490 ;
        RECT 2195.995 214.320 2196.285 214.490 ;
        RECT 2196.455 214.320 2196.745 214.490 ;
        RECT 2196.915 214.320 2197.205 214.490 ;
        RECT 2197.375 214.320 2197.665 214.490 ;
        RECT 2197.835 214.320 2198.125 214.490 ;
        RECT 2198.295 214.320 2198.585 214.490 ;
        RECT 2198.755 214.320 2199.045 214.490 ;
        RECT 2199.215 214.320 2199.505 214.490 ;
        RECT 2199.675 214.320 2199.965 214.490 ;
        RECT 2200.135 214.320 2200.425 214.490 ;
        RECT 2200.595 214.320 2200.885 214.490 ;
        RECT 2201.055 214.320 2201.345 214.490 ;
        RECT 2201.515 214.320 2201.805 214.490 ;
        RECT 2201.975 214.320 2202.265 214.490 ;
        RECT 2202.435 214.320 2202.725 214.490 ;
        RECT 2202.895 214.320 2203.185 214.490 ;
        RECT 2203.355 214.320 2203.645 214.490 ;
        RECT 2203.815 214.320 2204.105 214.490 ;
        RECT 2204.275 214.320 2204.565 214.490 ;
        RECT 2204.735 214.320 2205.025 214.490 ;
        RECT 2205.195 214.320 2205.485 214.490 ;
        RECT 2205.655 214.320 2205.945 214.490 ;
        RECT 2206.115 214.320 2206.405 214.490 ;
        RECT 2206.575 214.320 2206.865 214.490 ;
        RECT 2207.035 214.320 2207.325 214.490 ;
        RECT 2207.495 214.320 2207.785 214.490 ;
        RECT 2207.955 214.320 2208.245 214.490 ;
        RECT 2208.415 214.320 2208.705 214.490 ;
        RECT 2208.875 214.320 2209.165 214.490 ;
        RECT 2209.335 214.320 2209.625 214.490 ;
        RECT 2209.795 214.320 2210.085 214.490 ;
        RECT 2210.255 214.320 2210.545 214.490 ;
        RECT 2210.715 214.320 2211.005 214.490 ;
        RECT 2211.175 214.320 2211.465 214.490 ;
        RECT 2211.635 214.320 2211.925 214.490 ;
        RECT 2212.095 214.320 2212.385 214.490 ;
        RECT 2212.555 214.320 2212.845 214.490 ;
        RECT 2213.015 214.320 2213.305 214.490 ;
        RECT 2213.475 214.320 2213.765 214.490 ;
        RECT 2213.935 214.320 2214.225 214.490 ;
        RECT 2214.395 214.320 2214.685 214.490 ;
        RECT 2214.855 214.320 2215.145 214.490 ;
        RECT 2215.315 214.320 2215.605 214.490 ;
        RECT 2215.775 214.320 2216.065 214.490 ;
        RECT 2216.235 214.320 2216.525 214.490 ;
        RECT 2216.695 214.320 2216.985 214.490 ;
        RECT 2217.155 214.320 2217.445 214.490 ;
        RECT 2217.615 214.320 2217.905 214.490 ;
        RECT 2218.075 214.320 2218.365 214.490 ;
        RECT 2218.535 214.320 2218.825 214.490 ;
        RECT 2218.995 214.320 2219.285 214.490 ;
        RECT 2219.455 214.320 2219.745 214.490 ;
        RECT 2219.915 214.320 2220.205 214.490 ;
        RECT 2220.375 214.320 2220.665 214.490 ;
        RECT 2220.835 214.320 2221.125 214.490 ;
        RECT 2221.295 214.320 2221.585 214.490 ;
        RECT 2221.755 214.320 2222.045 214.490 ;
        RECT 2222.215 214.320 2222.505 214.490 ;
        RECT 2222.675 214.320 2222.965 214.490 ;
        RECT 2223.135 214.320 2223.425 214.490 ;
        RECT 2223.595 214.320 2223.885 214.490 ;
        RECT 2224.055 214.320 2224.345 214.490 ;
        RECT 2224.515 214.320 2224.805 214.490 ;
        RECT 2224.975 214.320 2225.265 214.490 ;
        RECT 2225.435 214.320 2225.725 214.490 ;
        RECT 2225.895 214.320 2226.185 214.490 ;
        RECT 2226.355 214.320 2226.645 214.490 ;
        RECT 2226.815 214.320 2227.105 214.490 ;
        RECT 2227.275 214.320 2227.565 214.490 ;
        RECT 2227.735 214.320 2228.025 214.490 ;
        RECT 2228.195 214.320 2228.485 214.490 ;
        RECT 2228.655 214.320 2228.945 214.490 ;
        RECT 2229.115 214.320 2229.405 214.490 ;
        RECT 2229.575 214.320 2229.865 214.490 ;
        RECT 2230.035 214.320 2230.325 214.490 ;
        RECT 2230.495 214.320 2230.785 214.490 ;
        RECT 2230.955 214.320 2231.245 214.490 ;
        RECT 2231.415 214.320 2231.705 214.490 ;
        RECT 2231.875 214.320 2232.165 214.490 ;
        RECT 2232.335 214.320 2232.625 214.490 ;
        RECT 2232.795 214.320 2233.085 214.490 ;
        RECT 2233.255 214.320 2233.545 214.490 ;
        RECT 2233.715 214.320 2234.005 214.490 ;
        RECT 2234.175 214.320 2234.465 214.490 ;
        RECT 2234.635 214.320 2234.925 214.490 ;
        RECT 2235.095 214.320 2235.385 214.490 ;
        RECT 2235.555 214.320 2235.845 214.490 ;
        RECT 2236.015 214.320 2236.305 214.490 ;
        RECT 2236.475 214.320 2236.765 214.490 ;
        RECT 2236.935 214.320 2237.225 214.490 ;
        RECT 2237.395 214.320 2237.685 214.490 ;
        RECT 2237.855 214.320 2238.145 214.490 ;
        RECT 2238.315 214.320 2238.605 214.490 ;
        RECT 2238.775 214.320 2239.065 214.490 ;
        RECT 2239.235 214.320 2239.525 214.490 ;
        RECT 2239.695 214.320 2239.985 214.490 ;
        RECT 2240.155 214.320 2240.445 214.490 ;
        RECT 2240.615 214.320 2240.905 214.490 ;
        RECT 2241.075 214.320 2241.365 214.490 ;
        RECT 2241.535 214.320 2241.825 214.490 ;
        RECT 2241.995 214.320 2242.285 214.490 ;
        RECT 2242.455 214.320 2242.745 214.490 ;
        RECT 2242.915 214.320 2243.205 214.490 ;
        RECT 2243.375 214.320 2243.665 214.490 ;
        RECT 2243.835 214.320 2244.125 214.490 ;
        RECT 2244.295 214.320 2244.585 214.490 ;
        RECT 2244.755 214.320 2245.045 214.490 ;
        RECT 2245.215 214.320 2245.505 214.490 ;
        RECT 2245.675 214.320 2245.965 214.490 ;
        RECT 2246.135 214.320 2246.425 214.490 ;
        RECT 2246.595 214.320 2246.885 214.490 ;
        RECT 2247.055 214.320 2247.345 214.490 ;
        RECT 2247.515 214.320 2247.805 214.490 ;
        RECT 2247.975 214.320 2248.265 214.490 ;
        RECT 2248.435 214.320 2248.725 214.490 ;
        RECT 2248.895 214.320 2249.185 214.490 ;
        RECT 2249.355 214.320 2249.645 214.490 ;
        RECT 2249.815 214.320 2250.105 214.490 ;
        RECT 2250.275 214.320 2250.565 214.490 ;
        RECT 2250.735 214.320 2251.025 214.490 ;
        RECT 2251.195 214.320 2251.485 214.490 ;
        RECT 2251.655 214.320 2251.945 214.490 ;
        RECT 2252.115 214.320 2252.405 214.490 ;
        RECT 2252.575 214.320 2252.865 214.490 ;
        RECT 2253.035 214.320 2253.325 214.490 ;
        RECT 2253.495 214.320 2253.785 214.490 ;
        RECT 2253.955 214.320 2254.245 214.490 ;
        RECT 2254.415 214.320 2254.705 214.490 ;
        RECT 2254.875 214.320 2255.165 214.490 ;
        RECT 2255.335 214.320 2255.625 214.490 ;
        RECT 2255.795 214.320 2256.085 214.490 ;
        RECT 2256.255 214.320 2256.545 214.490 ;
        RECT 2256.715 214.320 2257.005 214.490 ;
        RECT 2257.175 214.320 2257.465 214.490 ;
        RECT 2257.635 214.320 2257.925 214.490 ;
        RECT 2258.095 214.320 2258.385 214.490 ;
        RECT 2258.555 214.320 2258.845 214.490 ;
        RECT 2259.015 214.320 2259.305 214.490 ;
        RECT 2259.475 214.320 2259.765 214.490 ;
        RECT 2259.935 214.320 2260.225 214.490 ;
        RECT 2260.395 214.320 2260.685 214.490 ;
        RECT 2260.855 214.320 2261.145 214.490 ;
        RECT 2261.315 214.320 2261.605 214.490 ;
        RECT 2261.775 214.320 2262.065 214.490 ;
        RECT 2262.235 214.320 2262.525 214.490 ;
        RECT 2262.695 214.320 2262.985 214.490 ;
        RECT 2263.155 214.320 2263.445 214.490 ;
        RECT 2263.615 214.320 2263.905 214.490 ;
        RECT 2264.075 214.320 2264.365 214.490 ;
        RECT 2264.535 214.320 2264.825 214.490 ;
        RECT 2264.995 214.320 2265.285 214.490 ;
        RECT 2265.455 214.320 2265.745 214.490 ;
        RECT 2265.915 214.320 2266.205 214.490 ;
        RECT 2266.375 214.320 2266.665 214.490 ;
        RECT 2266.835 214.320 2267.125 214.490 ;
        RECT 2267.295 214.320 2267.585 214.490 ;
        RECT 2267.755 214.320 2268.045 214.490 ;
        RECT 2268.215 214.320 2268.505 214.490 ;
        RECT 2268.675 214.320 2268.965 214.490 ;
        RECT 2269.135 214.320 2269.425 214.490 ;
        RECT 2269.595 214.320 2269.885 214.490 ;
        RECT 2270.055 214.320 2270.345 214.490 ;
        RECT 2270.515 214.320 2270.805 214.490 ;
        RECT 2270.975 214.320 2271.265 214.490 ;
        RECT 2271.435 214.320 2271.725 214.490 ;
        RECT 2271.895 214.320 2272.040 214.490 ;
        RECT 669.085 213.155 669.375 214.320 ;
      LAYER li1 ;
        RECT 669.545 213.885 674.890 214.320 ;
        RECT 672.950 212.635 673.300 213.885 ;
      LAYER li1 ;
        RECT 675.065 213.155 675.355 214.320 ;
        RECT 675.535 213.300 675.865 214.150 ;
        RECT 676.035 213.520 676.205 214.320 ;
        RECT 676.375 213.300 676.705 214.150 ;
        RECT 676.875 213.520 677.045 214.320 ;
      LAYER li1 ;
        RECT 677.295 213.300 677.465 214.150 ;
      LAYER li1 ;
        RECT 677.635 213.520 677.965 214.320 ;
      LAYER li1 ;
        RECT 678.135 213.300 678.305 214.150 ;
      LAYER li1 ;
        RECT 678.475 213.520 678.805 214.320 ;
      LAYER li1 ;
        RECT 678.975 213.300 679.145 214.150 ;
      LAYER li1 ;
        RECT 679.315 213.520 679.645 214.320 ;
      LAYER li1 ;
        RECT 679.815 213.300 679.985 214.150 ;
      LAYER li1 ;
        RECT 675.535 213.130 677.035 213.300 ;
      LAYER li1 ;
        RECT 677.295 213.130 679.985 213.300 ;
      LAYER li1 ;
        RECT 680.155 213.170 680.485 214.320 ;
        RECT 681.045 213.155 681.335 214.320 ;
        RECT 681.515 213.300 681.845 214.150 ;
        RECT 682.015 213.520 682.185 214.320 ;
        RECT 682.355 213.300 682.685 214.150 ;
        RECT 682.855 213.520 683.025 214.320 ;
      LAYER li1 ;
        RECT 683.275 213.300 683.445 214.150 ;
      LAYER li1 ;
        RECT 683.615 213.520 683.945 214.320 ;
      LAYER li1 ;
        RECT 684.115 213.300 684.285 214.150 ;
      LAYER li1 ;
        RECT 684.455 213.520 684.785 214.320 ;
      LAYER li1 ;
        RECT 684.955 213.300 685.125 214.150 ;
      LAYER li1 ;
        RECT 685.295 213.520 685.625 214.320 ;
      LAYER li1 ;
        RECT 685.795 213.300 685.965 214.150 ;
      LAYER li1 ;
        RECT 681.515 213.130 683.015 213.300 ;
      LAYER li1 ;
        RECT 683.275 213.130 685.965 213.300 ;
      LAYER li1 ;
        RECT 686.135 213.170 686.465 214.320 ;
        RECT 687.025 213.155 687.315 214.320 ;
        RECT 687.495 213.300 687.825 214.150 ;
        RECT 687.995 213.520 688.165 214.320 ;
        RECT 688.335 213.300 688.665 214.150 ;
        RECT 688.835 213.520 689.005 214.320 ;
      LAYER li1 ;
        RECT 689.255 213.300 689.425 214.150 ;
      LAYER li1 ;
        RECT 689.595 213.520 689.925 214.320 ;
      LAYER li1 ;
        RECT 690.095 213.300 690.265 214.150 ;
      LAYER li1 ;
        RECT 690.435 213.520 690.765 214.320 ;
      LAYER li1 ;
        RECT 690.935 213.300 691.105 214.150 ;
      LAYER li1 ;
        RECT 691.275 213.520 691.605 214.320 ;
      LAYER li1 ;
        RECT 691.775 213.300 691.945 214.150 ;
      LAYER li1 ;
        RECT 687.495 213.130 688.995 213.300 ;
      LAYER li1 ;
        RECT 689.255 213.130 691.945 213.300 ;
      LAYER li1 ;
        RECT 692.115 213.170 692.445 214.320 ;
        RECT 693.005 213.155 693.295 214.320 ;
        RECT 693.475 213.300 693.805 214.150 ;
        RECT 693.975 213.520 694.145 214.320 ;
        RECT 694.315 213.300 694.645 214.150 ;
        RECT 694.815 213.520 694.985 214.320 ;
      LAYER li1 ;
        RECT 695.235 213.300 695.405 214.150 ;
      LAYER li1 ;
        RECT 695.575 213.520 695.905 214.320 ;
      LAYER li1 ;
        RECT 696.075 213.300 696.245 214.150 ;
      LAYER li1 ;
        RECT 696.415 213.520 696.745 214.320 ;
      LAYER li1 ;
        RECT 696.915 213.300 697.085 214.150 ;
      LAYER li1 ;
        RECT 697.255 213.520 697.585 214.320 ;
      LAYER li1 ;
        RECT 697.755 213.300 697.925 214.150 ;
      LAYER li1 ;
        RECT 693.475 213.130 694.975 213.300 ;
      LAYER li1 ;
        RECT 695.235 213.130 697.925 213.300 ;
      LAYER li1 ;
        RECT 698.095 213.170 698.425 214.320 ;
        RECT 698.985 213.155 699.275 214.320 ;
        RECT 699.455 213.300 699.785 214.150 ;
        RECT 699.955 213.520 700.125 214.320 ;
        RECT 700.295 213.300 700.625 214.150 ;
        RECT 700.795 213.520 700.965 214.320 ;
      LAYER li1 ;
        RECT 701.215 213.300 701.385 214.150 ;
      LAYER li1 ;
        RECT 701.555 213.520 701.885 214.320 ;
      LAYER li1 ;
        RECT 702.055 213.300 702.225 214.150 ;
      LAYER li1 ;
        RECT 702.395 213.520 702.725 214.320 ;
      LAYER li1 ;
        RECT 702.895 213.300 703.065 214.150 ;
      LAYER li1 ;
        RECT 703.235 213.520 703.565 214.320 ;
      LAYER li1 ;
        RECT 703.735 213.300 703.905 214.150 ;
      LAYER li1 ;
        RECT 699.455 213.130 700.955 213.300 ;
      LAYER li1 ;
        RECT 701.215 213.130 703.905 213.300 ;
      LAYER li1 ;
        RECT 704.075 213.170 704.405 214.320 ;
        RECT 704.965 213.155 705.255 214.320 ;
        RECT 705.435 213.300 705.765 214.150 ;
        RECT 705.935 213.520 706.105 214.320 ;
        RECT 706.275 213.300 706.605 214.150 ;
        RECT 706.775 213.520 706.945 214.320 ;
      LAYER li1 ;
        RECT 707.195 213.300 707.365 214.150 ;
      LAYER li1 ;
        RECT 707.535 213.520 707.865 214.320 ;
      LAYER li1 ;
        RECT 708.035 213.300 708.205 214.150 ;
      LAYER li1 ;
        RECT 708.375 213.520 708.705 214.320 ;
      LAYER li1 ;
        RECT 708.875 213.300 709.045 214.150 ;
      LAYER li1 ;
        RECT 709.215 213.520 709.545 214.320 ;
      LAYER li1 ;
        RECT 709.715 213.300 709.885 214.150 ;
      LAYER li1 ;
        RECT 705.435 213.130 706.935 213.300 ;
      LAYER li1 ;
        RECT 707.195 213.130 709.885 213.300 ;
      LAYER li1 ;
        RECT 710.055 213.170 710.385 214.320 ;
        RECT 710.945 213.155 711.235 214.320 ;
        RECT 711.415 213.300 711.745 214.150 ;
        RECT 711.915 213.520 712.085 214.320 ;
        RECT 712.255 213.300 712.585 214.150 ;
        RECT 712.755 213.520 712.925 214.320 ;
      LAYER li1 ;
        RECT 713.175 213.300 713.345 214.150 ;
      LAYER li1 ;
        RECT 713.515 213.520 713.845 214.320 ;
      LAYER li1 ;
        RECT 714.015 213.300 714.185 214.150 ;
      LAYER li1 ;
        RECT 714.355 213.520 714.685 214.320 ;
      LAYER li1 ;
        RECT 714.855 213.300 715.025 214.150 ;
      LAYER li1 ;
        RECT 715.195 213.520 715.525 214.320 ;
      LAYER li1 ;
        RECT 715.695 213.300 715.865 214.150 ;
      LAYER li1 ;
        RECT 711.415 213.130 712.915 213.300 ;
      LAYER li1 ;
        RECT 713.175 213.130 715.865 213.300 ;
      LAYER li1 ;
        RECT 716.035 213.170 716.365 214.320 ;
        RECT 716.925 213.155 717.215 214.320 ;
        RECT 717.395 213.300 717.725 214.150 ;
        RECT 717.895 213.520 718.065 214.320 ;
        RECT 718.235 213.300 718.565 214.150 ;
        RECT 718.735 213.520 718.905 214.320 ;
      LAYER li1 ;
        RECT 719.155 213.300 719.325 214.150 ;
      LAYER li1 ;
        RECT 719.495 213.520 719.825 214.320 ;
      LAYER li1 ;
        RECT 719.995 213.300 720.165 214.150 ;
      LAYER li1 ;
        RECT 720.335 213.520 720.665 214.320 ;
      LAYER li1 ;
        RECT 720.835 213.300 721.005 214.150 ;
      LAYER li1 ;
        RECT 721.175 213.520 721.505 214.320 ;
      LAYER li1 ;
        RECT 721.675 213.300 721.845 214.150 ;
      LAYER li1 ;
        RECT 717.395 213.130 718.895 213.300 ;
      LAYER li1 ;
        RECT 719.155 213.130 721.845 213.300 ;
      LAYER li1 ;
        RECT 722.015 213.170 722.345 214.320 ;
        RECT 722.905 213.155 723.195 214.320 ;
        RECT 723.375 213.300 723.705 214.150 ;
        RECT 723.875 213.520 724.045 214.320 ;
        RECT 724.215 213.300 724.545 214.150 ;
        RECT 724.715 213.520 724.885 214.320 ;
      LAYER li1 ;
        RECT 725.135 213.300 725.305 214.150 ;
      LAYER li1 ;
        RECT 725.475 213.520 725.805 214.320 ;
      LAYER li1 ;
        RECT 725.975 213.300 726.145 214.150 ;
      LAYER li1 ;
        RECT 726.315 213.520 726.645 214.320 ;
      LAYER li1 ;
        RECT 726.815 213.300 726.985 214.150 ;
      LAYER li1 ;
        RECT 727.155 213.520 727.485 214.320 ;
      LAYER li1 ;
        RECT 727.655 213.300 727.825 214.150 ;
      LAYER li1 ;
        RECT 723.375 213.130 724.875 213.300 ;
      LAYER li1 ;
        RECT 725.135 213.130 727.825 213.300 ;
      LAYER li1 ;
        RECT 727.995 213.170 728.325 214.320 ;
        RECT 728.885 213.155 729.175 214.320 ;
        RECT 729.355 213.300 729.685 214.150 ;
        RECT 729.855 213.520 730.025 214.320 ;
        RECT 730.195 213.300 730.525 214.150 ;
        RECT 730.695 213.520 730.865 214.320 ;
      LAYER li1 ;
        RECT 731.115 213.300 731.285 214.150 ;
      LAYER li1 ;
        RECT 731.455 213.520 731.785 214.320 ;
      LAYER li1 ;
        RECT 731.955 213.300 732.125 214.150 ;
      LAYER li1 ;
        RECT 732.295 213.520 732.625 214.320 ;
      LAYER li1 ;
        RECT 732.795 213.300 732.965 214.150 ;
      LAYER li1 ;
        RECT 733.135 213.520 733.465 214.320 ;
      LAYER li1 ;
        RECT 733.635 213.300 733.805 214.150 ;
      LAYER li1 ;
        RECT 729.355 213.130 730.855 213.300 ;
      LAYER li1 ;
        RECT 731.115 213.130 733.805 213.300 ;
      LAYER li1 ;
        RECT 733.975 213.170 734.305 214.320 ;
        RECT 734.865 213.155 735.155 214.320 ;
        RECT 735.335 213.300 735.665 214.150 ;
        RECT 735.835 213.520 736.005 214.320 ;
        RECT 736.175 213.300 736.505 214.150 ;
        RECT 736.675 213.520 736.845 214.320 ;
      LAYER li1 ;
        RECT 737.095 213.300 737.265 214.150 ;
      LAYER li1 ;
        RECT 737.435 213.520 737.765 214.320 ;
      LAYER li1 ;
        RECT 737.935 213.300 738.105 214.150 ;
      LAYER li1 ;
        RECT 738.275 213.520 738.605 214.320 ;
      LAYER li1 ;
        RECT 738.775 213.300 738.945 214.150 ;
      LAYER li1 ;
        RECT 739.115 213.520 739.445 214.320 ;
      LAYER li1 ;
        RECT 739.615 213.300 739.785 214.150 ;
      LAYER li1 ;
        RECT 735.335 213.130 736.835 213.300 ;
      LAYER li1 ;
        RECT 737.095 213.130 739.785 213.300 ;
      LAYER li1 ;
        RECT 739.955 213.170 740.285 214.320 ;
        RECT 740.845 213.155 741.135 214.320 ;
        RECT 741.315 213.300 741.645 214.150 ;
        RECT 741.815 213.520 741.985 214.320 ;
        RECT 742.155 213.300 742.485 214.150 ;
        RECT 742.655 213.520 742.825 214.320 ;
      LAYER li1 ;
        RECT 743.075 213.300 743.245 214.150 ;
      LAYER li1 ;
        RECT 743.415 213.520 743.745 214.320 ;
      LAYER li1 ;
        RECT 743.915 213.300 744.085 214.150 ;
      LAYER li1 ;
        RECT 744.255 213.520 744.585 214.320 ;
      LAYER li1 ;
        RECT 744.755 213.300 744.925 214.150 ;
      LAYER li1 ;
        RECT 745.095 213.520 745.425 214.320 ;
      LAYER li1 ;
        RECT 745.595 213.300 745.765 214.150 ;
      LAYER li1 ;
        RECT 741.315 213.130 742.815 213.300 ;
      LAYER li1 ;
        RECT 743.075 213.130 745.765 213.300 ;
      LAYER li1 ;
        RECT 745.935 213.170 746.265 214.320 ;
        RECT 746.825 213.155 747.115 214.320 ;
        RECT 747.295 213.300 747.625 214.150 ;
        RECT 747.795 213.520 747.965 214.320 ;
        RECT 748.135 213.300 748.465 214.150 ;
        RECT 748.635 213.520 748.805 214.320 ;
      LAYER li1 ;
        RECT 749.055 213.300 749.225 214.150 ;
      LAYER li1 ;
        RECT 749.395 213.520 749.725 214.320 ;
      LAYER li1 ;
        RECT 749.895 213.300 750.065 214.150 ;
      LAYER li1 ;
        RECT 750.235 213.520 750.565 214.320 ;
      LAYER li1 ;
        RECT 750.735 213.300 750.905 214.150 ;
      LAYER li1 ;
        RECT 751.075 213.520 751.405 214.320 ;
      LAYER li1 ;
        RECT 751.575 213.300 751.745 214.150 ;
      LAYER li1 ;
        RECT 747.295 213.130 748.795 213.300 ;
      LAYER li1 ;
        RECT 749.055 213.130 751.745 213.300 ;
      LAYER li1 ;
        RECT 751.915 213.170 752.245 214.320 ;
        RECT 752.805 213.155 753.095 214.320 ;
        RECT 753.275 213.300 753.605 214.150 ;
        RECT 753.775 213.520 753.945 214.320 ;
        RECT 754.115 213.300 754.445 214.150 ;
        RECT 754.615 213.520 754.785 214.320 ;
      LAYER li1 ;
        RECT 755.035 213.300 755.205 214.150 ;
      LAYER li1 ;
        RECT 755.375 213.520 755.705 214.320 ;
      LAYER li1 ;
        RECT 755.875 213.300 756.045 214.150 ;
      LAYER li1 ;
        RECT 756.215 213.520 756.545 214.320 ;
      LAYER li1 ;
        RECT 756.715 213.300 756.885 214.150 ;
      LAYER li1 ;
        RECT 757.055 213.520 757.385 214.320 ;
      LAYER li1 ;
        RECT 757.555 213.300 757.725 214.150 ;
      LAYER li1 ;
        RECT 753.275 213.130 754.775 213.300 ;
      LAYER li1 ;
        RECT 755.035 213.130 757.725 213.300 ;
      LAYER li1 ;
        RECT 757.895 213.170 758.225 214.320 ;
        RECT 758.785 213.155 759.075 214.320 ;
        RECT 759.255 213.300 759.585 214.150 ;
        RECT 759.755 213.520 759.925 214.320 ;
        RECT 760.095 213.300 760.425 214.150 ;
        RECT 760.595 213.520 760.765 214.320 ;
      LAYER li1 ;
        RECT 761.015 213.300 761.185 214.150 ;
      LAYER li1 ;
        RECT 761.355 213.520 761.685 214.320 ;
      LAYER li1 ;
        RECT 761.855 213.300 762.025 214.150 ;
      LAYER li1 ;
        RECT 762.195 213.520 762.525 214.320 ;
      LAYER li1 ;
        RECT 762.695 213.300 762.865 214.150 ;
      LAYER li1 ;
        RECT 763.035 213.520 763.365 214.320 ;
      LAYER li1 ;
        RECT 763.535 213.300 763.705 214.150 ;
      LAYER li1 ;
        RECT 759.255 213.130 760.755 213.300 ;
      LAYER li1 ;
        RECT 761.015 213.130 763.705 213.300 ;
      LAYER li1 ;
        RECT 763.875 213.170 764.205 214.320 ;
        RECT 764.765 213.155 765.055 214.320 ;
        RECT 765.235 213.300 765.565 214.150 ;
        RECT 765.735 213.520 765.905 214.320 ;
        RECT 766.075 213.300 766.405 214.150 ;
        RECT 766.575 213.520 766.745 214.320 ;
      LAYER li1 ;
        RECT 766.995 213.300 767.165 214.150 ;
      LAYER li1 ;
        RECT 767.335 213.520 767.665 214.320 ;
      LAYER li1 ;
        RECT 767.835 213.300 768.005 214.150 ;
      LAYER li1 ;
        RECT 768.175 213.520 768.505 214.320 ;
      LAYER li1 ;
        RECT 768.675 213.300 768.845 214.150 ;
      LAYER li1 ;
        RECT 769.015 213.520 769.345 214.320 ;
      LAYER li1 ;
        RECT 769.515 213.300 769.685 214.150 ;
      LAYER li1 ;
        RECT 765.235 213.130 766.735 213.300 ;
      LAYER li1 ;
        RECT 766.995 213.130 769.685 213.300 ;
      LAYER li1 ;
        RECT 769.855 213.170 770.185 214.320 ;
        RECT 770.745 213.155 771.035 214.320 ;
        RECT 771.215 213.300 771.545 214.150 ;
        RECT 771.715 213.520 771.885 214.320 ;
        RECT 772.055 213.300 772.385 214.150 ;
        RECT 772.555 213.520 772.725 214.320 ;
      LAYER li1 ;
        RECT 772.975 213.300 773.145 214.150 ;
      LAYER li1 ;
        RECT 773.315 213.520 773.645 214.320 ;
      LAYER li1 ;
        RECT 773.815 213.300 773.985 214.150 ;
      LAYER li1 ;
        RECT 774.155 213.520 774.485 214.320 ;
      LAYER li1 ;
        RECT 774.655 213.300 774.825 214.150 ;
      LAYER li1 ;
        RECT 774.995 213.520 775.325 214.320 ;
      LAYER li1 ;
        RECT 775.495 213.300 775.665 214.150 ;
      LAYER li1 ;
        RECT 771.215 213.130 772.715 213.300 ;
      LAYER li1 ;
        RECT 772.975 213.130 775.665 213.300 ;
      LAYER li1 ;
        RECT 775.835 213.170 776.165 214.320 ;
        RECT 776.725 213.155 777.015 214.320 ;
        RECT 777.195 213.300 777.525 214.150 ;
        RECT 777.695 213.520 777.865 214.320 ;
        RECT 778.035 213.300 778.365 214.150 ;
        RECT 778.535 213.520 778.705 214.320 ;
      LAYER li1 ;
        RECT 778.955 213.300 779.125 214.150 ;
      LAYER li1 ;
        RECT 779.295 213.520 779.625 214.320 ;
      LAYER li1 ;
        RECT 779.795 213.300 779.965 214.150 ;
      LAYER li1 ;
        RECT 780.135 213.520 780.465 214.320 ;
      LAYER li1 ;
        RECT 780.635 213.300 780.805 214.150 ;
      LAYER li1 ;
        RECT 780.975 213.520 781.305 214.320 ;
      LAYER li1 ;
        RECT 781.475 213.300 781.645 214.150 ;
      LAYER li1 ;
        RECT 777.195 213.130 778.695 213.300 ;
      LAYER li1 ;
        RECT 778.955 213.130 781.645 213.300 ;
      LAYER li1 ;
        RECT 781.815 213.170 782.145 214.320 ;
        RECT 782.705 213.155 782.995 214.320 ;
        RECT 783.175 213.300 783.505 214.150 ;
        RECT 783.675 213.520 783.845 214.320 ;
        RECT 784.015 213.300 784.345 214.150 ;
        RECT 784.515 213.520 784.685 214.320 ;
      LAYER li1 ;
        RECT 784.935 213.300 785.105 214.150 ;
      LAYER li1 ;
        RECT 785.275 213.520 785.605 214.320 ;
      LAYER li1 ;
        RECT 785.775 213.300 785.945 214.150 ;
      LAYER li1 ;
        RECT 786.115 213.520 786.445 214.320 ;
      LAYER li1 ;
        RECT 786.615 213.300 786.785 214.150 ;
      LAYER li1 ;
        RECT 786.955 213.520 787.285 214.320 ;
      LAYER li1 ;
        RECT 787.455 213.300 787.625 214.150 ;
      LAYER li1 ;
        RECT 783.175 213.130 784.675 213.300 ;
      LAYER li1 ;
        RECT 784.935 213.130 787.625 213.300 ;
      LAYER li1 ;
        RECT 787.795 213.170 788.125 214.320 ;
        RECT 788.685 213.155 788.975 214.320 ;
        RECT 789.535 213.170 789.865 214.320 ;
        RECT 790.375 213.520 790.705 214.320 ;
        RECT 791.215 213.520 791.545 214.320 ;
        RECT 792.055 213.520 792.385 214.320 ;
        RECT 792.975 213.520 793.145 214.320 ;
        RECT 793.315 213.300 793.645 214.150 ;
        RECT 793.815 213.520 793.985 214.320 ;
        RECT 794.155 213.300 794.485 214.150 ;
      LAYER li1 ;
        RECT 675.580 212.760 676.680 212.960 ;
      LAYER li1 ;
        RECT 676.860 212.930 677.035 213.130 ;
        RECT 676.860 212.760 679.485 212.930 ;
        RECT 676.860 212.590 677.035 212.760 ;
      LAYER li1 ;
        RECT 679.730 212.590 679.985 213.130 ;
        RECT 681.560 212.760 682.660 212.960 ;
      LAYER li1 ;
        RECT 682.840 212.930 683.015 213.130 ;
        RECT 682.840 212.760 685.465 212.930 ;
        RECT 682.840 212.590 683.015 212.760 ;
      LAYER li1 ;
        RECT 685.710 212.590 685.965 213.130 ;
        RECT 687.540 212.760 688.640 212.960 ;
      LAYER li1 ;
        RECT 688.820 212.930 688.995 213.130 ;
        RECT 688.820 212.760 691.445 212.930 ;
        RECT 688.820 212.590 688.995 212.760 ;
      LAYER li1 ;
        RECT 691.690 212.590 691.945 213.130 ;
        RECT 693.520 212.760 694.620 212.960 ;
      LAYER li1 ;
        RECT 694.800 212.930 694.975 213.130 ;
        RECT 694.800 212.760 697.425 212.930 ;
        RECT 694.800 212.590 694.975 212.760 ;
      LAYER li1 ;
        RECT 697.670 212.590 697.925 213.130 ;
        RECT 699.500 212.760 700.600 212.960 ;
      LAYER li1 ;
        RECT 700.780 212.930 700.955 213.130 ;
        RECT 700.780 212.760 703.405 212.930 ;
        RECT 700.780 212.590 700.955 212.760 ;
      LAYER li1 ;
        RECT 703.650 212.590 703.905 213.130 ;
        RECT 705.480 212.760 706.580 212.960 ;
      LAYER li1 ;
        RECT 706.760 212.930 706.935 213.130 ;
        RECT 706.760 212.760 709.385 212.930 ;
        RECT 706.760 212.590 706.935 212.760 ;
      LAYER li1 ;
        RECT 709.630 212.590 709.885 213.130 ;
        RECT 711.460 212.760 712.560 212.960 ;
      LAYER li1 ;
        RECT 712.740 212.930 712.915 213.130 ;
        RECT 712.740 212.760 715.365 212.930 ;
        RECT 712.740 212.590 712.915 212.760 ;
      LAYER li1 ;
        RECT 715.610 212.590 715.865 213.130 ;
        RECT 717.440 212.760 718.540 212.960 ;
      LAYER li1 ;
        RECT 718.720 212.930 718.895 213.130 ;
        RECT 718.720 212.760 721.345 212.930 ;
        RECT 718.720 212.590 718.895 212.760 ;
      LAYER li1 ;
        RECT 721.590 212.590 721.845 213.130 ;
        RECT 723.420 212.760 724.520 212.960 ;
      LAYER li1 ;
        RECT 724.700 212.930 724.875 213.130 ;
        RECT 724.700 212.760 727.325 212.930 ;
        RECT 724.700 212.590 724.875 212.760 ;
      LAYER li1 ;
        RECT 727.570 212.590 727.825 213.130 ;
        RECT 729.400 212.760 730.500 212.960 ;
      LAYER li1 ;
        RECT 730.680 212.930 730.855 213.130 ;
        RECT 730.680 212.760 733.305 212.930 ;
        RECT 730.680 212.590 730.855 212.760 ;
      LAYER li1 ;
        RECT 733.550 212.590 733.805 213.130 ;
        RECT 735.380 212.760 736.480 212.960 ;
      LAYER li1 ;
        RECT 736.660 212.930 736.835 213.130 ;
        RECT 736.660 212.760 739.285 212.930 ;
        RECT 736.660 212.590 736.835 212.760 ;
      LAYER li1 ;
        RECT 739.530 212.590 739.785 213.130 ;
        RECT 741.360 212.760 742.460 212.960 ;
      LAYER li1 ;
        RECT 742.640 212.930 742.815 213.130 ;
        RECT 742.640 212.760 745.265 212.930 ;
        RECT 742.640 212.590 742.815 212.760 ;
      LAYER li1 ;
        RECT 745.510 212.590 745.765 213.130 ;
        RECT 747.340 212.760 748.440 212.960 ;
      LAYER li1 ;
        RECT 748.620 212.930 748.795 213.130 ;
        RECT 748.620 212.760 751.245 212.930 ;
        RECT 748.620 212.590 748.795 212.760 ;
      LAYER li1 ;
        RECT 751.490 212.590 751.745 213.130 ;
        RECT 753.320 212.760 754.420 212.960 ;
      LAYER li1 ;
        RECT 754.600 212.930 754.775 213.130 ;
        RECT 754.600 212.760 757.225 212.930 ;
        RECT 754.600 212.590 754.775 212.760 ;
      LAYER li1 ;
        RECT 757.470 212.590 757.725 213.130 ;
        RECT 759.300 212.760 760.400 212.960 ;
      LAYER li1 ;
        RECT 760.580 212.930 760.755 213.130 ;
        RECT 760.580 212.760 763.205 212.930 ;
        RECT 760.580 212.590 760.755 212.760 ;
      LAYER li1 ;
        RECT 763.450 212.590 763.705 213.130 ;
      LAYER li1 ;
        RECT 766.560 212.930 766.735 213.130 ;
        RECT 766.560 212.760 769.185 212.930 ;
        RECT 766.560 212.590 766.735 212.760 ;
      LAYER li1 ;
        RECT 769.430 212.590 769.685 213.130 ;
      LAYER li1 ;
        RECT 772.540 212.930 772.715 213.130 ;
        RECT 772.540 212.760 775.165 212.930 ;
        RECT 772.540 212.590 772.715 212.760 ;
      LAYER li1 ;
        RECT 775.410 212.590 775.665 213.130 ;
      LAYER li1 ;
        RECT 778.520 212.930 778.695 213.130 ;
        RECT 778.520 212.760 781.145 212.930 ;
        RECT 778.520 212.590 778.695 212.760 ;
      LAYER li1 ;
        RECT 781.390 212.590 781.645 213.130 ;
      LAYER li1 ;
        RECT 784.500 212.930 784.675 213.130 ;
        RECT 784.500 212.760 787.125 212.930 ;
        RECT 784.500 212.590 784.675 212.760 ;
      LAYER li1 ;
        RECT 787.370 212.590 787.625 213.130 ;
      LAYER li1 ;
        RECT 792.985 213.130 794.485 213.300 ;
        RECT 794.665 213.155 794.955 214.320 ;
        RECT 2146.085 213.155 2146.375 214.320 ;
      LAYER li1 ;
        RECT 2146.545 213.885 2151.890 214.320 ;
      LAYER li1 ;
        RECT 792.985 212.930 793.160 213.130 ;
        RECT 790.535 212.760 793.160 212.930 ;
      LAYER li1 ;
        RECT 793.340 212.760 794.440 212.960 ;
      LAYER li1 ;
        RECT 669.085 211.770 669.375 212.495 ;
        RECT 675.065 211.770 675.355 212.495 ;
        RECT 675.615 212.420 677.035 212.590 ;
      LAYER li1 ;
        RECT 677.295 212.420 679.985 212.590 ;
      LAYER li1 ;
        RECT 675.615 211.940 675.785 212.420 ;
        RECT 675.955 211.770 676.285 212.250 ;
        RECT 676.455 211.945 676.625 212.420 ;
        RECT 676.795 211.770 677.125 212.250 ;
      LAYER li1 ;
        RECT 677.295 211.940 677.465 212.420 ;
      LAYER li1 ;
        RECT 677.635 211.770 677.965 212.250 ;
      LAYER li1 ;
        RECT 678.135 211.940 678.305 212.420 ;
      LAYER li1 ;
        RECT 678.475 211.770 678.805 212.250 ;
      LAYER li1 ;
        RECT 678.975 211.940 679.145 212.420 ;
      LAYER li1 ;
        RECT 679.315 211.770 679.645 212.250 ;
      LAYER li1 ;
        RECT 679.815 211.940 679.985 212.420 ;
      LAYER li1 ;
        RECT 680.155 211.770 680.485 212.570 ;
        RECT 681.045 211.770 681.335 212.495 ;
        RECT 681.595 212.420 683.015 212.590 ;
      LAYER li1 ;
        RECT 683.275 212.420 685.965 212.590 ;
      LAYER li1 ;
        RECT 681.595 211.940 681.765 212.420 ;
        RECT 681.935 211.770 682.265 212.250 ;
        RECT 682.435 211.945 682.605 212.420 ;
        RECT 682.775 211.770 683.105 212.250 ;
      LAYER li1 ;
        RECT 683.275 211.940 683.445 212.420 ;
      LAYER li1 ;
        RECT 683.615 211.770 683.945 212.250 ;
      LAYER li1 ;
        RECT 684.115 211.940 684.285 212.420 ;
      LAYER li1 ;
        RECT 684.455 211.770 684.785 212.250 ;
      LAYER li1 ;
        RECT 684.955 211.940 685.125 212.420 ;
      LAYER li1 ;
        RECT 685.295 211.770 685.625 212.250 ;
      LAYER li1 ;
        RECT 685.795 211.940 685.965 212.420 ;
      LAYER li1 ;
        RECT 686.135 211.770 686.465 212.570 ;
        RECT 687.025 211.770 687.315 212.495 ;
        RECT 687.575 212.420 688.995 212.590 ;
      LAYER li1 ;
        RECT 689.255 212.420 691.945 212.590 ;
      LAYER li1 ;
        RECT 687.575 211.940 687.745 212.420 ;
        RECT 687.915 211.770 688.245 212.250 ;
        RECT 688.415 211.945 688.585 212.420 ;
        RECT 688.755 211.770 689.085 212.250 ;
      LAYER li1 ;
        RECT 689.255 211.940 689.425 212.420 ;
      LAYER li1 ;
        RECT 689.595 211.770 689.925 212.250 ;
      LAYER li1 ;
        RECT 690.095 211.940 690.265 212.420 ;
      LAYER li1 ;
        RECT 690.435 211.770 690.765 212.250 ;
      LAYER li1 ;
        RECT 690.935 211.940 691.105 212.420 ;
      LAYER li1 ;
        RECT 691.275 211.770 691.605 212.250 ;
      LAYER li1 ;
        RECT 691.775 211.940 691.945 212.420 ;
      LAYER li1 ;
        RECT 692.115 211.770 692.445 212.570 ;
        RECT 693.005 211.770 693.295 212.495 ;
        RECT 693.555 212.420 694.975 212.590 ;
      LAYER li1 ;
        RECT 695.235 212.420 697.925 212.590 ;
      LAYER li1 ;
        RECT 693.555 211.940 693.725 212.420 ;
        RECT 693.895 211.770 694.225 212.250 ;
        RECT 694.395 211.945 694.565 212.420 ;
        RECT 694.735 211.770 695.065 212.250 ;
      LAYER li1 ;
        RECT 695.235 211.940 695.405 212.420 ;
      LAYER li1 ;
        RECT 695.575 211.770 695.905 212.250 ;
      LAYER li1 ;
        RECT 696.075 211.940 696.245 212.420 ;
      LAYER li1 ;
        RECT 696.415 211.770 696.745 212.250 ;
      LAYER li1 ;
        RECT 696.915 211.940 697.085 212.420 ;
      LAYER li1 ;
        RECT 697.255 211.770 697.585 212.250 ;
      LAYER li1 ;
        RECT 697.755 211.940 697.925 212.420 ;
      LAYER li1 ;
        RECT 698.095 211.770 698.425 212.570 ;
        RECT 698.985 211.770 699.275 212.495 ;
        RECT 699.535 212.420 700.955 212.590 ;
      LAYER li1 ;
        RECT 701.215 212.420 703.905 212.590 ;
      LAYER li1 ;
        RECT 699.535 211.940 699.705 212.420 ;
        RECT 699.875 211.770 700.205 212.250 ;
        RECT 700.375 211.945 700.545 212.420 ;
        RECT 700.715 211.770 701.045 212.250 ;
      LAYER li1 ;
        RECT 701.215 211.940 701.385 212.420 ;
      LAYER li1 ;
        RECT 701.555 211.770 701.885 212.250 ;
      LAYER li1 ;
        RECT 702.055 211.940 702.225 212.420 ;
      LAYER li1 ;
        RECT 702.395 211.770 702.725 212.250 ;
      LAYER li1 ;
        RECT 702.895 211.940 703.065 212.420 ;
      LAYER li1 ;
        RECT 703.235 211.770 703.565 212.250 ;
      LAYER li1 ;
        RECT 703.735 211.940 703.905 212.420 ;
      LAYER li1 ;
        RECT 704.075 211.770 704.405 212.570 ;
        RECT 704.965 211.770 705.255 212.495 ;
        RECT 705.515 212.420 706.935 212.590 ;
      LAYER li1 ;
        RECT 707.195 212.420 709.885 212.590 ;
      LAYER li1 ;
        RECT 705.515 211.940 705.685 212.420 ;
        RECT 705.855 211.770 706.185 212.250 ;
        RECT 706.355 211.945 706.525 212.420 ;
        RECT 706.695 211.770 707.025 212.250 ;
      LAYER li1 ;
        RECT 707.195 211.940 707.365 212.420 ;
      LAYER li1 ;
        RECT 707.535 211.770 707.865 212.250 ;
      LAYER li1 ;
        RECT 708.035 211.940 708.205 212.420 ;
      LAYER li1 ;
        RECT 708.375 211.770 708.705 212.250 ;
      LAYER li1 ;
        RECT 708.875 211.940 709.045 212.420 ;
      LAYER li1 ;
        RECT 709.215 211.770 709.545 212.250 ;
      LAYER li1 ;
        RECT 709.715 211.940 709.885 212.420 ;
      LAYER li1 ;
        RECT 710.055 211.770 710.385 212.570 ;
        RECT 710.945 211.770 711.235 212.495 ;
        RECT 711.495 212.420 712.915 212.590 ;
      LAYER li1 ;
        RECT 713.175 212.420 715.865 212.590 ;
      LAYER li1 ;
        RECT 711.495 211.940 711.665 212.420 ;
        RECT 711.835 211.770 712.165 212.250 ;
        RECT 712.335 211.945 712.505 212.420 ;
        RECT 712.675 211.770 713.005 212.250 ;
      LAYER li1 ;
        RECT 713.175 211.940 713.345 212.420 ;
      LAYER li1 ;
        RECT 713.515 211.770 713.845 212.250 ;
      LAYER li1 ;
        RECT 714.015 211.940 714.185 212.420 ;
      LAYER li1 ;
        RECT 714.355 211.770 714.685 212.250 ;
      LAYER li1 ;
        RECT 714.855 211.940 715.025 212.420 ;
      LAYER li1 ;
        RECT 715.195 211.770 715.525 212.250 ;
      LAYER li1 ;
        RECT 715.695 211.940 715.865 212.420 ;
      LAYER li1 ;
        RECT 716.035 211.770 716.365 212.570 ;
        RECT 716.925 211.770 717.215 212.495 ;
        RECT 717.475 212.420 718.895 212.590 ;
      LAYER li1 ;
        RECT 719.155 212.420 721.845 212.590 ;
      LAYER li1 ;
        RECT 717.475 211.940 717.645 212.420 ;
        RECT 717.815 211.770 718.145 212.250 ;
        RECT 718.315 211.945 718.485 212.420 ;
        RECT 718.655 211.770 718.985 212.250 ;
      LAYER li1 ;
        RECT 719.155 211.940 719.325 212.420 ;
      LAYER li1 ;
        RECT 719.495 211.770 719.825 212.250 ;
      LAYER li1 ;
        RECT 719.995 211.940 720.165 212.420 ;
      LAYER li1 ;
        RECT 720.335 211.770 720.665 212.250 ;
      LAYER li1 ;
        RECT 720.835 211.940 721.005 212.420 ;
      LAYER li1 ;
        RECT 721.175 211.770 721.505 212.250 ;
      LAYER li1 ;
        RECT 721.675 211.940 721.845 212.420 ;
      LAYER li1 ;
        RECT 722.015 211.770 722.345 212.570 ;
        RECT 722.905 211.770 723.195 212.495 ;
        RECT 723.455 212.420 724.875 212.590 ;
      LAYER li1 ;
        RECT 725.135 212.420 727.825 212.590 ;
      LAYER li1 ;
        RECT 723.455 211.940 723.625 212.420 ;
        RECT 723.795 211.770 724.125 212.250 ;
        RECT 724.295 211.945 724.465 212.420 ;
        RECT 724.635 211.770 724.965 212.250 ;
      LAYER li1 ;
        RECT 725.135 211.940 725.305 212.420 ;
      LAYER li1 ;
        RECT 725.475 211.770 725.805 212.250 ;
      LAYER li1 ;
        RECT 725.975 211.940 726.145 212.420 ;
      LAYER li1 ;
        RECT 726.315 211.770 726.645 212.250 ;
      LAYER li1 ;
        RECT 726.815 211.940 726.985 212.420 ;
      LAYER li1 ;
        RECT 727.155 211.770 727.485 212.250 ;
      LAYER li1 ;
        RECT 727.655 211.940 727.825 212.420 ;
      LAYER li1 ;
        RECT 727.995 211.770 728.325 212.570 ;
        RECT 728.885 211.770 729.175 212.495 ;
        RECT 729.435 212.420 730.855 212.590 ;
      LAYER li1 ;
        RECT 731.115 212.420 733.805 212.590 ;
      LAYER li1 ;
        RECT 729.435 211.940 729.605 212.420 ;
        RECT 729.775 211.770 730.105 212.250 ;
        RECT 730.275 211.945 730.445 212.420 ;
        RECT 730.615 211.770 730.945 212.250 ;
      LAYER li1 ;
        RECT 731.115 211.940 731.285 212.420 ;
      LAYER li1 ;
        RECT 731.455 211.770 731.785 212.250 ;
      LAYER li1 ;
        RECT 731.955 211.940 732.125 212.420 ;
      LAYER li1 ;
        RECT 732.295 211.770 732.625 212.250 ;
      LAYER li1 ;
        RECT 732.795 211.940 732.965 212.420 ;
      LAYER li1 ;
        RECT 733.135 211.770 733.465 212.250 ;
      LAYER li1 ;
        RECT 733.635 211.940 733.805 212.420 ;
      LAYER li1 ;
        RECT 733.975 211.770 734.305 212.570 ;
        RECT 734.865 211.770 735.155 212.495 ;
        RECT 735.415 212.420 736.835 212.590 ;
      LAYER li1 ;
        RECT 737.095 212.420 739.785 212.590 ;
      LAYER li1 ;
        RECT 735.415 211.940 735.585 212.420 ;
        RECT 735.755 211.770 736.085 212.250 ;
        RECT 736.255 211.945 736.425 212.420 ;
        RECT 736.595 211.770 736.925 212.250 ;
      LAYER li1 ;
        RECT 737.095 211.940 737.265 212.420 ;
      LAYER li1 ;
        RECT 737.435 211.770 737.765 212.250 ;
      LAYER li1 ;
        RECT 737.935 211.940 738.105 212.420 ;
      LAYER li1 ;
        RECT 738.275 211.770 738.605 212.250 ;
      LAYER li1 ;
        RECT 738.775 211.940 738.945 212.420 ;
      LAYER li1 ;
        RECT 739.115 211.770 739.445 212.250 ;
      LAYER li1 ;
        RECT 739.615 211.940 739.785 212.420 ;
      LAYER li1 ;
        RECT 739.955 211.770 740.285 212.570 ;
        RECT 740.845 211.770 741.135 212.495 ;
        RECT 741.395 212.420 742.815 212.590 ;
      LAYER li1 ;
        RECT 743.075 212.420 745.765 212.590 ;
      LAYER li1 ;
        RECT 741.395 211.940 741.565 212.420 ;
        RECT 741.735 211.770 742.065 212.250 ;
        RECT 742.235 211.945 742.405 212.420 ;
        RECT 742.575 211.770 742.905 212.250 ;
      LAYER li1 ;
        RECT 743.075 211.940 743.245 212.420 ;
      LAYER li1 ;
        RECT 743.415 211.770 743.745 212.250 ;
      LAYER li1 ;
        RECT 743.915 211.940 744.085 212.420 ;
      LAYER li1 ;
        RECT 744.255 211.770 744.585 212.250 ;
      LAYER li1 ;
        RECT 744.755 211.940 744.925 212.420 ;
      LAYER li1 ;
        RECT 745.095 211.770 745.425 212.250 ;
      LAYER li1 ;
        RECT 745.595 211.940 745.765 212.420 ;
      LAYER li1 ;
        RECT 745.935 211.770 746.265 212.570 ;
        RECT 746.825 211.770 747.115 212.495 ;
        RECT 747.375 212.420 748.795 212.590 ;
      LAYER li1 ;
        RECT 749.055 212.420 751.745 212.590 ;
      LAYER li1 ;
        RECT 747.375 211.940 747.545 212.420 ;
        RECT 747.715 211.770 748.045 212.250 ;
        RECT 748.215 211.945 748.385 212.420 ;
        RECT 748.555 211.770 748.885 212.250 ;
      LAYER li1 ;
        RECT 749.055 211.940 749.225 212.420 ;
      LAYER li1 ;
        RECT 749.395 211.770 749.725 212.250 ;
      LAYER li1 ;
        RECT 749.895 211.940 750.065 212.420 ;
      LAYER li1 ;
        RECT 750.235 211.770 750.565 212.250 ;
      LAYER li1 ;
        RECT 750.735 211.940 750.905 212.420 ;
      LAYER li1 ;
        RECT 751.075 211.770 751.405 212.250 ;
      LAYER li1 ;
        RECT 751.575 211.940 751.745 212.420 ;
      LAYER li1 ;
        RECT 751.915 211.770 752.245 212.570 ;
        RECT 752.805 211.770 753.095 212.495 ;
        RECT 753.355 212.420 754.775 212.590 ;
      LAYER li1 ;
        RECT 755.035 212.420 757.725 212.590 ;
      LAYER li1 ;
        RECT 753.355 211.940 753.525 212.420 ;
        RECT 753.695 211.770 754.025 212.250 ;
        RECT 754.195 211.945 754.365 212.420 ;
        RECT 754.535 211.770 754.865 212.250 ;
      LAYER li1 ;
        RECT 755.035 211.940 755.205 212.420 ;
      LAYER li1 ;
        RECT 755.375 211.770 755.705 212.250 ;
      LAYER li1 ;
        RECT 755.875 211.940 756.045 212.420 ;
      LAYER li1 ;
        RECT 756.215 211.770 756.545 212.250 ;
      LAYER li1 ;
        RECT 756.715 211.940 756.885 212.420 ;
      LAYER li1 ;
        RECT 757.055 211.770 757.385 212.250 ;
      LAYER li1 ;
        RECT 757.555 211.940 757.725 212.420 ;
      LAYER li1 ;
        RECT 757.895 211.770 758.225 212.570 ;
        RECT 758.785 211.770 759.075 212.495 ;
        RECT 759.335 212.420 760.755 212.590 ;
      LAYER li1 ;
        RECT 761.015 212.420 763.705 212.590 ;
      LAYER li1 ;
        RECT 759.335 211.940 759.505 212.420 ;
        RECT 759.675 211.770 760.005 212.250 ;
        RECT 760.175 211.945 760.345 212.420 ;
        RECT 760.515 211.770 760.845 212.250 ;
      LAYER li1 ;
        RECT 761.015 211.940 761.185 212.420 ;
      LAYER li1 ;
        RECT 761.355 211.770 761.685 212.250 ;
      LAYER li1 ;
        RECT 761.855 211.940 762.025 212.420 ;
      LAYER li1 ;
        RECT 762.195 211.770 762.525 212.250 ;
      LAYER li1 ;
        RECT 762.695 211.940 762.865 212.420 ;
      LAYER li1 ;
        RECT 763.035 211.770 763.365 212.250 ;
      LAYER li1 ;
        RECT 763.535 211.940 763.705 212.420 ;
      LAYER li1 ;
        RECT 763.875 211.770 764.205 212.570 ;
        RECT 764.765 211.770 765.055 212.495 ;
        RECT 765.315 212.420 766.735 212.590 ;
      LAYER li1 ;
        RECT 766.995 212.420 769.685 212.590 ;
      LAYER li1 ;
        RECT 765.315 211.940 765.485 212.420 ;
        RECT 765.655 211.770 765.985 212.250 ;
        RECT 766.155 211.945 766.325 212.420 ;
        RECT 766.495 211.770 766.825 212.250 ;
      LAYER li1 ;
        RECT 766.995 211.940 767.165 212.420 ;
      LAYER li1 ;
        RECT 767.335 211.770 767.665 212.250 ;
      LAYER li1 ;
        RECT 767.835 211.940 768.005 212.420 ;
      LAYER li1 ;
        RECT 768.175 211.770 768.505 212.250 ;
      LAYER li1 ;
        RECT 768.675 211.940 768.845 212.420 ;
      LAYER li1 ;
        RECT 769.015 211.770 769.345 212.250 ;
      LAYER li1 ;
        RECT 769.515 211.940 769.685 212.420 ;
      LAYER li1 ;
        RECT 769.855 211.770 770.185 212.570 ;
        RECT 770.745 211.770 771.035 212.495 ;
        RECT 771.295 212.420 772.715 212.590 ;
      LAYER li1 ;
        RECT 772.975 212.420 775.665 212.590 ;
      LAYER li1 ;
        RECT 771.295 211.940 771.465 212.420 ;
        RECT 771.635 211.770 771.965 212.250 ;
        RECT 772.135 211.945 772.305 212.420 ;
        RECT 772.475 211.770 772.805 212.250 ;
      LAYER li1 ;
        RECT 772.975 211.940 773.145 212.420 ;
      LAYER li1 ;
        RECT 773.315 211.770 773.645 212.250 ;
      LAYER li1 ;
        RECT 773.815 211.940 773.985 212.420 ;
      LAYER li1 ;
        RECT 774.155 211.770 774.485 212.250 ;
      LAYER li1 ;
        RECT 774.655 211.940 774.825 212.420 ;
      LAYER li1 ;
        RECT 774.995 211.770 775.325 212.250 ;
      LAYER li1 ;
        RECT 775.495 211.940 775.665 212.420 ;
      LAYER li1 ;
        RECT 775.835 211.770 776.165 212.570 ;
        RECT 776.725 211.770 777.015 212.495 ;
        RECT 777.275 212.420 778.695 212.590 ;
      LAYER li1 ;
        RECT 778.955 212.420 781.645 212.590 ;
      LAYER li1 ;
        RECT 777.275 211.940 777.445 212.420 ;
        RECT 777.615 211.770 777.945 212.250 ;
        RECT 778.115 211.945 778.285 212.420 ;
        RECT 778.455 211.770 778.785 212.250 ;
      LAYER li1 ;
        RECT 778.955 211.940 779.125 212.420 ;
      LAYER li1 ;
        RECT 779.295 211.770 779.625 212.250 ;
      LAYER li1 ;
        RECT 779.795 211.940 779.965 212.420 ;
      LAYER li1 ;
        RECT 780.135 211.770 780.465 212.250 ;
      LAYER li1 ;
        RECT 780.635 211.940 780.805 212.420 ;
      LAYER li1 ;
        RECT 780.975 211.770 781.305 212.250 ;
      LAYER li1 ;
        RECT 781.475 211.940 781.645 212.420 ;
      LAYER li1 ;
        RECT 781.815 211.770 782.145 212.570 ;
        RECT 782.705 211.770 782.995 212.495 ;
        RECT 783.255 212.420 784.675 212.590 ;
      LAYER li1 ;
        RECT 784.935 212.420 787.625 212.590 ;
      LAYER li1 ;
        RECT 792.985 212.590 793.160 212.760 ;
      LAYER li1 ;
        RECT 2149.950 212.635 2150.300 213.885 ;
      LAYER li1 ;
        RECT 2152.065 213.155 2152.355 214.320 ;
        RECT 2152.535 213.300 2152.865 214.150 ;
        RECT 2153.035 213.520 2153.205 214.320 ;
        RECT 2153.375 213.300 2153.705 214.150 ;
        RECT 2153.875 213.520 2154.045 214.320 ;
        RECT 2154.635 213.520 2154.965 214.320 ;
        RECT 2155.475 213.520 2155.805 214.320 ;
        RECT 2156.315 213.520 2156.645 214.320 ;
        RECT 2152.535 213.130 2154.035 213.300 ;
        RECT 2157.155 213.170 2157.485 214.320 ;
        RECT 2158.045 213.155 2158.335 214.320 ;
        RECT 2158.515 213.300 2158.845 214.150 ;
        RECT 2159.015 213.520 2159.185 214.320 ;
        RECT 2159.355 213.300 2159.685 214.150 ;
        RECT 2159.855 213.520 2160.025 214.320 ;
        RECT 2160.615 213.520 2160.945 214.320 ;
        RECT 2161.455 213.520 2161.785 214.320 ;
        RECT 2162.295 213.520 2162.625 214.320 ;
        RECT 2158.515 213.130 2160.015 213.300 ;
        RECT 2163.135 213.170 2163.465 214.320 ;
        RECT 2164.025 213.155 2164.315 214.320 ;
        RECT 2164.495 213.300 2164.825 214.150 ;
        RECT 2164.995 213.520 2165.165 214.320 ;
        RECT 2165.335 213.300 2165.665 214.150 ;
        RECT 2165.835 213.520 2166.005 214.320 ;
        RECT 2166.595 213.520 2166.925 214.320 ;
        RECT 2167.435 213.520 2167.765 214.320 ;
        RECT 2168.275 213.520 2168.605 214.320 ;
        RECT 2164.495 213.130 2165.995 213.300 ;
        RECT 2169.115 213.170 2169.445 214.320 ;
        RECT 2170.005 213.155 2170.295 214.320 ;
        RECT 2170.475 213.300 2170.805 214.150 ;
        RECT 2170.975 213.520 2171.145 214.320 ;
        RECT 2171.315 213.300 2171.645 214.150 ;
        RECT 2171.815 213.520 2171.985 214.320 ;
        RECT 2172.575 213.520 2172.905 214.320 ;
        RECT 2173.415 213.520 2173.745 214.320 ;
        RECT 2174.255 213.520 2174.585 214.320 ;
        RECT 2170.475 213.130 2171.975 213.300 ;
        RECT 2175.095 213.170 2175.425 214.320 ;
        RECT 2175.985 213.155 2176.275 214.320 ;
        RECT 2176.455 213.300 2176.785 214.150 ;
        RECT 2176.955 213.520 2177.125 214.320 ;
        RECT 2177.295 213.300 2177.625 214.150 ;
        RECT 2177.795 213.520 2177.965 214.320 ;
        RECT 2178.555 213.520 2178.885 214.320 ;
        RECT 2179.395 213.520 2179.725 214.320 ;
        RECT 2180.235 213.520 2180.565 214.320 ;
        RECT 2176.455 213.130 2177.955 213.300 ;
        RECT 2181.075 213.170 2181.405 214.320 ;
        RECT 2181.965 213.155 2182.255 214.320 ;
        RECT 2182.435 213.300 2182.765 214.150 ;
        RECT 2182.935 213.520 2183.105 214.320 ;
        RECT 2183.275 213.300 2183.605 214.150 ;
        RECT 2183.775 213.520 2183.945 214.320 ;
        RECT 2184.535 213.520 2184.865 214.320 ;
        RECT 2185.375 213.520 2185.705 214.320 ;
        RECT 2186.215 213.520 2186.545 214.320 ;
        RECT 2182.435 213.130 2183.935 213.300 ;
        RECT 2187.055 213.170 2187.385 214.320 ;
        RECT 2187.945 213.155 2188.235 214.320 ;
        RECT 2188.415 213.300 2188.745 214.150 ;
        RECT 2188.915 213.520 2189.085 214.320 ;
        RECT 2189.255 213.300 2189.585 214.150 ;
        RECT 2189.755 213.520 2189.925 214.320 ;
        RECT 2190.515 213.520 2190.845 214.320 ;
        RECT 2191.355 213.520 2191.685 214.320 ;
        RECT 2192.195 213.520 2192.525 214.320 ;
        RECT 2188.415 213.130 2189.915 213.300 ;
        RECT 2193.035 213.170 2193.365 214.320 ;
        RECT 2193.925 213.155 2194.215 214.320 ;
        RECT 2194.395 213.300 2194.725 214.150 ;
        RECT 2194.895 213.520 2195.065 214.320 ;
        RECT 2195.235 213.300 2195.565 214.150 ;
        RECT 2195.735 213.520 2195.905 214.320 ;
        RECT 2196.495 213.520 2196.825 214.320 ;
        RECT 2197.335 213.520 2197.665 214.320 ;
        RECT 2198.175 213.520 2198.505 214.320 ;
        RECT 2194.395 213.130 2195.895 213.300 ;
        RECT 2199.015 213.170 2199.345 214.320 ;
        RECT 2199.905 213.155 2200.195 214.320 ;
        RECT 2200.375 213.300 2200.705 214.150 ;
        RECT 2200.875 213.520 2201.045 214.320 ;
        RECT 2201.215 213.300 2201.545 214.150 ;
        RECT 2201.715 213.520 2201.885 214.320 ;
        RECT 2202.475 213.520 2202.805 214.320 ;
        RECT 2203.315 213.520 2203.645 214.320 ;
        RECT 2204.155 213.520 2204.485 214.320 ;
        RECT 2200.375 213.130 2201.875 213.300 ;
        RECT 2204.995 213.170 2205.325 214.320 ;
        RECT 2205.885 213.155 2206.175 214.320 ;
        RECT 2206.355 213.300 2206.685 214.150 ;
        RECT 2206.855 213.520 2207.025 214.320 ;
        RECT 2207.195 213.300 2207.525 214.150 ;
        RECT 2207.695 213.520 2207.865 214.320 ;
        RECT 2208.455 213.520 2208.785 214.320 ;
        RECT 2209.295 213.520 2209.625 214.320 ;
        RECT 2210.135 213.520 2210.465 214.320 ;
        RECT 2206.355 213.130 2207.855 213.300 ;
        RECT 2210.975 213.170 2211.305 214.320 ;
        RECT 2211.865 213.155 2212.155 214.320 ;
        RECT 2212.335 213.300 2212.665 214.150 ;
        RECT 2212.835 213.520 2213.005 214.320 ;
        RECT 2213.175 213.300 2213.505 214.150 ;
        RECT 2213.675 213.520 2213.845 214.320 ;
        RECT 2214.435 213.520 2214.765 214.320 ;
        RECT 2215.275 213.520 2215.605 214.320 ;
        RECT 2216.115 213.520 2216.445 214.320 ;
        RECT 2212.335 213.130 2213.835 213.300 ;
        RECT 2216.955 213.170 2217.285 214.320 ;
        RECT 2217.845 213.155 2218.135 214.320 ;
        RECT 2218.315 213.300 2218.645 214.150 ;
        RECT 2218.815 213.520 2218.985 214.320 ;
        RECT 2219.155 213.300 2219.485 214.150 ;
        RECT 2219.655 213.520 2219.825 214.320 ;
        RECT 2220.415 213.520 2220.745 214.320 ;
        RECT 2221.255 213.520 2221.585 214.320 ;
        RECT 2222.095 213.520 2222.425 214.320 ;
        RECT 2218.315 213.130 2219.815 213.300 ;
        RECT 2222.935 213.170 2223.265 214.320 ;
        RECT 2223.825 213.155 2224.115 214.320 ;
        RECT 2224.295 213.300 2224.625 214.150 ;
        RECT 2224.795 213.520 2224.965 214.320 ;
        RECT 2225.135 213.300 2225.465 214.150 ;
        RECT 2225.635 213.520 2225.805 214.320 ;
        RECT 2226.395 213.520 2226.725 214.320 ;
        RECT 2227.235 213.520 2227.565 214.320 ;
        RECT 2228.075 213.520 2228.405 214.320 ;
        RECT 2224.295 213.130 2225.795 213.300 ;
        RECT 2228.915 213.170 2229.245 214.320 ;
        RECT 2229.805 213.155 2230.095 214.320 ;
        RECT 2230.275 213.300 2230.605 214.150 ;
        RECT 2230.775 213.520 2230.945 214.320 ;
        RECT 2231.115 213.300 2231.445 214.150 ;
        RECT 2231.615 213.520 2231.785 214.320 ;
        RECT 2232.375 213.520 2232.705 214.320 ;
        RECT 2233.215 213.520 2233.545 214.320 ;
        RECT 2234.055 213.520 2234.385 214.320 ;
        RECT 2230.275 213.130 2231.775 213.300 ;
        RECT 2234.895 213.170 2235.225 214.320 ;
        RECT 2235.785 213.155 2236.075 214.320 ;
        RECT 2236.255 213.300 2236.585 214.150 ;
        RECT 2236.755 213.520 2236.925 214.320 ;
        RECT 2237.095 213.300 2237.425 214.150 ;
        RECT 2237.595 213.520 2237.765 214.320 ;
        RECT 2238.355 213.520 2238.685 214.320 ;
        RECT 2239.195 213.520 2239.525 214.320 ;
        RECT 2240.035 213.520 2240.365 214.320 ;
        RECT 2236.255 213.130 2237.755 213.300 ;
        RECT 2240.875 213.170 2241.205 214.320 ;
        RECT 2241.765 213.155 2242.055 214.320 ;
        RECT 2242.235 213.300 2242.565 214.150 ;
        RECT 2242.735 213.520 2242.905 214.320 ;
        RECT 2243.075 213.300 2243.405 214.150 ;
        RECT 2243.575 213.520 2243.745 214.320 ;
        RECT 2244.335 213.520 2244.665 214.320 ;
        RECT 2245.175 213.520 2245.505 214.320 ;
        RECT 2246.015 213.520 2246.345 214.320 ;
        RECT 2242.235 213.130 2243.735 213.300 ;
        RECT 2246.855 213.170 2247.185 214.320 ;
        RECT 2247.745 213.155 2248.035 214.320 ;
        RECT 2248.215 213.300 2248.545 214.150 ;
        RECT 2248.715 213.520 2248.885 214.320 ;
        RECT 2249.055 213.300 2249.385 214.150 ;
        RECT 2249.555 213.520 2249.725 214.320 ;
        RECT 2250.315 213.520 2250.645 214.320 ;
        RECT 2251.155 213.520 2251.485 214.320 ;
        RECT 2251.995 213.520 2252.325 214.320 ;
        RECT 2248.215 213.130 2249.715 213.300 ;
        RECT 2252.835 213.170 2253.165 214.320 ;
        RECT 2253.725 213.155 2254.015 214.320 ;
        RECT 2254.195 213.300 2254.525 214.150 ;
        RECT 2254.695 213.520 2254.865 214.320 ;
        RECT 2255.035 213.300 2255.365 214.150 ;
        RECT 2255.535 213.520 2255.705 214.320 ;
        RECT 2256.295 213.520 2256.625 214.320 ;
        RECT 2257.135 213.520 2257.465 214.320 ;
        RECT 2257.975 213.520 2258.305 214.320 ;
        RECT 2254.195 213.130 2255.695 213.300 ;
        RECT 2258.815 213.170 2259.145 214.320 ;
        RECT 2259.705 213.155 2259.995 214.320 ;
        RECT 2260.175 213.300 2260.505 214.150 ;
        RECT 2260.675 213.520 2260.845 214.320 ;
        RECT 2261.015 213.300 2261.345 214.150 ;
        RECT 2261.515 213.520 2261.685 214.320 ;
        RECT 2262.275 213.520 2262.605 214.320 ;
        RECT 2263.115 213.520 2263.445 214.320 ;
        RECT 2263.955 213.520 2264.285 214.320 ;
        RECT 2260.175 213.130 2261.675 213.300 ;
        RECT 2264.795 213.170 2265.125 214.320 ;
        RECT 2265.685 213.155 2265.975 214.320 ;
        RECT 2266.535 213.170 2266.865 214.320 ;
      LAYER li1 ;
        RECT 2267.035 213.300 2267.205 214.150 ;
      LAYER li1 ;
        RECT 2267.375 213.520 2267.705 214.320 ;
      LAYER li1 ;
        RECT 2267.875 213.300 2268.045 214.150 ;
      LAYER li1 ;
        RECT 2268.215 213.520 2268.545 214.320 ;
      LAYER li1 ;
        RECT 2268.715 213.300 2268.885 214.150 ;
      LAYER li1 ;
        RECT 2269.055 213.520 2269.385 214.320 ;
      LAYER li1 ;
        RECT 2269.555 213.300 2269.725 214.150 ;
      LAYER li1 ;
        RECT 2269.975 213.520 2270.145 214.320 ;
        RECT 2270.315 213.300 2270.645 214.150 ;
        RECT 2270.815 213.520 2270.985 214.320 ;
        RECT 2271.155 213.300 2271.485 214.150 ;
      LAYER li1 ;
        RECT 2152.580 212.760 2153.680 212.960 ;
      LAYER li1 ;
        RECT 2153.860 212.930 2154.035 213.130 ;
        RECT 2153.860 212.760 2156.485 212.930 ;
      LAYER li1 ;
        RECT 2158.560 212.760 2159.660 212.960 ;
      LAYER li1 ;
        RECT 2159.840 212.930 2160.015 213.130 ;
        RECT 2159.840 212.760 2162.465 212.930 ;
      LAYER li1 ;
        RECT 2164.540 212.760 2165.640 212.960 ;
      LAYER li1 ;
        RECT 2165.820 212.930 2165.995 213.130 ;
        RECT 2165.820 212.760 2168.445 212.930 ;
      LAYER li1 ;
        RECT 2170.520 212.760 2171.620 212.960 ;
      LAYER li1 ;
        RECT 2171.800 212.930 2171.975 213.130 ;
        RECT 2171.800 212.760 2174.425 212.930 ;
      LAYER li1 ;
        RECT 2176.500 212.760 2177.600 212.960 ;
      LAYER li1 ;
        RECT 2177.780 212.930 2177.955 213.130 ;
        RECT 2177.780 212.760 2180.405 212.930 ;
      LAYER li1 ;
        RECT 2182.480 212.760 2183.580 212.960 ;
      LAYER li1 ;
        RECT 2183.760 212.930 2183.935 213.130 ;
        RECT 2183.760 212.760 2186.385 212.930 ;
      LAYER li1 ;
        RECT 2188.460 212.760 2189.560 212.960 ;
      LAYER li1 ;
        RECT 2189.740 212.930 2189.915 213.130 ;
        RECT 2189.740 212.760 2192.365 212.930 ;
      LAYER li1 ;
        RECT 2194.440 212.760 2195.540 212.960 ;
      LAYER li1 ;
        RECT 2195.720 212.930 2195.895 213.130 ;
        RECT 2195.720 212.760 2198.345 212.930 ;
      LAYER li1 ;
        RECT 2200.420 212.760 2201.520 212.960 ;
      LAYER li1 ;
        RECT 2201.700 212.930 2201.875 213.130 ;
        RECT 2201.700 212.760 2204.325 212.930 ;
      LAYER li1 ;
        RECT 2206.400 212.760 2207.500 212.960 ;
      LAYER li1 ;
        RECT 2207.680 212.930 2207.855 213.130 ;
        RECT 2207.680 212.760 2210.305 212.930 ;
      LAYER li1 ;
        RECT 2212.380 212.760 2213.480 212.960 ;
      LAYER li1 ;
        RECT 2213.660 212.930 2213.835 213.130 ;
        RECT 2213.660 212.760 2216.285 212.930 ;
      LAYER li1 ;
        RECT 2218.360 212.760 2219.460 212.960 ;
      LAYER li1 ;
        RECT 2219.640 212.930 2219.815 213.130 ;
        RECT 2219.640 212.760 2222.265 212.930 ;
      LAYER li1 ;
        RECT 2224.340 212.760 2225.440 212.960 ;
      LAYER li1 ;
        RECT 2225.620 212.930 2225.795 213.130 ;
        RECT 2225.620 212.760 2228.245 212.930 ;
      LAYER li1 ;
        RECT 2230.320 212.760 2231.420 212.960 ;
      LAYER li1 ;
        RECT 2231.600 212.930 2231.775 213.130 ;
        RECT 2231.600 212.760 2234.225 212.930 ;
      LAYER li1 ;
        RECT 2236.300 212.760 2237.400 212.960 ;
      LAYER li1 ;
        RECT 2237.580 212.930 2237.755 213.130 ;
        RECT 2237.580 212.760 2240.205 212.930 ;
      LAYER li1 ;
        RECT 2242.280 212.760 2243.380 212.960 ;
      LAYER li1 ;
        RECT 2243.560 212.930 2243.735 213.130 ;
        RECT 2243.560 212.760 2246.185 212.930 ;
      LAYER li1 ;
        RECT 2248.260 212.760 2249.360 212.960 ;
      LAYER li1 ;
        RECT 2249.540 212.930 2249.715 213.130 ;
        RECT 2249.540 212.760 2252.165 212.930 ;
      LAYER li1 ;
        RECT 2254.240 212.760 2255.340 212.960 ;
      LAYER li1 ;
        RECT 2255.520 212.930 2255.695 213.130 ;
        RECT 2255.520 212.760 2258.145 212.930 ;
      LAYER li1 ;
        RECT 2260.220 212.760 2261.320 212.960 ;
      LAYER li1 ;
        RECT 2261.500 212.930 2261.675 213.130 ;
      LAYER li1 ;
        RECT 2267.035 213.130 2269.725 213.300 ;
      LAYER li1 ;
        RECT 2269.985 213.130 2271.485 213.300 ;
        RECT 2271.665 213.155 2271.955 214.320 ;
        RECT 2261.500 212.760 2264.125 212.930 ;
        RECT 2153.860 212.590 2154.035 212.760 ;
        RECT 2159.840 212.590 2160.015 212.760 ;
        RECT 2165.820 212.590 2165.995 212.760 ;
        RECT 2171.800 212.590 2171.975 212.760 ;
        RECT 2177.780 212.590 2177.955 212.760 ;
        RECT 2183.760 212.590 2183.935 212.760 ;
        RECT 2189.740 212.590 2189.915 212.760 ;
        RECT 2195.720 212.590 2195.895 212.760 ;
        RECT 2201.700 212.590 2201.875 212.760 ;
        RECT 2207.680 212.590 2207.855 212.760 ;
        RECT 2213.660 212.590 2213.835 212.760 ;
        RECT 2219.640 212.590 2219.815 212.760 ;
        RECT 2225.620 212.590 2225.795 212.760 ;
        RECT 2231.600 212.590 2231.775 212.760 ;
        RECT 2237.580 212.590 2237.755 212.760 ;
        RECT 2243.560 212.590 2243.735 212.760 ;
        RECT 2249.540 212.590 2249.715 212.760 ;
        RECT 2255.520 212.590 2255.695 212.760 ;
        RECT 2261.500 212.590 2261.675 212.760 ;
        RECT 783.255 211.940 783.425 212.420 ;
        RECT 783.595 211.770 783.925 212.250 ;
        RECT 784.095 211.945 784.265 212.420 ;
        RECT 784.435 211.770 784.765 212.250 ;
      LAYER li1 ;
        RECT 784.935 211.940 785.105 212.420 ;
      LAYER li1 ;
        RECT 785.275 211.770 785.605 212.250 ;
      LAYER li1 ;
        RECT 785.775 211.940 785.945 212.420 ;
      LAYER li1 ;
        RECT 786.115 211.770 786.445 212.250 ;
      LAYER li1 ;
        RECT 786.615 211.940 786.785 212.420 ;
      LAYER li1 ;
        RECT 786.955 211.770 787.285 212.250 ;
      LAYER li1 ;
        RECT 787.455 211.940 787.625 212.420 ;
      LAYER li1 ;
        RECT 787.795 211.770 788.125 212.570 ;
        RECT 788.685 211.770 788.975 212.495 ;
        RECT 789.535 211.770 789.865 212.570 ;
        RECT 792.985 212.420 794.405 212.590 ;
        RECT 790.375 211.770 790.705 212.250 ;
        RECT 791.215 211.770 791.545 212.250 ;
        RECT 792.055 211.770 792.385 212.250 ;
        RECT 792.895 211.770 793.225 212.250 ;
        RECT 793.395 211.945 793.565 212.420 ;
        RECT 793.735 211.770 794.065 212.250 ;
        RECT 794.235 211.940 794.405 212.420 ;
        RECT 794.665 211.770 794.955 212.495 ;
        RECT 2146.085 211.770 2146.375 212.495 ;
        RECT 2152.065 211.770 2152.355 212.495 ;
        RECT 2152.615 212.420 2154.035 212.590 ;
        RECT 2152.615 211.940 2152.785 212.420 ;
        RECT 2152.955 211.770 2153.285 212.250 ;
        RECT 2153.455 211.945 2153.625 212.420 ;
        RECT 2153.795 211.770 2154.125 212.250 ;
        RECT 2154.635 211.770 2154.965 212.250 ;
        RECT 2155.475 211.770 2155.805 212.250 ;
        RECT 2156.315 211.770 2156.645 212.250 ;
        RECT 2157.155 211.770 2157.485 212.570 ;
        RECT 2158.045 211.770 2158.335 212.495 ;
        RECT 2158.595 212.420 2160.015 212.590 ;
        RECT 2158.595 211.940 2158.765 212.420 ;
        RECT 2158.935 211.770 2159.265 212.250 ;
        RECT 2159.435 211.945 2159.605 212.420 ;
        RECT 2159.775 211.770 2160.105 212.250 ;
        RECT 2160.615 211.770 2160.945 212.250 ;
        RECT 2161.455 211.770 2161.785 212.250 ;
        RECT 2162.295 211.770 2162.625 212.250 ;
        RECT 2163.135 211.770 2163.465 212.570 ;
        RECT 2164.025 211.770 2164.315 212.495 ;
        RECT 2164.575 212.420 2165.995 212.590 ;
        RECT 2164.575 211.940 2164.745 212.420 ;
        RECT 2164.915 211.770 2165.245 212.250 ;
        RECT 2165.415 211.945 2165.585 212.420 ;
        RECT 2165.755 211.770 2166.085 212.250 ;
        RECT 2166.595 211.770 2166.925 212.250 ;
        RECT 2167.435 211.770 2167.765 212.250 ;
        RECT 2168.275 211.770 2168.605 212.250 ;
        RECT 2169.115 211.770 2169.445 212.570 ;
        RECT 2170.005 211.770 2170.295 212.495 ;
        RECT 2170.555 212.420 2171.975 212.590 ;
        RECT 2170.555 211.940 2170.725 212.420 ;
        RECT 2170.895 211.770 2171.225 212.250 ;
        RECT 2171.395 211.945 2171.565 212.420 ;
        RECT 2171.735 211.770 2172.065 212.250 ;
        RECT 2172.575 211.770 2172.905 212.250 ;
        RECT 2173.415 211.770 2173.745 212.250 ;
        RECT 2174.255 211.770 2174.585 212.250 ;
        RECT 2175.095 211.770 2175.425 212.570 ;
        RECT 2175.985 211.770 2176.275 212.495 ;
        RECT 2176.535 212.420 2177.955 212.590 ;
        RECT 2176.535 211.940 2176.705 212.420 ;
        RECT 2176.875 211.770 2177.205 212.250 ;
        RECT 2177.375 211.945 2177.545 212.420 ;
        RECT 2177.715 211.770 2178.045 212.250 ;
        RECT 2178.555 211.770 2178.885 212.250 ;
        RECT 2179.395 211.770 2179.725 212.250 ;
        RECT 2180.235 211.770 2180.565 212.250 ;
        RECT 2181.075 211.770 2181.405 212.570 ;
        RECT 2181.965 211.770 2182.255 212.495 ;
        RECT 2182.515 212.420 2183.935 212.590 ;
        RECT 2182.515 211.940 2182.685 212.420 ;
        RECT 2182.855 211.770 2183.185 212.250 ;
        RECT 2183.355 211.945 2183.525 212.420 ;
        RECT 2183.695 211.770 2184.025 212.250 ;
        RECT 2184.535 211.770 2184.865 212.250 ;
        RECT 2185.375 211.770 2185.705 212.250 ;
        RECT 2186.215 211.770 2186.545 212.250 ;
        RECT 2187.055 211.770 2187.385 212.570 ;
        RECT 2187.945 211.770 2188.235 212.495 ;
        RECT 2188.495 212.420 2189.915 212.590 ;
        RECT 2188.495 211.940 2188.665 212.420 ;
        RECT 2188.835 211.770 2189.165 212.250 ;
        RECT 2189.335 211.945 2189.505 212.420 ;
        RECT 2189.675 211.770 2190.005 212.250 ;
        RECT 2190.515 211.770 2190.845 212.250 ;
        RECT 2191.355 211.770 2191.685 212.250 ;
        RECT 2192.195 211.770 2192.525 212.250 ;
        RECT 2193.035 211.770 2193.365 212.570 ;
        RECT 2193.925 211.770 2194.215 212.495 ;
        RECT 2194.475 212.420 2195.895 212.590 ;
        RECT 2194.475 211.940 2194.645 212.420 ;
        RECT 2194.815 211.770 2195.145 212.250 ;
        RECT 2195.315 211.945 2195.485 212.420 ;
        RECT 2195.655 211.770 2195.985 212.250 ;
        RECT 2196.495 211.770 2196.825 212.250 ;
        RECT 2197.335 211.770 2197.665 212.250 ;
        RECT 2198.175 211.770 2198.505 212.250 ;
        RECT 2199.015 211.770 2199.345 212.570 ;
        RECT 2199.905 211.770 2200.195 212.495 ;
        RECT 2200.455 212.420 2201.875 212.590 ;
        RECT 2200.455 211.940 2200.625 212.420 ;
        RECT 2200.795 211.770 2201.125 212.250 ;
        RECT 2201.295 211.945 2201.465 212.420 ;
        RECT 2201.635 211.770 2201.965 212.250 ;
        RECT 2202.475 211.770 2202.805 212.250 ;
        RECT 2203.315 211.770 2203.645 212.250 ;
        RECT 2204.155 211.770 2204.485 212.250 ;
        RECT 2204.995 211.770 2205.325 212.570 ;
        RECT 2205.885 211.770 2206.175 212.495 ;
        RECT 2206.435 212.420 2207.855 212.590 ;
        RECT 2206.435 211.940 2206.605 212.420 ;
        RECT 2206.775 211.770 2207.105 212.250 ;
        RECT 2207.275 211.945 2207.445 212.420 ;
        RECT 2207.615 211.770 2207.945 212.250 ;
        RECT 2208.455 211.770 2208.785 212.250 ;
        RECT 2209.295 211.770 2209.625 212.250 ;
        RECT 2210.135 211.770 2210.465 212.250 ;
        RECT 2210.975 211.770 2211.305 212.570 ;
        RECT 2211.865 211.770 2212.155 212.495 ;
        RECT 2212.415 212.420 2213.835 212.590 ;
        RECT 2212.415 211.940 2212.585 212.420 ;
        RECT 2212.755 211.770 2213.085 212.250 ;
        RECT 2213.255 211.945 2213.425 212.420 ;
        RECT 2213.595 211.770 2213.925 212.250 ;
        RECT 2214.435 211.770 2214.765 212.250 ;
        RECT 2215.275 211.770 2215.605 212.250 ;
        RECT 2216.115 211.770 2216.445 212.250 ;
        RECT 2216.955 211.770 2217.285 212.570 ;
        RECT 2217.845 211.770 2218.135 212.495 ;
        RECT 2218.395 212.420 2219.815 212.590 ;
        RECT 2218.395 211.940 2218.565 212.420 ;
        RECT 2218.735 211.770 2219.065 212.250 ;
        RECT 2219.235 211.945 2219.405 212.420 ;
        RECT 2219.575 211.770 2219.905 212.250 ;
        RECT 2220.415 211.770 2220.745 212.250 ;
        RECT 2221.255 211.770 2221.585 212.250 ;
        RECT 2222.095 211.770 2222.425 212.250 ;
        RECT 2222.935 211.770 2223.265 212.570 ;
        RECT 2223.825 211.770 2224.115 212.495 ;
        RECT 2224.375 212.420 2225.795 212.590 ;
        RECT 2224.375 211.940 2224.545 212.420 ;
        RECT 2224.715 211.770 2225.045 212.250 ;
        RECT 2225.215 211.945 2225.385 212.420 ;
        RECT 2225.555 211.770 2225.885 212.250 ;
        RECT 2226.395 211.770 2226.725 212.250 ;
        RECT 2227.235 211.770 2227.565 212.250 ;
        RECT 2228.075 211.770 2228.405 212.250 ;
        RECT 2228.915 211.770 2229.245 212.570 ;
        RECT 2229.805 211.770 2230.095 212.495 ;
        RECT 2230.355 212.420 2231.775 212.590 ;
        RECT 2230.355 211.940 2230.525 212.420 ;
        RECT 2230.695 211.770 2231.025 212.250 ;
        RECT 2231.195 211.945 2231.365 212.420 ;
        RECT 2231.535 211.770 2231.865 212.250 ;
        RECT 2232.375 211.770 2232.705 212.250 ;
        RECT 2233.215 211.770 2233.545 212.250 ;
        RECT 2234.055 211.770 2234.385 212.250 ;
        RECT 2234.895 211.770 2235.225 212.570 ;
        RECT 2235.785 211.770 2236.075 212.495 ;
        RECT 2236.335 212.420 2237.755 212.590 ;
        RECT 2236.335 211.940 2236.505 212.420 ;
        RECT 2236.675 211.770 2237.005 212.250 ;
        RECT 2237.175 211.945 2237.345 212.420 ;
        RECT 2237.515 211.770 2237.845 212.250 ;
        RECT 2238.355 211.770 2238.685 212.250 ;
        RECT 2239.195 211.770 2239.525 212.250 ;
        RECT 2240.035 211.770 2240.365 212.250 ;
        RECT 2240.875 211.770 2241.205 212.570 ;
        RECT 2241.765 211.770 2242.055 212.495 ;
        RECT 2242.315 212.420 2243.735 212.590 ;
        RECT 2242.315 211.940 2242.485 212.420 ;
        RECT 2242.655 211.770 2242.985 212.250 ;
        RECT 2243.155 211.945 2243.325 212.420 ;
        RECT 2243.495 211.770 2243.825 212.250 ;
        RECT 2244.335 211.770 2244.665 212.250 ;
        RECT 2245.175 211.770 2245.505 212.250 ;
        RECT 2246.015 211.770 2246.345 212.250 ;
        RECT 2246.855 211.770 2247.185 212.570 ;
        RECT 2247.745 211.770 2248.035 212.495 ;
        RECT 2248.295 212.420 2249.715 212.590 ;
        RECT 2248.295 211.940 2248.465 212.420 ;
        RECT 2248.635 211.770 2248.965 212.250 ;
        RECT 2249.135 211.945 2249.305 212.420 ;
        RECT 2249.475 211.770 2249.805 212.250 ;
        RECT 2250.315 211.770 2250.645 212.250 ;
        RECT 2251.155 211.770 2251.485 212.250 ;
        RECT 2251.995 211.770 2252.325 212.250 ;
        RECT 2252.835 211.770 2253.165 212.570 ;
        RECT 2253.725 211.770 2254.015 212.495 ;
        RECT 2254.275 212.420 2255.695 212.590 ;
        RECT 2254.275 211.940 2254.445 212.420 ;
        RECT 2254.615 211.770 2254.945 212.250 ;
        RECT 2255.115 211.945 2255.285 212.420 ;
        RECT 2255.455 211.770 2255.785 212.250 ;
        RECT 2256.295 211.770 2256.625 212.250 ;
        RECT 2257.135 211.770 2257.465 212.250 ;
        RECT 2257.975 211.770 2258.305 212.250 ;
        RECT 2258.815 211.770 2259.145 212.570 ;
        RECT 2259.705 211.770 2259.995 212.495 ;
        RECT 2260.255 212.420 2261.675 212.590 ;
      LAYER li1 ;
        RECT 2267.035 212.590 2267.290 213.130 ;
      LAYER li1 ;
        RECT 2269.985 212.930 2270.160 213.130 ;
        RECT 2267.535 212.760 2270.160 212.930 ;
        RECT 2269.985 212.590 2270.160 212.760 ;
        RECT 2260.255 211.940 2260.425 212.420 ;
        RECT 2260.595 211.770 2260.925 212.250 ;
        RECT 2261.095 211.945 2261.265 212.420 ;
        RECT 2261.435 211.770 2261.765 212.250 ;
        RECT 2262.275 211.770 2262.605 212.250 ;
        RECT 2263.115 211.770 2263.445 212.250 ;
        RECT 2263.955 211.770 2264.285 212.250 ;
        RECT 2264.795 211.770 2265.125 212.570 ;
        RECT 2265.685 211.770 2265.975 212.495 ;
        RECT 2266.535 211.770 2266.865 212.570 ;
      LAYER li1 ;
        RECT 2267.035 212.420 2269.725 212.590 ;
      LAYER li1 ;
        RECT 2269.985 212.420 2271.405 212.590 ;
      LAYER li1 ;
        RECT 2267.035 211.940 2267.205 212.420 ;
      LAYER li1 ;
        RECT 2267.375 211.770 2267.705 212.250 ;
      LAYER li1 ;
        RECT 2267.875 211.940 2268.045 212.420 ;
      LAYER li1 ;
        RECT 2268.215 211.770 2268.545 212.250 ;
      LAYER li1 ;
        RECT 2268.715 211.940 2268.885 212.420 ;
      LAYER li1 ;
        RECT 2269.055 211.770 2269.385 212.250 ;
      LAYER li1 ;
        RECT 2269.555 211.940 2269.725 212.420 ;
      LAYER li1 ;
        RECT 2269.895 211.770 2270.225 212.250 ;
        RECT 2270.395 211.945 2270.565 212.420 ;
        RECT 2270.735 211.770 2271.065 212.250 ;
        RECT 2271.235 211.940 2271.405 212.420 ;
        RECT 2271.665 211.770 2271.955 212.495 ;
        RECT 669.000 211.600 669.145 211.770 ;
        RECT 669.315 211.600 669.460 211.770 ;
        RECT 674.980 211.600 675.125 211.770 ;
        RECT 675.295 211.600 675.585 211.770 ;
        RECT 675.755 211.600 676.045 211.770 ;
        RECT 676.215 211.600 676.505 211.770 ;
        RECT 676.675 211.600 676.965 211.770 ;
        RECT 677.135 211.600 677.425 211.770 ;
        RECT 677.595 211.600 677.885 211.770 ;
        RECT 678.055 211.600 678.345 211.770 ;
        RECT 678.515 211.600 678.805 211.770 ;
        RECT 678.975 211.600 679.265 211.770 ;
        RECT 679.435 211.600 679.725 211.770 ;
        RECT 679.895 211.600 680.185 211.770 ;
        RECT 680.355 211.600 680.645 211.770 ;
        RECT 680.815 211.600 681.105 211.770 ;
        RECT 681.275 211.600 681.565 211.770 ;
        RECT 681.735 211.600 682.025 211.770 ;
        RECT 682.195 211.600 682.485 211.770 ;
        RECT 682.655 211.600 682.945 211.770 ;
        RECT 683.115 211.600 683.405 211.770 ;
        RECT 683.575 211.600 683.865 211.770 ;
        RECT 684.035 211.600 684.325 211.770 ;
        RECT 684.495 211.600 684.785 211.770 ;
        RECT 684.955 211.600 685.245 211.770 ;
        RECT 685.415 211.600 685.705 211.770 ;
        RECT 685.875 211.600 686.165 211.770 ;
        RECT 686.335 211.600 686.625 211.770 ;
        RECT 686.795 211.600 687.085 211.770 ;
        RECT 687.255 211.600 687.545 211.770 ;
        RECT 687.715 211.600 688.005 211.770 ;
        RECT 688.175 211.600 688.465 211.770 ;
        RECT 688.635 211.600 688.925 211.770 ;
        RECT 689.095 211.600 689.385 211.770 ;
        RECT 689.555 211.600 689.845 211.770 ;
        RECT 690.015 211.600 690.305 211.770 ;
        RECT 690.475 211.600 690.765 211.770 ;
        RECT 690.935 211.600 691.225 211.770 ;
        RECT 691.395 211.600 691.685 211.770 ;
        RECT 691.855 211.600 692.145 211.770 ;
        RECT 692.315 211.600 692.605 211.770 ;
        RECT 692.775 211.600 693.065 211.770 ;
        RECT 693.235 211.600 693.525 211.770 ;
        RECT 693.695 211.600 693.985 211.770 ;
        RECT 694.155 211.600 694.445 211.770 ;
        RECT 694.615 211.600 694.905 211.770 ;
        RECT 695.075 211.600 695.365 211.770 ;
        RECT 695.535 211.600 695.825 211.770 ;
        RECT 695.995 211.600 696.285 211.770 ;
        RECT 696.455 211.600 696.745 211.770 ;
        RECT 696.915 211.600 697.205 211.770 ;
        RECT 697.375 211.600 697.665 211.770 ;
        RECT 697.835 211.600 698.125 211.770 ;
        RECT 698.295 211.600 698.585 211.770 ;
        RECT 698.755 211.600 699.045 211.770 ;
        RECT 699.215 211.600 699.505 211.770 ;
        RECT 699.675 211.600 699.965 211.770 ;
        RECT 700.135 211.600 700.425 211.770 ;
        RECT 700.595 211.600 700.885 211.770 ;
        RECT 701.055 211.600 701.345 211.770 ;
        RECT 701.515 211.600 701.805 211.770 ;
        RECT 701.975 211.600 702.265 211.770 ;
        RECT 702.435 211.600 702.725 211.770 ;
        RECT 702.895 211.600 703.185 211.770 ;
        RECT 703.355 211.600 703.645 211.770 ;
        RECT 703.815 211.600 704.105 211.770 ;
        RECT 704.275 211.600 704.565 211.770 ;
        RECT 704.735 211.600 705.025 211.770 ;
        RECT 705.195 211.600 705.485 211.770 ;
        RECT 705.655 211.600 705.945 211.770 ;
        RECT 706.115 211.600 706.405 211.770 ;
        RECT 706.575 211.600 706.865 211.770 ;
        RECT 707.035 211.600 707.325 211.770 ;
        RECT 707.495 211.600 707.785 211.770 ;
        RECT 707.955 211.600 708.245 211.770 ;
        RECT 708.415 211.600 708.705 211.770 ;
        RECT 708.875 211.600 709.165 211.770 ;
        RECT 709.335 211.600 709.625 211.770 ;
        RECT 709.795 211.600 710.085 211.770 ;
        RECT 710.255 211.600 710.545 211.770 ;
        RECT 710.715 211.600 711.005 211.770 ;
        RECT 711.175 211.600 711.465 211.770 ;
        RECT 711.635 211.600 711.925 211.770 ;
        RECT 712.095 211.600 712.385 211.770 ;
        RECT 712.555 211.600 712.845 211.770 ;
        RECT 713.015 211.600 713.305 211.770 ;
        RECT 713.475 211.600 713.765 211.770 ;
        RECT 713.935 211.600 714.225 211.770 ;
        RECT 714.395 211.600 714.685 211.770 ;
        RECT 714.855 211.600 715.145 211.770 ;
        RECT 715.315 211.600 715.605 211.770 ;
        RECT 715.775 211.600 716.065 211.770 ;
        RECT 716.235 211.600 716.525 211.770 ;
        RECT 716.695 211.600 716.985 211.770 ;
        RECT 717.155 211.600 717.445 211.770 ;
        RECT 717.615 211.600 717.905 211.770 ;
        RECT 718.075 211.600 718.365 211.770 ;
        RECT 718.535 211.600 718.825 211.770 ;
        RECT 718.995 211.600 719.285 211.770 ;
        RECT 719.455 211.600 719.745 211.770 ;
        RECT 719.915 211.600 720.205 211.770 ;
        RECT 720.375 211.600 720.665 211.770 ;
        RECT 720.835 211.600 721.125 211.770 ;
        RECT 721.295 211.600 721.585 211.770 ;
        RECT 721.755 211.600 722.045 211.770 ;
        RECT 722.215 211.600 722.505 211.770 ;
        RECT 722.675 211.600 722.965 211.770 ;
        RECT 723.135 211.600 723.425 211.770 ;
        RECT 723.595 211.600 723.885 211.770 ;
        RECT 724.055 211.600 724.345 211.770 ;
        RECT 724.515 211.600 724.805 211.770 ;
        RECT 724.975 211.600 725.265 211.770 ;
        RECT 725.435 211.600 725.725 211.770 ;
        RECT 725.895 211.600 726.185 211.770 ;
        RECT 726.355 211.600 726.645 211.770 ;
        RECT 726.815 211.600 727.105 211.770 ;
        RECT 727.275 211.600 727.565 211.770 ;
        RECT 727.735 211.600 728.025 211.770 ;
        RECT 728.195 211.600 728.485 211.770 ;
        RECT 728.655 211.600 728.945 211.770 ;
        RECT 729.115 211.600 729.405 211.770 ;
        RECT 729.575 211.600 729.865 211.770 ;
        RECT 730.035 211.600 730.325 211.770 ;
        RECT 730.495 211.600 730.785 211.770 ;
        RECT 730.955 211.600 731.245 211.770 ;
        RECT 731.415 211.600 731.705 211.770 ;
        RECT 731.875 211.600 732.165 211.770 ;
        RECT 732.335 211.600 732.625 211.770 ;
        RECT 732.795 211.600 733.085 211.770 ;
        RECT 733.255 211.600 733.545 211.770 ;
        RECT 733.715 211.600 734.005 211.770 ;
        RECT 734.175 211.600 734.465 211.770 ;
        RECT 734.635 211.600 734.925 211.770 ;
        RECT 735.095 211.600 735.385 211.770 ;
        RECT 735.555 211.600 735.845 211.770 ;
        RECT 736.015 211.600 736.305 211.770 ;
        RECT 736.475 211.600 736.765 211.770 ;
        RECT 736.935 211.600 737.225 211.770 ;
        RECT 737.395 211.600 737.685 211.770 ;
        RECT 737.855 211.600 738.145 211.770 ;
        RECT 738.315 211.600 738.605 211.770 ;
        RECT 738.775 211.600 739.065 211.770 ;
        RECT 739.235 211.600 739.525 211.770 ;
        RECT 739.695 211.600 739.985 211.770 ;
        RECT 740.155 211.600 740.445 211.770 ;
        RECT 740.615 211.600 740.905 211.770 ;
        RECT 741.075 211.600 741.365 211.770 ;
        RECT 741.535 211.600 741.825 211.770 ;
        RECT 741.995 211.600 742.285 211.770 ;
        RECT 742.455 211.600 742.745 211.770 ;
        RECT 742.915 211.600 743.205 211.770 ;
        RECT 743.375 211.600 743.665 211.770 ;
        RECT 743.835 211.600 744.125 211.770 ;
        RECT 744.295 211.600 744.585 211.770 ;
        RECT 744.755 211.600 745.045 211.770 ;
        RECT 745.215 211.600 745.505 211.770 ;
        RECT 745.675 211.600 745.965 211.770 ;
        RECT 746.135 211.600 746.425 211.770 ;
        RECT 746.595 211.600 746.885 211.770 ;
        RECT 747.055 211.600 747.345 211.770 ;
        RECT 747.515 211.600 747.805 211.770 ;
        RECT 747.975 211.600 748.265 211.770 ;
        RECT 748.435 211.600 748.725 211.770 ;
        RECT 748.895 211.600 749.185 211.770 ;
        RECT 749.355 211.600 749.645 211.770 ;
        RECT 749.815 211.600 750.105 211.770 ;
        RECT 750.275 211.600 750.565 211.770 ;
        RECT 750.735 211.600 751.025 211.770 ;
        RECT 751.195 211.600 751.485 211.770 ;
        RECT 751.655 211.600 751.945 211.770 ;
        RECT 752.115 211.600 752.405 211.770 ;
        RECT 752.575 211.600 752.865 211.770 ;
        RECT 753.035 211.600 753.325 211.770 ;
        RECT 753.495 211.600 753.785 211.770 ;
        RECT 753.955 211.600 754.245 211.770 ;
        RECT 754.415 211.600 754.705 211.770 ;
        RECT 754.875 211.600 755.165 211.770 ;
        RECT 755.335 211.600 755.625 211.770 ;
        RECT 755.795 211.600 756.085 211.770 ;
        RECT 756.255 211.600 756.545 211.770 ;
        RECT 756.715 211.600 757.005 211.770 ;
        RECT 757.175 211.600 757.465 211.770 ;
        RECT 757.635 211.600 757.925 211.770 ;
        RECT 758.095 211.600 758.385 211.770 ;
        RECT 758.555 211.600 758.845 211.770 ;
        RECT 759.015 211.600 759.305 211.770 ;
        RECT 759.475 211.600 759.765 211.770 ;
        RECT 759.935 211.600 760.225 211.770 ;
        RECT 760.395 211.600 760.685 211.770 ;
        RECT 760.855 211.600 761.145 211.770 ;
        RECT 761.315 211.600 761.605 211.770 ;
        RECT 761.775 211.600 762.065 211.770 ;
        RECT 762.235 211.600 762.525 211.770 ;
        RECT 762.695 211.600 762.985 211.770 ;
        RECT 763.155 211.600 763.445 211.770 ;
        RECT 763.615 211.600 763.905 211.770 ;
        RECT 764.075 211.600 764.365 211.770 ;
        RECT 764.535 211.600 764.825 211.770 ;
        RECT 764.995 211.600 765.285 211.770 ;
        RECT 765.455 211.600 765.745 211.770 ;
        RECT 765.915 211.600 766.205 211.770 ;
        RECT 766.375 211.600 766.665 211.770 ;
        RECT 766.835 211.600 767.125 211.770 ;
        RECT 767.295 211.600 767.585 211.770 ;
        RECT 767.755 211.600 768.045 211.770 ;
        RECT 768.215 211.600 768.505 211.770 ;
        RECT 768.675 211.600 768.965 211.770 ;
        RECT 769.135 211.600 769.425 211.770 ;
        RECT 769.595 211.600 769.885 211.770 ;
        RECT 770.055 211.600 770.345 211.770 ;
        RECT 770.515 211.600 770.805 211.770 ;
        RECT 770.975 211.600 771.265 211.770 ;
        RECT 771.435 211.600 771.725 211.770 ;
        RECT 771.895 211.600 772.185 211.770 ;
        RECT 772.355 211.600 772.645 211.770 ;
        RECT 772.815 211.600 773.105 211.770 ;
        RECT 773.275 211.600 773.565 211.770 ;
        RECT 773.735 211.600 774.025 211.770 ;
        RECT 774.195 211.600 774.485 211.770 ;
        RECT 774.655 211.600 774.945 211.770 ;
        RECT 775.115 211.600 775.405 211.770 ;
        RECT 775.575 211.600 775.865 211.770 ;
        RECT 776.035 211.600 776.325 211.770 ;
        RECT 776.495 211.600 776.785 211.770 ;
        RECT 776.955 211.600 777.245 211.770 ;
        RECT 777.415 211.600 777.705 211.770 ;
        RECT 777.875 211.600 778.165 211.770 ;
        RECT 778.335 211.600 778.625 211.770 ;
        RECT 778.795 211.600 779.085 211.770 ;
        RECT 779.255 211.600 779.545 211.770 ;
        RECT 779.715 211.600 780.005 211.770 ;
        RECT 780.175 211.600 780.465 211.770 ;
        RECT 780.635 211.600 780.925 211.770 ;
        RECT 781.095 211.600 781.385 211.770 ;
        RECT 781.555 211.600 781.845 211.770 ;
        RECT 782.015 211.600 782.305 211.770 ;
        RECT 782.475 211.600 782.765 211.770 ;
        RECT 782.935 211.600 783.225 211.770 ;
        RECT 783.395 211.600 783.685 211.770 ;
        RECT 783.855 211.600 784.145 211.770 ;
        RECT 784.315 211.600 784.605 211.770 ;
        RECT 784.775 211.600 785.065 211.770 ;
        RECT 785.235 211.600 785.525 211.770 ;
        RECT 785.695 211.600 785.985 211.770 ;
        RECT 786.155 211.600 786.445 211.770 ;
        RECT 786.615 211.600 786.905 211.770 ;
        RECT 787.075 211.600 787.365 211.770 ;
        RECT 787.535 211.600 787.825 211.770 ;
        RECT 787.995 211.600 788.285 211.770 ;
        RECT 788.455 211.600 788.745 211.770 ;
        RECT 788.915 211.600 789.205 211.770 ;
        RECT 789.375 211.600 789.665 211.770 ;
        RECT 789.835 211.600 790.125 211.770 ;
        RECT 790.295 211.600 790.585 211.770 ;
        RECT 790.755 211.600 791.045 211.770 ;
        RECT 791.215 211.600 791.505 211.770 ;
        RECT 791.675 211.600 791.965 211.770 ;
        RECT 792.135 211.600 792.425 211.770 ;
        RECT 792.595 211.600 792.885 211.770 ;
        RECT 793.055 211.600 793.345 211.770 ;
        RECT 793.515 211.600 793.805 211.770 ;
        RECT 793.975 211.600 794.265 211.770 ;
        RECT 794.435 211.600 794.725 211.770 ;
        RECT 794.895 211.600 795.040 211.770 ;
        RECT 2146.000 211.600 2146.145 211.770 ;
        RECT 2146.315 211.600 2146.460 211.770 ;
        RECT 2151.980 211.600 2152.125 211.770 ;
        RECT 2152.295 211.600 2152.585 211.770 ;
        RECT 2152.755 211.600 2153.045 211.770 ;
        RECT 2153.215 211.600 2153.505 211.770 ;
        RECT 2153.675 211.600 2153.965 211.770 ;
        RECT 2154.135 211.600 2154.425 211.770 ;
        RECT 2154.595 211.600 2154.885 211.770 ;
        RECT 2155.055 211.600 2155.345 211.770 ;
        RECT 2155.515 211.600 2155.805 211.770 ;
        RECT 2155.975 211.600 2156.265 211.770 ;
        RECT 2156.435 211.600 2156.725 211.770 ;
        RECT 2156.895 211.600 2157.185 211.770 ;
        RECT 2157.355 211.600 2157.645 211.770 ;
        RECT 2157.815 211.600 2158.105 211.770 ;
        RECT 2158.275 211.600 2158.565 211.770 ;
        RECT 2158.735 211.600 2159.025 211.770 ;
        RECT 2159.195 211.600 2159.485 211.770 ;
        RECT 2159.655 211.600 2159.945 211.770 ;
        RECT 2160.115 211.600 2160.405 211.770 ;
        RECT 2160.575 211.600 2160.865 211.770 ;
        RECT 2161.035 211.600 2161.325 211.770 ;
        RECT 2161.495 211.600 2161.785 211.770 ;
        RECT 2161.955 211.600 2162.245 211.770 ;
        RECT 2162.415 211.600 2162.705 211.770 ;
        RECT 2162.875 211.600 2163.165 211.770 ;
        RECT 2163.335 211.600 2163.625 211.770 ;
        RECT 2163.795 211.600 2164.085 211.770 ;
        RECT 2164.255 211.600 2164.545 211.770 ;
        RECT 2164.715 211.600 2165.005 211.770 ;
        RECT 2165.175 211.600 2165.465 211.770 ;
        RECT 2165.635 211.600 2165.925 211.770 ;
        RECT 2166.095 211.600 2166.385 211.770 ;
        RECT 2166.555 211.600 2166.845 211.770 ;
        RECT 2167.015 211.600 2167.305 211.770 ;
        RECT 2167.475 211.600 2167.765 211.770 ;
        RECT 2167.935 211.600 2168.225 211.770 ;
        RECT 2168.395 211.600 2168.685 211.770 ;
        RECT 2168.855 211.600 2169.145 211.770 ;
        RECT 2169.315 211.600 2169.605 211.770 ;
        RECT 2169.775 211.600 2170.065 211.770 ;
        RECT 2170.235 211.600 2170.525 211.770 ;
        RECT 2170.695 211.600 2170.985 211.770 ;
        RECT 2171.155 211.600 2171.445 211.770 ;
        RECT 2171.615 211.600 2171.905 211.770 ;
        RECT 2172.075 211.600 2172.365 211.770 ;
        RECT 2172.535 211.600 2172.825 211.770 ;
        RECT 2172.995 211.600 2173.285 211.770 ;
        RECT 2173.455 211.600 2173.745 211.770 ;
        RECT 2173.915 211.600 2174.205 211.770 ;
        RECT 2174.375 211.600 2174.665 211.770 ;
        RECT 2174.835 211.600 2175.125 211.770 ;
        RECT 2175.295 211.600 2175.585 211.770 ;
        RECT 2175.755 211.600 2176.045 211.770 ;
        RECT 2176.215 211.600 2176.505 211.770 ;
        RECT 2176.675 211.600 2176.965 211.770 ;
        RECT 2177.135 211.600 2177.425 211.770 ;
        RECT 2177.595 211.600 2177.885 211.770 ;
        RECT 2178.055 211.600 2178.345 211.770 ;
        RECT 2178.515 211.600 2178.805 211.770 ;
        RECT 2178.975 211.600 2179.265 211.770 ;
        RECT 2179.435 211.600 2179.725 211.770 ;
        RECT 2179.895 211.600 2180.185 211.770 ;
        RECT 2180.355 211.600 2180.645 211.770 ;
        RECT 2180.815 211.600 2181.105 211.770 ;
        RECT 2181.275 211.600 2181.565 211.770 ;
        RECT 2181.735 211.600 2182.025 211.770 ;
        RECT 2182.195 211.600 2182.485 211.770 ;
        RECT 2182.655 211.600 2182.945 211.770 ;
        RECT 2183.115 211.600 2183.405 211.770 ;
        RECT 2183.575 211.600 2183.865 211.770 ;
        RECT 2184.035 211.600 2184.325 211.770 ;
        RECT 2184.495 211.600 2184.785 211.770 ;
        RECT 2184.955 211.600 2185.245 211.770 ;
        RECT 2185.415 211.600 2185.705 211.770 ;
        RECT 2185.875 211.600 2186.165 211.770 ;
        RECT 2186.335 211.600 2186.625 211.770 ;
        RECT 2186.795 211.600 2187.085 211.770 ;
        RECT 2187.255 211.600 2187.545 211.770 ;
        RECT 2187.715 211.600 2188.005 211.770 ;
        RECT 2188.175 211.600 2188.465 211.770 ;
        RECT 2188.635 211.600 2188.925 211.770 ;
        RECT 2189.095 211.600 2189.385 211.770 ;
        RECT 2189.555 211.600 2189.845 211.770 ;
        RECT 2190.015 211.600 2190.305 211.770 ;
        RECT 2190.475 211.600 2190.765 211.770 ;
        RECT 2190.935 211.600 2191.225 211.770 ;
        RECT 2191.395 211.600 2191.685 211.770 ;
        RECT 2191.855 211.600 2192.145 211.770 ;
        RECT 2192.315 211.600 2192.605 211.770 ;
        RECT 2192.775 211.600 2193.065 211.770 ;
        RECT 2193.235 211.600 2193.525 211.770 ;
        RECT 2193.695 211.600 2193.985 211.770 ;
        RECT 2194.155 211.600 2194.445 211.770 ;
        RECT 2194.615 211.600 2194.905 211.770 ;
        RECT 2195.075 211.600 2195.365 211.770 ;
        RECT 2195.535 211.600 2195.825 211.770 ;
        RECT 2195.995 211.600 2196.285 211.770 ;
        RECT 2196.455 211.600 2196.745 211.770 ;
        RECT 2196.915 211.600 2197.205 211.770 ;
        RECT 2197.375 211.600 2197.665 211.770 ;
        RECT 2197.835 211.600 2198.125 211.770 ;
        RECT 2198.295 211.600 2198.585 211.770 ;
        RECT 2198.755 211.600 2199.045 211.770 ;
        RECT 2199.215 211.600 2199.505 211.770 ;
        RECT 2199.675 211.600 2199.965 211.770 ;
        RECT 2200.135 211.600 2200.425 211.770 ;
        RECT 2200.595 211.600 2200.885 211.770 ;
        RECT 2201.055 211.600 2201.345 211.770 ;
        RECT 2201.515 211.600 2201.805 211.770 ;
        RECT 2201.975 211.600 2202.265 211.770 ;
        RECT 2202.435 211.600 2202.725 211.770 ;
        RECT 2202.895 211.600 2203.185 211.770 ;
        RECT 2203.355 211.600 2203.645 211.770 ;
        RECT 2203.815 211.600 2204.105 211.770 ;
        RECT 2204.275 211.600 2204.565 211.770 ;
        RECT 2204.735 211.600 2205.025 211.770 ;
        RECT 2205.195 211.600 2205.485 211.770 ;
        RECT 2205.655 211.600 2205.945 211.770 ;
        RECT 2206.115 211.600 2206.405 211.770 ;
        RECT 2206.575 211.600 2206.865 211.770 ;
        RECT 2207.035 211.600 2207.325 211.770 ;
        RECT 2207.495 211.600 2207.785 211.770 ;
        RECT 2207.955 211.600 2208.245 211.770 ;
        RECT 2208.415 211.600 2208.705 211.770 ;
        RECT 2208.875 211.600 2209.165 211.770 ;
        RECT 2209.335 211.600 2209.625 211.770 ;
        RECT 2209.795 211.600 2210.085 211.770 ;
        RECT 2210.255 211.600 2210.545 211.770 ;
        RECT 2210.715 211.600 2211.005 211.770 ;
        RECT 2211.175 211.600 2211.465 211.770 ;
        RECT 2211.635 211.600 2211.925 211.770 ;
        RECT 2212.095 211.600 2212.385 211.770 ;
        RECT 2212.555 211.600 2212.845 211.770 ;
        RECT 2213.015 211.600 2213.305 211.770 ;
        RECT 2213.475 211.600 2213.765 211.770 ;
        RECT 2213.935 211.600 2214.225 211.770 ;
        RECT 2214.395 211.600 2214.685 211.770 ;
        RECT 2214.855 211.600 2215.145 211.770 ;
        RECT 2215.315 211.600 2215.605 211.770 ;
        RECT 2215.775 211.600 2216.065 211.770 ;
        RECT 2216.235 211.600 2216.525 211.770 ;
        RECT 2216.695 211.600 2216.985 211.770 ;
        RECT 2217.155 211.600 2217.445 211.770 ;
        RECT 2217.615 211.600 2217.905 211.770 ;
        RECT 2218.075 211.600 2218.365 211.770 ;
        RECT 2218.535 211.600 2218.825 211.770 ;
        RECT 2218.995 211.600 2219.285 211.770 ;
        RECT 2219.455 211.600 2219.745 211.770 ;
        RECT 2219.915 211.600 2220.205 211.770 ;
        RECT 2220.375 211.600 2220.665 211.770 ;
        RECT 2220.835 211.600 2221.125 211.770 ;
        RECT 2221.295 211.600 2221.585 211.770 ;
        RECT 2221.755 211.600 2222.045 211.770 ;
        RECT 2222.215 211.600 2222.505 211.770 ;
        RECT 2222.675 211.600 2222.965 211.770 ;
        RECT 2223.135 211.600 2223.425 211.770 ;
        RECT 2223.595 211.600 2223.885 211.770 ;
        RECT 2224.055 211.600 2224.345 211.770 ;
        RECT 2224.515 211.600 2224.805 211.770 ;
        RECT 2224.975 211.600 2225.265 211.770 ;
        RECT 2225.435 211.600 2225.725 211.770 ;
        RECT 2225.895 211.600 2226.185 211.770 ;
        RECT 2226.355 211.600 2226.645 211.770 ;
        RECT 2226.815 211.600 2227.105 211.770 ;
        RECT 2227.275 211.600 2227.565 211.770 ;
        RECT 2227.735 211.600 2228.025 211.770 ;
        RECT 2228.195 211.600 2228.485 211.770 ;
        RECT 2228.655 211.600 2228.945 211.770 ;
        RECT 2229.115 211.600 2229.405 211.770 ;
        RECT 2229.575 211.600 2229.865 211.770 ;
        RECT 2230.035 211.600 2230.325 211.770 ;
        RECT 2230.495 211.600 2230.785 211.770 ;
        RECT 2230.955 211.600 2231.245 211.770 ;
        RECT 2231.415 211.600 2231.705 211.770 ;
        RECT 2231.875 211.600 2232.165 211.770 ;
        RECT 2232.335 211.600 2232.625 211.770 ;
        RECT 2232.795 211.600 2233.085 211.770 ;
        RECT 2233.255 211.600 2233.545 211.770 ;
        RECT 2233.715 211.600 2234.005 211.770 ;
        RECT 2234.175 211.600 2234.465 211.770 ;
        RECT 2234.635 211.600 2234.925 211.770 ;
        RECT 2235.095 211.600 2235.385 211.770 ;
        RECT 2235.555 211.600 2235.845 211.770 ;
        RECT 2236.015 211.600 2236.305 211.770 ;
        RECT 2236.475 211.600 2236.765 211.770 ;
        RECT 2236.935 211.600 2237.225 211.770 ;
        RECT 2237.395 211.600 2237.685 211.770 ;
        RECT 2237.855 211.600 2238.145 211.770 ;
        RECT 2238.315 211.600 2238.605 211.770 ;
        RECT 2238.775 211.600 2239.065 211.770 ;
        RECT 2239.235 211.600 2239.525 211.770 ;
        RECT 2239.695 211.600 2239.985 211.770 ;
        RECT 2240.155 211.600 2240.445 211.770 ;
        RECT 2240.615 211.600 2240.905 211.770 ;
        RECT 2241.075 211.600 2241.365 211.770 ;
        RECT 2241.535 211.600 2241.825 211.770 ;
        RECT 2241.995 211.600 2242.285 211.770 ;
        RECT 2242.455 211.600 2242.745 211.770 ;
        RECT 2242.915 211.600 2243.205 211.770 ;
        RECT 2243.375 211.600 2243.665 211.770 ;
        RECT 2243.835 211.600 2244.125 211.770 ;
        RECT 2244.295 211.600 2244.585 211.770 ;
        RECT 2244.755 211.600 2245.045 211.770 ;
        RECT 2245.215 211.600 2245.505 211.770 ;
        RECT 2245.675 211.600 2245.965 211.770 ;
        RECT 2246.135 211.600 2246.425 211.770 ;
        RECT 2246.595 211.600 2246.885 211.770 ;
        RECT 2247.055 211.600 2247.345 211.770 ;
        RECT 2247.515 211.600 2247.805 211.770 ;
        RECT 2247.975 211.600 2248.265 211.770 ;
        RECT 2248.435 211.600 2248.725 211.770 ;
        RECT 2248.895 211.600 2249.185 211.770 ;
        RECT 2249.355 211.600 2249.645 211.770 ;
        RECT 2249.815 211.600 2250.105 211.770 ;
        RECT 2250.275 211.600 2250.565 211.770 ;
        RECT 2250.735 211.600 2251.025 211.770 ;
        RECT 2251.195 211.600 2251.485 211.770 ;
        RECT 2251.655 211.600 2251.945 211.770 ;
        RECT 2252.115 211.600 2252.405 211.770 ;
        RECT 2252.575 211.600 2252.865 211.770 ;
        RECT 2253.035 211.600 2253.325 211.770 ;
        RECT 2253.495 211.600 2253.785 211.770 ;
        RECT 2253.955 211.600 2254.245 211.770 ;
        RECT 2254.415 211.600 2254.705 211.770 ;
        RECT 2254.875 211.600 2255.165 211.770 ;
        RECT 2255.335 211.600 2255.625 211.770 ;
        RECT 2255.795 211.600 2256.085 211.770 ;
        RECT 2256.255 211.600 2256.545 211.770 ;
        RECT 2256.715 211.600 2257.005 211.770 ;
        RECT 2257.175 211.600 2257.465 211.770 ;
        RECT 2257.635 211.600 2257.925 211.770 ;
        RECT 2258.095 211.600 2258.385 211.770 ;
        RECT 2258.555 211.600 2258.845 211.770 ;
        RECT 2259.015 211.600 2259.305 211.770 ;
        RECT 2259.475 211.600 2259.765 211.770 ;
        RECT 2259.935 211.600 2260.225 211.770 ;
        RECT 2260.395 211.600 2260.685 211.770 ;
        RECT 2260.855 211.600 2261.145 211.770 ;
        RECT 2261.315 211.600 2261.605 211.770 ;
        RECT 2261.775 211.600 2262.065 211.770 ;
        RECT 2262.235 211.600 2262.525 211.770 ;
        RECT 2262.695 211.600 2262.985 211.770 ;
        RECT 2263.155 211.600 2263.445 211.770 ;
        RECT 2263.615 211.600 2263.905 211.770 ;
        RECT 2264.075 211.600 2264.365 211.770 ;
        RECT 2264.535 211.600 2264.825 211.770 ;
        RECT 2264.995 211.600 2265.285 211.770 ;
        RECT 2265.455 211.600 2265.745 211.770 ;
        RECT 2265.915 211.600 2266.205 211.770 ;
        RECT 2266.375 211.600 2266.665 211.770 ;
        RECT 2266.835 211.600 2267.125 211.770 ;
        RECT 2267.295 211.600 2267.585 211.770 ;
        RECT 2267.755 211.600 2268.045 211.770 ;
        RECT 2268.215 211.600 2268.505 211.770 ;
        RECT 2268.675 211.600 2268.965 211.770 ;
        RECT 2269.135 211.600 2269.425 211.770 ;
        RECT 2269.595 211.600 2269.885 211.770 ;
        RECT 2270.055 211.600 2270.345 211.770 ;
        RECT 2270.515 211.600 2270.805 211.770 ;
        RECT 2270.975 211.600 2271.265 211.770 ;
        RECT 2271.435 211.600 2271.725 211.770 ;
        RECT 2271.895 211.600 2272.040 211.770 ;
      LAYER mcon ;
        RECT 835.260 4984.800 836.350 4984.970 ;
        RECT 841.240 4984.800 842.330 4984.970 ;
        RECT 847.220 4984.800 848.310 4984.970 ;
        RECT 836.170 4981.400 836.340 4982.250 ;
        RECT 842.150 4981.400 842.320 4982.250 ;
        RECT 848.130 4981.400 848.300 4982.250 ;
        RECT 2087.580 4983.025 2087.750 4983.875 ;
        RECT 3311.355 4985.675 3311.525 4986.525 ;
        RECT 3309.945 4982.955 3311.035 4983.125 ;
        RECT 3314.585 4982.615 3314.755 4983.465 ;
        RECT 3320.565 4982.615 3320.735 4983.465 ;
        RECT 3326.545 4982.615 3326.715 4983.465 ;
        RECT 3332.525 4982.615 3332.695 4983.465 ;
        RECT 202.610 4455.510 203.460 4455.680 ;
        RECT 206.010 4456.000 206.180 4457.090 ;
        RECT 202.950 4451.370 203.120 4452.460 ;
        RECT 205.670 4452.280 206.520 4452.450 ;
        RECT 202.610 4449.530 203.460 4449.700 ;
        RECT 206.010 4450.020 206.180 4451.110 ;
        RECT 202.950 4445.390 203.120 4446.480 ;
        RECT 205.670 4446.300 206.520 4446.470 ;
        RECT 202.610 4443.550 203.460 4443.720 ;
        RECT 206.010 4444.040 206.180 4445.130 ;
        RECT 202.950 4439.410 203.120 4440.500 ;
        RECT 205.670 4440.320 206.520 4440.490 ;
        RECT 202.950 4433.430 203.120 4434.520 ;
        RECT 205.670 4434.340 206.520 4434.510 ;
        RECT 202.950 4427.450 203.120 4428.540 ;
        RECT 205.670 4428.360 206.520 4428.530 ;
        RECT 3381.690 3637.200 3381.860 3638.290 ;
        RECT 3381.350 3633.480 3382.200 3633.650 ;
        RECT 3384.750 3632.570 3384.920 3633.660 ;
        RECT 3381.690 3631.220 3381.860 3632.310 ;
        RECT 3381.350 3627.500 3382.200 3627.670 ;
        RECT 3384.750 3626.590 3384.920 3627.680 ;
        RECT 3381.690 3625.240 3381.860 3626.330 ;
        RECT 3381.350 3621.520 3382.200 3621.690 ;
        RECT 3384.750 3620.610 3384.920 3621.700 ;
        RECT 3381.690 3619.260 3381.860 3620.350 ;
        RECT 3381.350 3615.540 3382.200 3615.710 ;
        RECT 3384.750 3614.630 3384.920 3615.720 ;
        RECT 3381.350 3609.560 3382.200 3609.730 ;
        RECT 3384.750 3608.650 3384.920 3609.740 ;
        RECT 3381.350 3603.580 3382.200 3603.750 ;
        RECT 3384.750 3602.670 3384.920 3603.760 ;
        RECT 202.735 3049.280 203.585 3049.450 ;
        RECT 206.135 3049.770 206.305 3050.860 ;
        RECT 203.075 3045.140 203.245 3046.230 ;
        RECT 205.795 3046.050 206.645 3046.220 ;
        RECT 202.735 3043.300 203.585 3043.470 ;
        RECT 206.135 3043.790 206.305 3044.880 ;
        RECT 203.075 3039.160 203.245 3040.250 ;
        RECT 205.795 3040.070 206.645 3040.240 ;
        RECT 202.735 3037.320 203.585 3037.490 ;
        RECT 206.135 3037.810 206.305 3038.900 ;
        RECT 203.075 3033.180 203.245 3034.270 ;
        RECT 205.795 3034.090 206.645 3034.260 ;
        RECT 202.735 3031.340 203.585 3031.510 ;
        RECT 206.135 3031.830 206.305 3032.920 ;
        RECT 203.075 3027.200 203.245 3028.290 ;
        RECT 205.795 3028.110 206.645 3028.280 ;
        RECT 202.735 3025.360 203.585 3025.530 ;
        RECT 206.135 3025.850 206.305 3026.940 ;
        RECT 203.075 3021.220 203.245 3022.310 ;
        RECT 205.795 3022.130 206.645 3022.300 ;
        RECT 203.075 3015.240 203.245 3016.330 ;
        RECT 205.795 3016.150 206.645 3016.320 ;
        RECT 203.075 3009.260 203.245 3010.350 ;
        RECT 205.795 3010.170 206.645 3010.340 ;
        RECT 203.075 3003.280 203.245 3004.370 ;
        RECT 205.795 3004.190 206.645 3004.360 ;
        RECT 203.075 2997.300 203.245 2998.390 ;
        RECT 205.795 2998.210 206.645 2998.380 ;
        RECT 203.075 2991.320 203.245 2992.410 ;
        RECT 205.795 2992.230 206.645 2992.400 ;
        RECT 203.075 2985.340 203.245 2986.430 ;
        RECT 205.795 2986.250 206.645 2986.420 ;
        RECT 3381.690 2267.080 3381.860 2268.170 ;
        RECT 3381.690 2261.100 3381.860 2262.190 ;
        RECT 3381.690 2255.120 3381.860 2256.210 ;
        RECT 3381.690 2249.140 3381.860 2250.230 ;
        RECT 3381.690 2243.160 3381.860 2244.250 ;
        RECT 3381.690 2237.180 3381.860 2238.270 ;
        RECT 202.845 1761.375 203.695 1761.545 ;
        RECT 206.245 1761.865 206.415 1762.955 ;
        RECT 203.185 1757.235 203.355 1758.325 ;
        RECT 205.905 1758.145 206.755 1758.315 ;
        RECT 202.845 1755.395 203.695 1755.565 ;
        RECT 206.245 1755.885 206.415 1756.975 ;
        RECT 203.185 1751.255 203.355 1752.345 ;
        RECT 205.855 1752.165 206.705 1752.335 ;
        RECT 202.845 1749.415 203.695 1749.585 ;
        RECT 206.245 1749.905 206.415 1750.995 ;
        RECT 203.185 1745.275 203.355 1746.365 ;
        RECT 205.905 1746.185 206.755 1746.355 ;
        RECT 202.845 1743.435 203.695 1743.605 ;
        RECT 206.245 1743.925 206.415 1745.015 ;
        RECT 203.185 1739.295 203.355 1740.385 ;
        RECT 205.905 1740.205 206.755 1740.375 ;
        RECT 202.845 1737.455 203.695 1737.625 ;
        RECT 206.245 1737.945 206.415 1739.035 ;
        RECT 203.185 1733.315 203.355 1734.405 ;
        RECT 205.905 1734.225 206.755 1734.395 ;
        RECT 202.845 1731.475 203.695 1731.645 ;
        RECT 206.245 1731.965 206.415 1733.055 ;
        RECT 203.185 1727.335 203.355 1728.425 ;
        RECT 205.905 1728.245 206.755 1728.415 ;
        RECT 202.845 1725.495 203.695 1725.665 ;
        RECT 206.245 1725.985 206.415 1727.075 ;
        RECT 203.185 1721.355 203.355 1722.445 ;
        RECT 205.905 1722.265 206.755 1722.435 ;
        RECT 202.845 1719.515 203.695 1719.685 ;
        RECT 206.245 1720.005 206.415 1721.095 ;
        RECT 203.185 1715.375 203.355 1716.465 ;
        RECT 205.905 1716.285 206.755 1716.455 ;
        RECT 202.845 1713.535 203.695 1713.705 ;
        RECT 206.245 1714.025 206.415 1715.115 ;
        RECT 203.185 1709.395 203.355 1710.485 ;
        RECT 205.905 1710.305 206.755 1710.475 ;
        RECT 202.845 1707.555 203.695 1707.725 ;
        RECT 206.245 1708.045 206.415 1709.135 ;
        RECT 203.185 1703.415 203.355 1704.505 ;
        RECT 205.905 1704.325 206.755 1704.495 ;
        RECT 202.845 1701.575 203.695 1701.745 ;
        RECT 206.245 1702.065 206.415 1703.155 ;
        RECT 203.185 1697.435 203.355 1698.525 ;
        RECT 205.905 1698.345 206.755 1698.515 ;
        RECT 203.185 1691.455 203.355 1692.545 ;
        RECT 205.905 1692.365 206.755 1692.535 ;
        RECT 203.185 1685.475 203.355 1686.565 ;
        RECT 205.905 1686.385 206.755 1686.555 ;
        RECT 203.185 1679.495 203.355 1680.585 ;
        RECT 205.905 1680.405 206.755 1680.575 ;
        RECT 203.185 1673.515 203.355 1674.605 ;
        RECT 205.905 1674.425 206.755 1674.595 ;
        RECT 670.520 215.510 670.690 216.360 ;
        RECT 674.240 215.850 675.330 216.020 ;
        RECT 676.500 215.510 676.670 216.360 ;
        RECT 680.220 215.850 681.310 216.020 ;
        RECT 682.480 215.510 682.650 216.360 ;
        RECT 686.200 215.850 687.290 216.020 ;
        RECT 688.460 215.510 688.630 216.360 ;
        RECT 692.180 215.850 693.270 216.020 ;
        RECT 694.440 215.510 694.610 216.360 ;
        RECT 698.160 215.850 699.250 216.020 ;
        RECT 700.420 215.510 700.590 216.360 ;
        RECT 704.140 215.850 705.230 216.020 ;
        RECT 706.400 215.510 706.570 216.360 ;
        RECT 710.120 215.850 711.210 216.020 ;
        RECT 712.380 215.510 712.550 216.360 ;
        RECT 716.100 215.850 717.190 216.020 ;
        RECT 718.360 215.510 718.530 216.360 ;
        RECT 722.080 215.850 723.170 216.020 ;
        RECT 724.340 215.510 724.510 216.360 ;
        RECT 728.060 215.850 729.150 216.020 ;
        RECT 730.320 215.510 730.490 216.360 ;
        RECT 734.040 215.850 735.130 216.020 ;
        RECT 736.300 215.510 736.470 216.360 ;
        RECT 740.020 215.850 741.110 216.020 ;
        RECT 742.280 215.510 742.450 216.360 ;
        RECT 746.000 215.850 747.090 216.020 ;
        RECT 748.260 215.510 748.430 216.360 ;
        RECT 751.980 215.850 753.070 216.020 ;
        RECT 754.240 215.510 754.410 216.360 ;
        RECT 757.960 215.850 759.050 216.020 ;
        RECT 763.940 215.850 765.030 216.020 ;
        RECT 769.920 215.850 771.010 216.020 ;
        RECT 775.900 215.850 776.990 216.020 ;
        RECT 781.880 215.850 782.970 216.020 ;
        RECT 787.860 215.850 788.950 216.020 ;
        RECT 793.840 215.850 794.930 216.020 ;
        RECT 2147.520 215.510 2147.690 216.360 ;
        RECT 2153.500 215.510 2153.670 216.360 ;
        RECT 2159.480 215.510 2159.650 216.360 ;
        RECT 2165.460 215.510 2165.630 216.360 ;
        RECT 2171.440 215.510 2171.610 216.360 ;
        RECT 2177.420 215.510 2177.590 216.360 ;
        RECT 2183.400 215.510 2183.570 216.360 ;
        RECT 2189.380 215.510 2189.550 216.360 ;
        RECT 2195.360 215.510 2195.530 216.360 ;
        RECT 2201.340 215.510 2201.510 216.360 ;
        RECT 2207.320 215.510 2207.490 216.360 ;
        RECT 2213.300 215.510 2213.470 216.360 ;
        RECT 2219.280 215.510 2219.450 216.360 ;
        RECT 2225.260 215.510 2225.430 216.360 ;
        RECT 2231.240 215.510 2231.410 216.360 ;
        RECT 2237.220 215.510 2237.390 216.360 ;
        RECT 2243.200 215.510 2243.370 216.360 ;
        RECT 2249.180 215.510 2249.350 216.360 ;
        RECT 2255.160 215.510 2255.330 216.360 ;
        RECT 2261.140 215.510 2261.310 216.360 ;
        RECT 2267.120 215.510 2267.290 216.360 ;
        RECT 675.590 212.790 676.680 212.960 ;
        RECT 679.730 212.450 679.900 213.300 ;
        RECT 681.570 212.790 682.660 212.960 ;
        RECT 685.710 212.450 685.880 213.300 ;
        RECT 687.550 212.790 688.640 212.960 ;
        RECT 691.690 212.450 691.860 213.300 ;
        RECT 693.530 212.790 694.620 212.960 ;
        RECT 697.670 212.450 697.840 213.300 ;
        RECT 699.510 212.790 700.600 212.960 ;
        RECT 703.650 212.450 703.820 213.300 ;
        RECT 705.490 212.790 706.580 212.960 ;
        RECT 709.630 212.450 709.800 213.300 ;
        RECT 711.470 212.790 712.560 212.960 ;
        RECT 715.610 212.450 715.780 213.300 ;
        RECT 717.450 212.790 718.540 212.960 ;
        RECT 721.590 212.450 721.760 213.300 ;
        RECT 723.430 212.790 724.520 212.960 ;
        RECT 727.570 212.450 727.740 213.300 ;
        RECT 729.410 212.790 730.500 212.960 ;
        RECT 733.550 212.450 733.720 213.300 ;
        RECT 735.390 212.790 736.480 212.960 ;
        RECT 739.530 212.450 739.700 213.300 ;
        RECT 741.370 212.790 742.460 212.960 ;
        RECT 745.510 212.450 745.680 213.300 ;
        RECT 747.350 212.790 748.440 212.960 ;
        RECT 751.490 212.450 751.660 213.300 ;
        RECT 753.330 212.790 754.420 212.960 ;
        RECT 757.470 212.450 757.640 213.300 ;
        RECT 759.310 212.790 760.400 212.960 ;
        RECT 763.450 212.450 763.620 213.300 ;
        RECT 769.430 212.450 769.600 213.300 ;
        RECT 775.410 212.450 775.580 213.300 ;
        RECT 781.390 212.450 781.560 213.300 ;
        RECT 787.370 212.450 787.540 213.300 ;
        RECT 793.340 212.790 794.430 212.960 ;
        RECT 2152.590 212.790 2153.680 212.960 ;
        RECT 2158.570 212.790 2159.660 212.960 ;
        RECT 2164.550 212.790 2165.640 212.960 ;
        RECT 2170.530 212.790 2171.620 212.960 ;
        RECT 2176.510 212.790 2177.600 212.960 ;
        RECT 2182.490 212.790 2183.580 212.960 ;
        RECT 2188.470 212.790 2189.560 212.960 ;
        RECT 2194.450 212.790 2195.540 212.960 ;
        RECT 2200.430 212.790 2201.520 212.960 ;
        RECT 2206.410 212.790 2207.500 212.960 ;
        RECT 2212.390 212.790 2213.480 212.960 ;
        RECT 2218.370 212.790 2219.460 212.960 ;
        RECT 2224.350 212.790 2225.440 212.960 ;
        RECT 2230.330 212.790 2231.420 212.960 ;
        RECT 2236.310 212.790 2237.400 212.960 ;
        RECT 2242.290 212.790 2243.380 212.960 ;
        RECT 2248.270 212.790 2249.360 212.960 ;
        RECT 2254.250 212.790 2255.340 212.960 ;
        RECT 2260.230 212.790 2261.320 212.960 ;
        RECT 2267.120 212.450 2267.290 213.300 ;
      LAYER met1 ;
        RECT 2087.510 4986.375 2088.720 4986.635 ;
        RECT 3311.315 4985.615 3311.575 4986.585 ;
        RECT 3314.515 4985.965 3315.725 4986.225 ;
        RECT 3320.495 4985.965 3321.705 4986.225 ;
        RECT 3326.475 4985.965 3327.685 4986.225 ;
        RECT 3332.455 4985.965 3333.665 4986.225 ;
        RECT 835.200 4984.750 836.410 4985.010 ;
        RECT 841.180 4984.750 842.390 4985.010 ;
        RECT 847.160 4984.750 848.370 4985.010 ;
        RECT 2087.540 4982.965 2087.800 4983.935 ;
        RECT 3309.885 4982.905 3311.095 4983.165 ;
        RECT 3314.545 4982.555 3314.805 4983.525 ;
        RECT 3320.525 4982.555 3320.785 4983.525 ;
        RECT 3326.505 4982.555 3326.765 4983.525 ;
        RECT 3332.485 4982.555 3332.745 4983.525 ;
        RECT 836.120 4981.340 836.380 4982.310 ;
        RECT 842.100 4981.340 842.360 4982.310 ;
        RECT 848.080 4981.340 848.340 4982.310 ;
        RECT 211.175 4977.145 848.420 4977.285 ;
        RECT 205.970 4455.940 206.230 4457.150 ;
        RECT 211.175 4456.785 211.315 4977.145 ;
        RECT 848.100 4977.025 848.420 4977.145 ;
        RECT 211.055 4456.465 211.315 4456.785 ;
        RECT 211.455 4976.865 847.800 4977.005 ;
        RECT 211.455 4455.815 211.595 4976.865 ;
        RECT 847.480 4976.745 847.800 4976.865 ;
        RECT 3310.250 4976.795 3310.570 4976.915 ;
        RECT 2087.460 4976.655 3310.570 4976.795 ;
        RECT 3314.465 4976.795 3376.660 4976.935 ;
        RECT 3314.465 4976.675 3314.785 4976.795 ;
        RECT 2087.460 4976.535 2087.780 4976.655 ;
        RECT 3311.220 4976.515 3311.540 4976.635 ;
        RECT 2088.055 4976.375 3311.540 4976.515 ;
        RECT 3315.085 4976.515 3376.380 4976.655 ;
        RECT 3315.085 4976.395 3315.405 4976.515 ;
        RECT 2088.080 4976.255 2088.400 4976.375 ;
        RECT 202.550 4455.460 203.520 4455.720 ;
        RECT 211.335 4455.495 211.595 4455.815 ;
        RECT 212.295 4976.025 842.440 4976.165 ;
        RECT 202.910 4451.310 203.170 4452.520 ;
        RECT 205.610 4452.230 206.580 4452.490 ;
        RECT 211.035 4452.250 211.295 4452.570 ;
        RECT 205.970 4449.960 206.230 4451.170 ;
        RECT 202.550 4449.480 203.520 4449.740 ;
        RECT 202.910 4445.330 203.170 4446.540 ;
        RECT 205.610 4446.250 206.580 4446.510 ;
        RECT 205.970 4443.980 206.230 4445.190 ;
        RECT 202.550 4443.500 203.520 4443.760 ;
        RECT 202.910 4439.350 203.170 4440.560 ;
        RECT 205.610 4440.270 206.580 4440.530 ;
        RECT 202.910 4433.370 203.170 4434.580 ;
        RECT 205.610 4434.290 206.580 4434.550 ;
        RECT 202.910 4427.390 203.170 4428.600 ;
        RECT 205.610 4428.310 206.580 4428.570 ;
        RECT 206.095 3049.710 206.355 3050.920 ;
        RECT 211.035 3050.555 211.175 4452.250 ;
        RECT 210.915 3050.235 211.175 3050.555 ;
        RECT 211.315 4451.630 211.575 4451.950 ;
        RECT 211.315 3049.585 211.455 4451.630 ;
        RECT 212.295 4450.685 212.435 4976.025 ;
        RECT 842.120 4975.905 842.440 4976.025 ;
        RECT 212.175 4450.365 212.435 4450.685 ;
        RECT 212.575 4975.745 841.820 4975.885 ;
        RECT 212.575 4449.835 212.715 4975.745 ;
        RECT 841.500 4975.625 841.820 4975.745 ;
        RECT 3320.445 4975.675 3375.400 4975.815 ;
        RECT 3320.445 4975.555 3320.765 4975.675 ;
        RECT 3321.065 4975.395 3375.120 4975.535 ;
        RECT 3321.065 4975.275 3321.385 4975.395 ;
        RECT 212.455 4449.515 212.715 4449.835 ;
        RECT 213.415 4974.905 836.460 4975.045 ;
        RECT 202.675 3049.230 203.645 3049.490 ;
        RECT 211.195 3049.265 211.455 3049.585 ;
        RECT 212.155 4446.270 212.415 4446.590 ;
        RECT 203.035 3045.080 203.295 3046.290 ;
        RECT 205.735 3046.000 206.705 3046.260 ;
        RECT 210.895 3046.020 211.155 3046.340 ;
        RECT 206.095 3043.730 206.355 3044.940 ;
        RECT 202.675 3043.250 203.645 3043.510 ;
        RECT 203.035 3039.100 203.295 3040.310 ;
        RECT 205.735 3040.020 206.705 3040.280 ;
        RECT 206.095 3037.750 206.355 3038.960 ;
        RECT 202.675 3037.270 203.645 3037.530 ;
        RECT 203.035 3033.120 203.295 3034.330 ;
        RECT 205.735 3034.040 206.705 3034.300 ;
        RECT 206.095 3031.770 206.355 3032.980 ;
        RECT 202.675 3031.290 203.645 3031.550 ;
        RECT 203.035 3027.140 203.295 3028.350 ;
        RECT 205.735 3028.060 206.705 3028.320 ;
        RECT 206.095 3025.790 206.355 3027.000 ;
        RECT 202.675 3025.310 203.645 3025.570 ;
        RECT 203.035 3021.160 203.295 3022.370 ;
        RECT 205.735 3022.080 206.705 3022.340 ;
        RECT 203.035 3015.180 203.295 3016.390 ;
        RECT 205.735 3016.100 206.705 3016.360 ;
        RECT 203.035 3009.200 203.295 3010.410 ;
        RECT 205.735 3010.120 206.705 3010.380 ;
        RECT 203.035 3003.220 203.295 3004.430 ;
        RECT 205.735 3004.140 206.705 3004.400 ;
        RECT 203.035 2997.240 203.295 2998.450 ;
        RECT 205.735 2998.160 206.705 2998.420 ;
        RECT 203.035 2991.260 203.295 2992.470 ;
        RECT 205.735 2992.180 206.705 2992.440 ;
        RECT 203.035 2985.280 203.295 2986.490 ;
        RECT 205.735 2986.200 206.705 2986.460 ;
        RECT 206.205 1761.805 206.465 1763.015 ;
        RECT 210.895 1762.650 211.035 3046.020 ;
        RECT 210.775 1762.330 211.035 1762.650 ;
        RECT 211.175 3045.400 211.435 3045.720 ;
        RECT 211.175 1761.680 211.315 3045.400 ;
        RECT 212.155 3044.455 212.295 4446.270 ;
        RECT 212.035 3044.135 212.295 3044.455 ;
        RECT 212.435 4445.650 212.695 4445.970 ;
        RECT 212.435 3043.605 212.575 4445.650 ;
        RECT 213.415 4444.825 213.555 4974.905 ;
        RECT 836.140 4974.785 836.460 4974.905 ;
        RECT 213.295 4444.505 213.555 4444.825 ;
        RECT 213.695 4974.625 835.840 4974.765 ;
        RECT 213.695 4443.855 213.835 4974.625 ;
        RECT 835.520 4974.505 835.840 4974.625 ;
        RECT 3326.425 4974.555 3374.280 4974.695 ;
        RECT 3326.425 4974.435 3326.745 4974.555 ;
        RECT 3327.045 4974.275 3374.000 4974.415 ;
        RECT 3327.045 4974.155 3327.365 4974.275 ;
        RECT 3332.405 4973.435 3373.160 4973.575 ;
        RECT 3332.405 4973.315 3332.725 4973.435 ;
        RECT 3333.000 4973.155 3372.880 4973.295 ;
        RECT 3333.025 4973.035 3333.345 4973.155 ;
        RECT 213.575 4443.535 213.835 4443.855 ;
        RECT 212.315 3043.285 212.575 3043.605 ;
        RECT 213.275 4440.290 213.535 4440.610 ;
        RECT 202.785 1761.325 203.755 1761.585 ;
        RECT 211.055 1761.360 211.315 1761.680 ;
        RECT 212.015 3040.040 212.275 3040.360 ;
        RECT 203.145 1757.175 203.405 1758.385 ;
        RECT 205.845 1758.095 206.815 1758.355 ;
        RECT 210.755 1758.115 211.015 1758.435 ;
        RECT 206.205 1755.825 206.465 1757.035 ;
        RECT 202.785 1755.345 203.755 1755.605 ;
        RECT 203.145 1751.195 203.405 1752.405 ;
        RECT 205.795 1752.115 206.765 1752.375 ;
        RECT 206.205 1749.845 206.465 1751.055 ;
        RECT 202.785 1749.365 203.755 1749.625 ;
        RECT 203.145 1745.215 203.405 1746.425 ;
        RECT 205.845 1746.135 206.815 1746.395 ;
        RECT 206.205 1743.865 206.465 1745.075 ;
        RECT 202.785 1743.385 203.755 1743.645 ;
        RECT 203.145 1739.235 203.405 1740.445 ;
        RECT 205.845 1740.155 206.815 1740.415 ;
        RECT 206.205 1737.885 206.465 1739.095 ;
        RECT 202.785 1737.405 203.755 1737.665 ;
        RECT 203.145 1733.255 203.405 1734.465 ;
        RECT 205.845 1734.175 206.815 1734.435 ;
        RECT 206.205 1731.905 206.465 1733.115 ;
        RECT 202.785 1731.425 203.755 1731.685 ;
        RECT 203.145 1727.275 203.405 1728.485 ;
        RECT 205.845 1728.195 206.815 1728.455 ;
        RECT 206.205 1725.925 206.465 1727.135 ;
        RECT 202.785 1725.445 203.755 1725.705 ;
        RECT 203.145 1721.295 203.405 1722.505 ;
        RECT 205.845 1722.215 206.815 1722.475 ;
        RECT 206.205 1719.945 206.465 1721.155 ;
        RECT 202.785 1719.465 203.755 1719.725 ;
        RECT 203.145 1715.315 203.405 1716.525 ;
        RECT 205.845 1716.235 206.815 1716.495 ;
        RECT 206.205 1713.965 206.465 1715.175 ;
        RECT 202.785 1713.485 203.755 1713.745 ;
        RECT 203.145 1709.335 203.405 1710.545 ;
        RECT 205.845 1710.255 206.815 1710.515 ;
        RECT 206.205 1707.985 206.465 1709.195 ;
        RECT 202.785 1707.505 203.755 1707.765 ;
        RECT 203.145 1703.355 203.405 1704.565 ;
        RECT 205.845 1704.275 206.815 1704.535 ;
        RECT 206.205 1702.005 206.465 1703.215 ;
        RECT 202.785 1701.525 203.755 1701.785 ;
        RECT 203.145 1697.375 203.405 1698.585 ;
        RECT 205.845 1698.295 206.815 1698.555 ;
        RECT 203.145 1691.395 203.405 1692.605 ;
        RECT 205.845 1692.315 206.815 1692.575 ;
        RECT 203.145 1685.415 203.405 1686.625 ;
        RECT 205.845 1686.335 206.815 1686.595 ;
        RECT 203.145 1679.435 203.405 1680.645 ;
        RECT 205.845 1680.355 206.815 1680.615 ;
        RECT 203.145 1673.455 203.405 1674.665 ;
        RECT 205.845 1674.375 206.815 1674.635 ;
        RECT 210.755 225.940 210.895 1758.115 ;
        RECT 211.035 1757.495 211.295 1757.815 ;
        RECT 211.035 226.220 211.175 1757.495 ;
        RECT 212.015 1756.550 212.155 3040.040 ;
        RECT 211.895 1756.230 212.155 1756.550 ;
        RECT 212.295 3039.420 212.555 3039.740 ;
        RECT 212.295 1755.700 212.435 3039.420 ;
        RECT 213.275 3038.595 213.415 4440.290 ;
        RECT 213.155 3038.275 213.415 3038.595 ;
        RECT 213.555 4439.670 213.815 4439.990 ;
        RECT 213.555 3037.625 213.695 4439.670 ;
        RECT 213.435 3037.305 213.695 3037.625 ;
        RECT 214.395 4434.310 214.655 4434.630 ;
        RECT 212.175 1755.380 212.435 1755.700 ;
        RECT 213.135 3034.060 213.395 3034.380 ;
        RECT 211.875 1752.135 212.135 1752.455 ;
        RECT 211.875 226.780 212.015 1752.135 ;
        RECT 212.155 1751.515 212.415 1751.835 ;
        RECT 212.155 227.060 212.295 1751.515 ;
        RECT 213.135 1750.690 213.275 3034.060 ;
        RECT 213.015 1750.370 213.275 1750.690 ;
        RECT 213.415 3033.440 213.675 3033.760 ;
        RECT 213.415 1749.720 213.555 3033.440 ;
        RECT 214.395 3032.495 214.535 4434.310 ;
        RECT 214.275 3032.175 214.535 3032.495 ;
        RECT 214.675 4433.690 214.935 4434.010 ;
        RECT 214.675 3031.645 214.815 4433.690 ;
        RECT 214.555 3031.325 214.815 3031.645 ;
        RECT 215.515 4428.330 215.775 4428.650 ;
        RECT 213.295 1749.400 213.555 1749.720 ;
        RECT 214.255 3028.080 214.515 3028.400 ;
        RECT 212.995 1746.155 213.255 1746.475 ;
        RECT 212.995 227.620 213.135 1746.155 ;
        RECT 213.275 1745.535 213.535 1745.855 ;
        RECT 213.275 227.900 213.415 1745.535 ;
        RECT 214.255 1744.590 214.395 3028.080 ;
        RECT 214.135 1744.270 214.395 1744.590 ;
        RECT 214.535 3027.460 214.795 3027.780 ;
        RECT 214.535 1743.740 214.675 3027.460 ;
        RECT 215.515 3026.635 215.655 4428.330 ;
        RECT 215.395 3026.315 215.655 3026.635 ;
        RECT 215.795 4427.710 216.055 4428.030 ;
        RECT 215.795 3025.665 215.935 4427.710 ;
        RECT 3372.740 3619.075 3372.880 4973.155 ;
        RECT 3373.020 3620.045 3373.160 4973.435 ;
        RECT 3373.860 3625.055 3374.000 4974.275 ;
        RECT 3374.140 3626.025 3374.280 4974.555 ;
        RECT 3374.980 3631.035 3375.120 4975.395 ;
        RECT 3375.260 3632.005 3375.400 4975.675 ;
        RECT 3376.240 3637.015 3376.380 4976.515 ;
        RECT 3376.520 3637.865 3376.660 4976.795 ;
        RECT 3376.520 3637.545 3376.780 3637.865 ;
        RECT 3381.640 3637.140 3381.900 3638.350 ;
        RECT 3376.240 3636.695 3376.500 3637.015 ;
        RECT 3384.350 3636.660 3385.320 3636.920 ;
        RECT 3376.540 3633.450 3376.800 3633.770 ;
        RECT 3376.260 3632.830 3376.520 3633.150 ;
        RECT 3375.260 3631.685 3375.520 3632.005 ;
        RECT 3374.980 3630.715 3375.240 3631.035 ;
        RECT 3375.280 3627.470 3375.540 3627.790 ;
        RECT 3375.000 3626.850 3375.260 3627.170 ;
        RECT 3374.140 3625.705 3374.400 3626.025 ;
        RECT 3373.860 3624.735 3374.120 3625.055 ;
        RECT 3374.160 3621.490 3374.420 3621.810 ;
        RECT 3373.880 3620.870 3374.140 3621.190 ;
        RECT 3373.020 3619.725 3373.280 3620.045 ;
        RECT 3372.740 3618.755 3373.000 3619.075 ;
        RECT 3373.040 3615.510 3373.300 3615.830 ;
        RECT 3372.760 3614.890 3373.020 3615.210 ;
        RECT 3371.920 3609.530 3372.180 3609.850 ;
        RECT 3371.640 3608.910 3371.900 3609.230 ;
        RECT 3370.800 3603.550 3371.060 3603.870 ;
        RECT 3370.640 3603.250 3370.780 3603.275 ;
        RECT 3370.520 3602.930 3370.780 3603.250 ;
        RECT 215.675 3025.345 215.935 3025.665 ;
        RECT 214.415 1743.420 214.675 1743.740 ;
        RECT 215.375 3022.100 215.635 3022.420 ;
        RECT 214.115 1740.175 214.375 1740.495 ;
        RECT 214.115 228.460 214.255 1740.175 ;
        RECT 214.395 1739.555 214.655 1739.875 ;
        RECT 214.395 228.740 214.535 1739.555 ;
        RECT 215.375 1738.730 215.515 3022.100 ;
        RECT 215.255 1738.410 215.515 1738.730 ;
        RECT 215.655 3021.480 215.915 3021.800 ;
        RECT 215.655 1737.760 215.795 3021.480 ;
        RECT 215.535 1737.440 215.795 1737.760 ;
        RECT 216.495 3016.120 216.755 3016.440 ;
        RECT 215.235 1734.195 215.495 1734.515 ;
        RECT 215.235 229.300 215.375 1734.195 ;
        RECT 215.515 1733.575 215.775 1733.895 ;
        RECT 215.515 229.580 215.655 1733.575 ;
        RECT 216.495 1732.750 216.635 3016.120 ;
        RECT 216.375 1732.430 216.635 1732.750 ;
        RECT 216.775 3015.500 217.035 3015.820 ;
        RECT 216.775 1731.780 216.915 3015.500 ;
        RECT 216.655 1731.460 216.915 1731.780 ;
        RECT 217.615 3010.140 217.875 3010.460 ;
        RECT 216.355 1728.215 216.615 1728.535 ;
        RECT 216.355 230.140 216.495 1728.215 ;
        RECT 216.635 1727.595 216.895 1727.915 ;
        RECT 216.635 230.420 216.775 1727.595 ;
        RECT 217.615 1726.770 217.755 3010.140 ;
        RECT 217.495 1726.450 217.755 1726.770 ;
        RECT 217.895 3009.520 218.155 3009.840 ;
        RECT 217.895 1725.800 218.035 3009.520 ;
        RECT 217.775 1725.480 218.035 1725.800 ;
        RECT 218.735 3004.160 218.995 3004.480 ;
        RECT 217.475 1722.235 217.735 1722.555 ;
        RECT 217.475 230.980 217.615 1722.235 ;
        RECT 217.755 1721.615 218.015 1721.935 ;
        RECT 217.755 231.260 217.895 1721.615 ;
        RECT 218.735 1720.790 218.875 3004.160 ;
        RECT 218.615 1720.470 218.875 1720.790 ;
        RECT 219.015 3003.540 219.275 3003.860 ;
        RECT 219.015 1719.820 219.155 3003.540 ;
        RECT 218.895 1719.500 219.155 1719.820 ;
        RECT 219.855 2998.180 220.115 2998.500 ;
        RECT 218.595 1716.255 218.855 1716.575 ;
        RECT 218.595 231.820 218.735 1716.255 ;
        RECT 218.875 1715.635 219.135 1715.955 ;
        RECT 218.875 232.100 219.015 1715.635 ;
        RECT 219.855 1714.810 219.995 2998.180 ;
        RECT 219.735 1714.490 219.995 1714.810 ;
        RECT 220.135 2997.560 220.395 2997.880 ;
        RECT 220.135 1713.840 220.275 2997.560 ;
        RECT 220.015 1713.520 220.275 1713.840 ;
        RECT 220.975 2992.200 221.235 2992.520 ;
        RECT 219.715 1710.275 219.975 1710.595 ;
        RECT 219.715 232.660 219.855 1710.275 ;
        RECT 219.995 1709.655 220.255 1709.975 ;
        RECT 219.995 232.940 220.135 1709.655 ;
        RECT 220.975 1708.830 221.115 2992.200 ;
        RECT 220.855 1708.510 221.115 1708.830 ;
        RECT 221.255 2991.580 221.515 2991.900 ;
        RECT 221.255 1707.860 221.395 2991.580 ;
        RECT 221.135 1707.540 221.395 1707.860 ;
        RECT 222.095 2986.220 222.355 2986.540 ;
        RECT 220.835 1704.295 221.095 1704.615 ;
        RECT 220.835 233.500 220.975 1704.295 ;
        RECT 221.115 1703.675 221.375 1703.995 ;
        RECT 221.115 233.780 221.255 1703.675 ;
        RECT 222.095 1702.850 222.235 2986.220 ;
        RECT 221.975 1702.530 222.235 1702.850 ;
        RECT 222.375 2985.600 222.635 2985.920 ;
        RECT 222.375 1701.880 222.515 2985.600 ;
        RECT 3370.640 2236.995 3370.780 3602.930 ;
        RECT 3370.920 2237.965 3371.060 3603.550 ;
        RECT 3371.760 2242.975 3371.900 3608.910 ;
        RECT 3372.040 2243.945 3372.180 3609.530 ;
        RECT 3372.880 2248.955 3373.020 3614.890 ;
        RECT 3373.160 2249.805 3373.300 3615.510 ;
        RECT 3374.000 2254.935 3374.140 3620.870 ;
        RECT 3374.280 2255.905 3374.420 3621.490 ;
        RECT 3375.120 2260.915 3375.260 3626.850 ;
        RECT 3375.400 2261.765 3375.540 3627.470 ;
        RECT 3376.380 2266.895 3376.520 3632.830 ;
        RECT 3376.660 2267.865 3376.800 3633.450 ;
        RECT 3381.290 3633.430 3382.260 3633.690 ;
        RECT 3384.700 3632.510 3384.960 3633.720 ;
        RECT 3381.640 3631.160 3381.900 3632.370 ;
        RECT 3384.350 3630.680 3385.320 3630.940 ;
        RECT 3381.290 3627.450 3382.260 3627.710 ;
        RECT 3384.700 3626.530 3384.960 3627.740 ;
        RECT 3381.640 3625.180 3381.900 3626.390 ;
        RECT 3384.350 3624.700 3385.320 3624.960 ;
        RECT 3381.290 3621.470 3382.260 3621.730 ;
        RECT 3384.700 3620.550 3384.960 3621.760 ;
        RECT 3381.640 3619.200 3381.900 3620.410 ;
        RECT 3384.350 3618.720 3385.320 3618.980 ;
        RECT 3381.290 3615.490 3382.260 3615.750 ;
        RECT 3384.700 3614.570 3384.960 3615.780 ;
        RECT 3381.290 3609.510 3382.260 3609.770 ;
        RECT 3384.700 3608.590 3384.960 3609.800 ;
        RECT 3381.290 3603.530 3382.260 3603.790 ;
        RECT 3384.700 3602.610 3384.960 3603.820 ;
        RECT 3376.660 2267.545 3376.920 2267.865 ;
        RECT 3381.640 2267.020 3381.900 2268.230 ;
        RECT 3376.380 2266.575 3376.640 2266.895 ;
        RECT 3384.350 2266.540 3385.320 2266.800 ;
        RECT 3375.400 2261.445 3375.660 2261.765 ;
        RECT 3381.640 2261.040 3381.900 2262.250 ;
        RECT 3375.120 2260.595 3375.380 2260.915 ;
        RECT 3384.350 2260.560 3385.320 2260.820 ;
        RECT 3374.280 2255.585 3374.540 2255.905 ;
        RECT 3381.640 2255.060 3381.900 2256.270 ;
        RECT 3374.000 2254.615 3374.260 2254.935 ;
        RECT 3384.350 2254.580 3385.320 2254.840 ;
        RECT 3373.160 2249.485 3373.420 2249.805 ;
        RECT 3381.640 2249.080 3381.900 2250.290 ;
        RECT 3372.880 2248.635 3373.140 2248.955 ;
        RECT 3384.350 2248.600 3385.320 2248.860 ;
        RECT 3372.040 2243.625 3372.300 2243.945 ;
        RECT 3381.640 2243.100 3381.900 2244.310 ;
        RECT 3371.760 2242.655 3372.020 2242.975 ;
        RECT 3384.350 2242.620 3385.320 2242.880 ;
        RECT 3370.920 2237.645 3371.180 2237.965 ;
        RECT 3381.640 2237.120 3381.900 2238.330 ;
        RECT 3370.640 2236.675 3370.900 2236.995 ;
        RECT 3384.350 2236.640 3385.320 2236.900 ;
        RECT 222.255 1701.560 222.515 1701.880 ;
        RECT 221.955 1698.315 222.215 1698.635 ;
        RECT 221.955 234.340 222.095 1698.315 ;
        RECT 222.235 1697.695 222.495 1698.015 ;
        RECT 222.235 234.620 222.375 1697.695 ;
        RECT 223.075 1692.335 223.335 1692.655 ;
        RECT 223.075 235.180 223.215 1692.335 ;
        RECT 223.355 1691.715 223.615 1692.035 ;
        RECT 223.355 235.460 223.495 1691.715 ;
        RECT 224.195 1686.355 224.455 1686.675 ;
        RECT 224.195 236.020 224.335 1686.355 ;
        RECT 224.475 1685.735 224.735 1686.055 ;
        RECT 224.475 236.300 224.615 1685.735 ;
        RECT 225.315 1680.375 225.575 1680.695 ;
        RECT 225.315 236.860 225.455 1680.375 ;
        RECT 225.595 1679.755 225.855 1680.075 ;
        RECT 225.595 237.140 225.735 1679.755 ;
        RECT 226.435 1674.395 226.695 1674.715 ;
        RECT 226.435 237.700 226.575 1674.395 ;
        RECT 226.715 1673.775 226.975 1674.095 ;
        RECT 226.715 237.980 226.855 1673.775 ;
        RECT 2147.490 238.120 2147.810 238.240 ;
        RECT 670.490 237.980 670.810 238.100 ;
        RECT 226.715 237.840 670.810 237.980 ;
        RECT 674.705 237.980 706.345 238.120 ;
        RECT 674.705 237.860 675.025 237.980 ;
        RECT 675.850 237.700 676.170 237.820 ;
        RECT 226.435 237.560 676.170 237.700 ;
        RECT 679.715 237.700 706.065 237.840 ;
        RECT 679.715 237.580 680.035 237.700 ;
        RECT 676.470 237.140 676.790 237.260 ;
        RECT 225.595 237.000 676.790 237.140 ;
        RECT 680.685 237.140 705.505 237.280 ;
        RECT 680.685 237.020 681.005 237.140 ;
        RECT 681.830 236.860 682.150 236.980 ;
        RECT 225.315 236.720 682.150 236.860 ;
        RECT 685.695 236.860 705.225 237.000 ;
        RECT 685.695 236.740 686.015 236.860 ;
        RECT 682.450 236.300 682.770 236.420 ;
        RECT 224.475 236.160 682.770 236.300 ;
        RECT 686.665 236.300 704.665 236.440 ;
        RECT 686.665 236.180 686.985 236.300 ;
        RECT 687.810 236.020 688.130 236.140 ;
        RECT 224.195 235.880 688.130 236.020 ;
        RECT 691.675 236.020 704.385 236.160 ;
        RECT 691.675 235.900 691.995 236.020 ;
        RECT 688.430 235.460 688.750 235.580 ;
        RECT 223.355 235.320 688.750 235.460 ;
        RECT 692.645 235.460 703.825 235.600 ;
        RECT 692.645 235.340 692.965 235.460 ;
        RECT 693.790 235.180 694.110 235.300 ;
        RECT 223.075 235.040 694.110 235.180 ;
        RECT 697.655 235.180 703.545 235.320 ;
        RECT 697.655 235.060 697.975 235.180 ;
        RECT 694.410 234.620 694.730 234.740 ;
        RECT 222.235 234.480 694.730 234.620 ;
        RECT 698.625 234.620 703.255 234.760 ;
        RECT 698.625 234.500 698.945 234.620 ;
        RECT 699.770 234.340 700.090 234.460 ;
        RECT 221.955 234.200 700.090 234.340 ;
        RECT 700.390 233.780 700.710 233.900 ;
        RECT 221.115 233.640 700.710 233.780 ;
        RECT 220.835 233.360 702.925 233.500 ;
        RECT 219.995 232.800 702.630 232.940 ;
        RECT 219.715 232.520 702.310 232.660 ;
        RECT 218.875 231.960 702.015 232.100 ;
        RECT 218.595 231.680 701.735 231.820 ;
        RECT 217.755 231.120 701.435 231.260 ;
        RECT 217.475 230.840 701.155 230.980 ;
        RECT 701.015 230.420 701.155 230.840 ;
        RECT 701.295 230.700 701.435 231.120 ;
        RECT 701.595 230.980 701.735 231.680 ;
        RECT 701.875 231.260 702.015 231.960 ;
        RECT 702.170 231.540 702.310 232.520 ;
        RECT 702.490 231.820 702.630 232.800 ;
        RECT 702.785 232.100 702.925 233.360 ;
        RECT 703.115 233.080 703.255 234.620 ;
        RECT 703.405 233.360 703.545 235.180 ;
        RECT 703.685 233.640 703.825 235.460 ;
        RECT 704.245 233.920 704.385 236.020 ;
        RECT 704.525 234.200 704.665 236.300 ;
        RECT 705.085 234.480 705.225 236.860 ;
        RECT 705.365 234.760 705.505 237.140 ;
        RECT 705.925 235.040 706.065 237.700 ;
        RECT 706.205 235.320 706.345 237.980 ;
        RECT 778.015 237.980 2147.810 238.120 ;
        RECT 778.015 235.320 778.155 237.980 ;
        RECT 2152.850 237.840 2153.170 237.960 ;
        RECT 706.205 235.180 778.155 235.320 ;
        RECT 778.295 237.700 2153.170 237.840 ;
        RECT 778.295 235.040 778.435 237.700 ;
        RECT 2153.470 237.280 2153.790 237.400 ;
        RECT 705.925 234.900 778.435 235.040 ;
        RECT 778.855 237.140 2153.790 237.280 ;
        RECT 778.855 234.760 778.995 237.140 ;
        RECT 2158.830 237.000 2159.150 237.120 ;
        RECT 705.365 234.620 778.995 234.760 ;
        RECT 779.135 236.860 2159.150 237.000 ;
        RECT 779.135 234.480 779.275 236.860 ;
        RECT 2159.450 236.440 2159.770 236.560 ;
        RECT 705.085 234.340 779.275 234.480 ;
        RECT 779.695 236.300 2159.770 236.440 ;
        RECT 779.695 234.200 779.835 236.300 ;
        RECT 2164.810 236.160 2165.130 236.280 ;
        RECT 704.525 234.060 779.835 234.200 ;
        RECT 779.975 236.020 2165.130 236.160 ;
        RECT 779.975 233.920 780.115 236.020 ;
        RECT 2165.430 235.600 2165.750 235.720 ;
        RECT 704.245 233.780 780.115 233.920 ;
        RECT 780.535 235.460 2165.750 235.600 ;
        RECT 780.535 233.640 780.675 235.460 ;
        RECT 2170.790 235.320 2171.110 235.440 ;
        RECT 703.685 233.500 780.675 233.640 ;
        RECT 780.815 235.180 2171.110 235.320 ;
        RECT 780.815 233.360 780.955 235.180 ;
        RECT 2171.410 234.760 2171.730 234.880 ;
        RECT 703.405 233.220 780.955 233.360 ;
        RECT 781.375 234.620 2171.730 234.760 ;
        RECT 781.375 233.080 781.515 234.620 ;
        RECT 2176.770 234.480 2177.090 234.600 ;
        RECT 703.115 232.940 781.515 233.080 ;
        RECT 781.655 234.340 2177.090 234.480 ;
        RECT 781.655 232.800 781.795 234.340 ;
        RECT 2177.390 233.920 2177.710 234.040 ;
        RECT 703.635 232.660 781.795 232.800 ;
        RECT 782.215 233.780 2177.710 233.920 ;
        RECT 703.635 232.540 703.955 232.660 ;
        RECT 782.215 232.520 782.355 233.780 ;
        RECT 2182.750 233.640 2183.070 233.760 ;
        RECT 704.485 232.380 782.355 232.520 ;
        RECT 782.495 233.500 2183.070 233.640 ;
        RECT 704.485 232.260 704.805 232.380 ;
        RECT 782.495 232.240 782.635 233.500 ;
        RECT 2183.370 233.080 2183.690 233.200 ;
        RECT 705.750 232.100 706.070 232.220 ;
        RECT 702.785 231.960 706.070 232.100 ;
        RECT 709.615 232.100 782.635 232.240 ;
        RECT 783.055 232.940 2183.690 233.080 ;
        RECT 709.615 231.980 709.935 232.100 ;
        RECT 783.055 231.960 783.195 232.940 ;
        RECT 2188.730 232.800 2189.050 232.920 ;
        RECT 706.370 231.820 706.690 231.940 ;
        RECT 702.490 231.680 706.690 231.820 ;
        RECT 710.585 231.820 783.195 231.960 ;
        RECT 783.335 232.660 2189.050 232.800 ;
        RECT 710.585 231.700 710.905 231.820 ;
        RECT 783.335 231.680 783.475 232.660 ;
        RECT 2189.350 232.240 2189.670 232.360 ;
        RECT 711.730 231.540 712.050 231.660 ;
        RECT 702.170 231.400 712.050 231.540 ;
        RECT 715.595 231.540 783.475 231.680 ;
        RECT 783.895 232.100 2189.670 232.240 ;
        RECT 715.595 231.420 715.915 231.540 ;
        RECT 783.895 231.400 784.035 232.100 ;
        RECT 2194.710 231.960 2195.030 232.080 ;
        RECT 712.350 231.260 712.670 231.380 ;
        RECT 701.875 231.120 712.670 231.260 ;
        RECT 716.445 231.260 784.035 231.400 ;
        RECT 784.175 231.820 2195.030 231.960 ;
        RECT 716.445 231.140 716.765 231.260 ;
        RECT 784.175 231.120 784.315 231.820 ;
        RECT 2195.330 231.400 2195.650 231.520 ;
        RECT 717.710 230.980 718.030 231.100 ;
        RECT 701.595 230.840 718.030 230.980 ;
        RECT 721.575 230.980 784.315 231.120 ;
        RECT 784.735 231.260 2195.650 231.400 ;
        RECT 721.575 230.860 721.895 230.980 ;
        RECT 784.735 230.840 784.875 231.260 ;
        RECT 2200.690 231.120 2201.010 231.240 ;
        RECT 718.330 230.700 718.650 230.820 ;
        RECT 701.295 230.560 718.650 230.700 ;
        RECT 722.545 230.700 784.875 230.840 ;
        RECT 785.015 230.980 2201.010 231.120 ;
        RECT 722.545 230.580 722.865 230.700 ;
        RECT 785.015 230.560 785.155 230.980 ;
        RECT 2201.310 230.560 2201.630 230.680 ;
        RECT 723.690 230.420 724.010 230.540 ;
        RECT 216.635 230.280 700.840 230.420 ;
        RECT 701.015 230.280 724.010 230.420 ;
        RECT 727.555 230.420 785.155 230.560 ;
        RECT 785.360 230.420 2201.630 230.560 ;
        RECT 727.555 230.300 727.875 230.420 ;
        RECT 785.360 230.280 785.500 230.420 ;
        RECT 2206.670 230.280 2206.990 230.400 ;
        RECT 700.700 230.140 700.840 230.280 ;
        RECT 724.310 230.140 724.630 230.260 ;
        RECT 216.355 230.000 700.545 230.140 ;
        RECT 700.700 230.000 724.630 230.140 ;
        RECT 728.525 230.140 785.500 230.280 ;
        RECT 785.865 230.140 2206.990 230.280 ;
        RECT 728.525 230.020 728.845 230.140 ;
        RECT 785.865 230.000 786.005 230.140 ;
        RECT 700.405 229.860 700.545 230.000 ;
        RECT 729.670 229.860 729.990 229.980 ;
        RECT 700.405 229.720 729.990 229.860 ;
        RECT 733.535 229.860 786.005 230.000 ;
        RECT 733.535 229.740 733.855 229.860 ;
        RECT 2207.290 229.720 2207.610 229.840 ;
        RECT 730.290 229.580 730.610 229.700 ;
        RECT 215.515 229.440 730.610 229.580 ;
        RECT 734.505 229.580 2207.610 229.720 ;
        RECT 734.505 229.460 734.825 229.580 ;
        RECT 2212.650 229.440 2212.970 229.560 ;
        RECT 735.650 229.300 735.970 229.420 ;
        RECT 215.235 229.160 735.970 229.300 ;
        RECT 739.515 229.300 2212.970 229.440 ;
        RECT 739.515 229.180 739.835 229.300 ;
        RECT 2213.270 228.880 2213.590 229.000 ;
        RECT 736.270 228.740 736.590 228.860 ;
        RECT 214.395 228.600 736.590 228.740 ;
        RECT 740.485 228.740 2213.590 228.880 ;
        RECT 740.485 228.620 740.805 228.740 ;
        RECT 2218.630 228.600 2218.950 228.720 ;
        RECT 741.630 228.460 741.950 228.580 ;
        RECT 214.115 228.320 741.950 228.460 ;
        RECT 745.495 228.460 2218.950 228.600 ;
        RECT 745.495 228.340 745.815 228.460 ;
        RECT 2219.250 228.040 2219.570 228.160 ;
        RECT 742.250 227.900 742.570 228.020 ;
        RECT 213.275 227.760 742.570 227.900 ;
        RECT 746.465 227.900 2219.570 228.040 ;
        RECT 746.465 227.780 746.785 227.900 ;
        RECT 2224.610 227.760 2224.930 227.880 ;
        RECT 747.610 227.620 747.930 227.740 ;
        RECT 212.995 227.480 747.930 227.620 ;
        RECT 751.475 227.620 2224.930 227.760 ;
        RECT 751.475 227.500 751.795 227.620 ;
        RECT 2225.230 227.200 2225.550 227.320 ;
        RECT 748.230 227.060 748.550 227.180 ;
        RECT 212.155 226.920 748.550 227.060 ;
        RECT 752.445 227.060 2225.550 227.200 ;
        RECT 752.445 226.940 752.765 227.060 ;
        RECT 2230.590 226.920 2230.910 227.040 ;
        RECT 753.590 226.780 753.910 226.900 ;
        RECT 211.875 226.640 753.910 226.780 ;
        RECT 757.455 226.780 2230.910 226.920 ;
        RECT 757.455 226.660 757.775 226.780 ;
        RECT 2231.210 226.360 2231.530 226.480 ;
        RECT 754.210 226.220 754.530 226.340 ;
        RECT 211.035 226.080 754.530 226.220 ;
        RECT 758.425 226.220 2231.530 226.360 ;
        RECT 758.425 226.100 758.745 226.220 ;
        RECT 2236.570 226.080 2236.890 226.200 ;
        RECT 759.570 225.940 759.890 226.060 ;
        RECT 210.755 225.800 759.890 225.940 ;
        RECT 763.435 225.940 2236.890 226.080 ;
        RECT 763.435 225.820 763.755 225.940 ;
        RECT 2237.190 225.520 2237.510 225.640 ;
        RECT 764.405 225.380 2237.510 225.520 ;
        RECT 764.405 225.260 764.725 225.380 ;
        RECT 2242.550 225.240 2242.870 225.360 ;
        RECT 769.415 225.100 2242.870 225.240 ;
        RECT 769.415 224.980 769.735 225.100 ;
        RECT 2243.170 224.680 2243.490 224.800 ;
        RECT 770.385 224.540 2243.490 224.680 ;
        RECT 770.385 224.420 770.705 224.540 ;
        RECT 2248.530 224.400 2248.850 224.520 ;
        RECT 775.395 224.260 2248.850 224.400 ;
        RECT 775.395 224.140 775.715 224.260 ;
        RECT 2249.150 223.840 2249.470 223.960 ;
        RECT 776.245 223.700 2249.470 223.840 ;
        RECT 776.245 223.580 776.565 223.700 ;
        RECT 2254.510 223.560 2254.830 223.680 ;
        RECT 781.375 223.420 2254.830 223.560 ;
        RECT 781.375 223.300 781.695 223.420 ;
        RECT 2255.130 223.000 2255.450 223.120 ;
        RECT 782.345 222.860 2255.450 223.000 ;
        RECT 782.345 222.740 782.665 222.860 ;
        RECT 2260.490 222.720 2260.810 222.840 ;
        RECT 787.355 222.580 2260.810 222.720 ;
        RECT 787.355 222.460 787.675 222.580 ;
        RECT 2261.110 222.160 2261.430 222.280 ;
        RECT 788.205 222.020 2261.430 222.160 ;
        RECT 788.205 221.900 788.525 222.020 ;
        RECT 2266.470 221.600 2266.790 221.720 ;
        RECT 793.335 221.460 2266.790 221.600 ;
        RECT 793.335 221.340 793.655 221.460 ;
        RECT 2267.090 221.040 2267.410 221.160 ;
        RECT 794.305 220.900 2267.410 221.040 ;
        RECT 794.305 220.780 794.625 220.900 ;
        RECT 670.470 215.450 670.730 216.420 ;
        RECT 674.180 215.810 675.390 216.070 ;
        RECT 676.450 215.450 676.710 216.420 ;
        RECT 680.160 215.810 681.370 216.070 ;
        RECT 682.430 215.450 682.690 216.420 ;
        RECT 686.140 215.810 687.350 216.070 ;
        RECT 688.410 215.450 688.670 216.420 ;
        RECT 692.120 215.810 693.330 216.070 ;
        RECT 694.390 215.450 694.650 216.420 ;
        RECT 698.100 215.810 699.310 216.070 ;
        RECT 700.370 215.450 700.630 216.420 ;
        RECT 704.080 215.810 705.290 216.070 ;
        RECT 706.350 215.450 706.610 216.420 ;
        RECT 710.060 215.810 711.270 216.070 ;
        RECT 712.330 215.450 712.590 216.420 ;
        RECT 716.040 215.810 717.250 216.070 ;
        RECT 718.310 215.450 718.570 216.420 ;
        RECT 722.020 215.810 723.230 216.070 ;
        RECT 724.290 215.450 724.550 216.420 ;
        RECT 728.000 215.810 729.210 216.070 ;
        RECT 730.270 215.450 730.530 216.420 ;
        RECT 733.980 215.810 735.190 216.070 ;
        RECT 736.250 215.450 736.510 216.420 ;
        RECT 739.960 215.810 741.170 216.070 ;
        RECT 742.230 215.450 742.490 216.420 ;
        RECT 745.940 215.810 747.150 216.070 ;
        RECT 748.210 215.450 748.470 216.420 ;
        RECT 751.920 215.810 753.130 216.070 ;
        RECT 754.190 215.450 754.450 216.420 ;
        RECT 757.900 215.810 759.110 216.070 ;
        RECT 763.880 215.810 765.090 216.070 ;
        RECT 769.860 215.810 771.070 216.070 ;
        RECT 775.840 215.810 777.050 216.070 ;
        RECT 781.820 215.810 783.030 216.070 ;
        RECT 787.800 215.810 789.010 216.070 ;
        RECT 793.780 215.810 794.990 216.070 ;
        RECT 2147.470 215.450 2147.730 216.420 ;
        RECT 2153.450 215.450 2153.710 216.420 ;
        RECT 2159.430 215.450 2159.690 216.420 ;
        RECT 2165.410 215.450 2165.670 216.420 ;
        RECT 2171.390 215.450 2171.650 216.420 ;
        RECT 2177.370 215.450 2177.630 216.420 ;
        RECT 2183.350 215.450 2183.610 216.420 ;
        RECT 2189.330 215.450 2189.590 216.420 ;
        RECT 2195.310 215.450 2195.570 216.420 ;
        RECT 2201.290 215.450 2201.550 216.420 ;
        RECT 2207.270 215.450 2207.530 216.420 ;
        RECT 2213.250 215.450 2213.510 216.420 ;
        RECT 2219.230 215.450 2219.490 216.420 ;
        RECT 2225.210 215.450 2225.470 216.420 ;
        RECT 2231.190 215.450 2231.450 216.420 ;
        RECT 2237.170 215.450 2237.430 216.420 ;
        RECT 2243.150 215.450 2243.410 216.420 ;
        RECT 2249.130 215.450 2249.390 216.420 ;
        RECT 2255.110 215.450 2255.370 216.420 ;
        RECT 2261.090 215.450 2261.350 216.420 ;
        RECT 2267.070 215.450 2267.330 216.420 ;
        RECT 675.530 212.750 676.740 213.010 ;
        RECT 679.680 212.390 679.940 213.360 ;
        RECT 681.510 212.750 682.720 213.010 ;
        RECT 685.660 212.390 685.920 213.360 ;
        RECT 687.490 212.750 688.700 213.010 ;
        RECT 691.640 212.390 691.900 213.360 ;
        RECT 693.470 212.750 694.680 213.010 ;
        RECT 697.620 212.390 697.880 213.360 ;
        RECT 699.450 212.750 700.660 213.010 ;
        RECT 703.600 212.390 703.860 213.360 ;
        RECT 705.430 212.750 706.640 213.010 ;
        RECT 709.580 212.390 709.840 213.360 ;
        RECT 711.410 212.750 712.620 213.010 ;
        RECT 715.560 212.390 715.820 213.360 ;
        RECT 717.390 212.750 718.600 213.010 ;
        RECT 721.540 212.390 721.800 213.360 ;
        RECT 723.370 212.750 724.580 213.010 ;
        RECT 727.520 212.390 727.780 213.360 ;
        RECT 729.350 212.750 730.560 213.010 ;
        RECT 733.500 212.390 733.760 213.360 ;
        RECT 735.330 212.750 736.540 213.010 ;
        RECT 739.480 212.390 739.740 213.360 ;
        RECT 741.310 212.750 742.520 213.010 ;
        RECT 745.460 212.390 745.720 213.360 ;
        RECT 747.290 212.750 748.500 213.010 ;
        RECT 751.440 212.390 751.700 213.360 ;
        RECT 753.270 212.750 754.480 213.010 ;
        RECT 757.420 212.390 757.680 213.360 ;
        RECT 759.250 212.750 760.460 213.010 ;
        RECT 763.400 212.390 763.660 213.360 ;
        RECT 769.380 212.390 769.640 213.360 ;
        RECT 775.360 212.390 775.620 213.360 ;
        RECT 781.340 212.390 781.600 213.360 ;
        RECT 787.320 212.390 787.580 213.360 ;
        RECT 793.280 212.750 794.490 213.010 ;
        RECT 2152.530 212.750 2153.740 213.010 ;
        RECT 2158.510 212.750 2159.720 213.010 ;
        RECT 2164.490 212.750 2165.700 213.010 ;
        RECT 2170.470 212.750 2171.680 213.010 ;
        RECT 2176.450 212.750 2177.660 213.010 ;
        RECT 2182.430 212.750 2183.640 213.010 ;
        RECT 2188.410 212.750 2189.620 213.010 ;
        RECT 2194.390 212.750 2195.600 213.010 ;
        RECT 2200.370 212.750 2201.580 213.010 ;
        RECT 2206.350 212.750 2207.560 213.010 ;
        RECT 2212.330 212.750 2213.540 213.010 ;
        RECT 2218.310 212.750 2219.520 213.010 ;
        RECT 2224.290 212.750 2225.500 213.010 ;
        RECT 2230.270 212.750 2231.480 213.010 ;
        RECT 2236.250 212.750 2237.460 213.010 ;
        RECT 2242.230 212.750 2243.440 213.010 ;
        RECT 2248.210 212.750 2249.420 213.010 ;
        RECT 2254.190 212.750 2255.400 213.010 ;
        RECT 2260.170 212.750 2261.380 213.010 ;
        RECT 2267.080 212.390 2267.340 213.360 ;
      LAYER via ;
        RECT 2087.570 4986.375 2088.660 4986.635 ;
        RECT 3311.315 4985.675 3311.575 4986.525 ;
        RECT 3314.575 4985.965 3315.665 4986.225 ;
        RECT 3320.555 4985.965 3321.645 4986.225 ;
        RECT 3326.535 4985.965 3327.625 4986.225 ;
        RECT 3332.515 4985.965 3333.605 4986.225 ;
        RECT 835.260 4984.750 836.350 4985.010 ;
        RECT 841.240 4984.750 842.330 4985.010 ;
        RECT 847.220 4984.750 848.310 4985.010 ;
        RECT 2087.540 4983.025 2087.800 4983.875 ;
        RECT 3309.945 4982.905 3311.035 4983.165 ;
        RECT 3314.545 4982.615 3314.805 4983.465 ;
        RECT 3320.525 4982.615 3320.785 4983.465 ;
        RECT 3326.505 4982.615 3326.765 4983.465 ;
        RECT 3332.485 4982.615 3332.745 4983.465 ;
        RECT 836.120 4981.400 836.380 4982.250 ;
        RECT 842.100 4981.400 842.360 4982.250 ;
        RECT 848.080 4981.400 848.340 4982.250 ;
        RECT 205.970 4456.000 206.230 4457.090 ;
        RECT 848.130 4977.025 848.390 4977.285 ;
        RECT 211.055 4456.495 211.315 4456.755 ;
        RECT 847.510 4976.745 847.770 4977.005 ;
        RECT 2087.490 4976.535 2087.750 4976.795 ;
        RECT 3310.280 4976.655 3310.540 4976.915 ;
        RECT 3314.495 4976.675 3314.755 4976.935 ;
        RECT 2088.110 4976.255 2088.370 4976.515 ;
        RECT 3311.250 4976.375 3311.510 4976.635 ;
        RECT 3315.115 4976.395 3315.375 4976.655 ;
        RECT 202.610 4455.460 203.460 4455.720 ;
        RECT 211.335 4455.525 211.595 4455.785 ;
        RECT 202.910 4451.370 203.170 4452.460 ;
        RECT 205.670 4452.230 206.520 4452.490 ;
        RECT 211.035 4452.280 211.295 4452.540 ;
        RECT 205.970 4450.020 206.230 4451.110 ;
        RECT 202.610 4449.480 203.460 4449.740 ;
        RECT 202.910 4445.390 203.170 4446.480 ;
        RECT 205.670 4446.250 206.520 4446.510 ;
        RECT 205.970 4444.040 206.230 4445.130 ;
        RECT 202.610 4443.500 203.460 4443.760 ;
        RECT 202.910 4439.410 203.170 4440.500 ;
        RECT 205.670 4440.270 206.520 4440.530 ;
        RECT 202.910 4433.430 203.170 4434.520 ;
        RECT 205.670 4434.290 206.520 4434.550 ;
        RECT 202.910 4427.450 203.170 4428.540 ;
        RECT 205.670 4428.310 206.520 4428.570 ;
        RECT 206.095 3049.770 206.355 3050.860 ;
        RECT 210.915 3050.265 211.175 3050.525 ;
        RECT 211.315 4451.660 211.575 4451.920 ;
        RECT 842.150 4975.905 842.410 4976.165 ;
        RECT 212.175 4450.395 212.435 4450.655 ;
        RECT 841.530 4975.625 841.790 4975.885 ;
        RECT 3320.475 4975.555 3320.735 4975.815 ;
        RECT 3321.095 4975.275 3321.355 4975.535 ;
        RECT 212.455 4449.545 212.715 4449.805 ;
        RECT 202.735 3049.230 203.585 3049.490 ;
        RECT 211.195 3049.295 211.455 3049.555 ;
        RECT 212.155 4446.300 212.415 4446.560 ;
        RECT 203.035 3045.140 203.295 3046.230 ;
        RECT 205.795 3046.000 206.645 3046.260 ;
        RECT 210.895 3046.050 211.155 3046.310 ;
        RECT 206.095 3043.790 206.355 3044.880 ;
        RECT 202.735 3043.250 203.585 3043.510 ;
        RECT 203.035 3039.160 203.295 3040.250 ;
        RECT 205.795 3040.020 206.645 3040.280 ;
        RECT 206.095 3037.810 206.355 3038.900 ;
        RECT 202.735 3037.270 203.585 3037.530 ;
        RECT 203.035 3033.180 203.295 3034.270 ;
        RECT 205.795 3034.040 206.645 3034.300 ;
        RECT 206.095 3031.830 206.355 3032.920 ;
        RECT 202.735 3031.290 203.585 3031.550 ;
        RECT 203.035 3027.200 203.295 3028.290 ;
        RECT 205.795 3028.060 206.645 3028.320 ;
        RECT 206.095 3025.850 206.355 3026.940 ;
        RECT 202.735 3025.310 203.585 3025.570 ;
        RECT 203.035 3021.220 203.295 3022.310 ;
        RECT 205.795 3022.080 206.645 3022.340 ;
        RECT 203.035 3015.240 203.295 3016.330 ;
        RECT 205.795 3016.100 206.645 3016.360 ;
        RECT 203.035 3009.260 203.295 3010.350 ;
        RECT 205.795 3010.120 206.645 3010.380 ;
        RECT 203.035 3003.280 203.295 3004.370 ;
        RECT 205.795 3004.140 206.645 3004.400 ;
        RECT 203.035 2997.300 203.295 2998.390 ;
        RECT 205.795 2998.160 206.645 2998.420 ;
        RECT 203.035 2991.320 203.295 2992.410 ;
        RECT 205.795 2992.180 206.645 2992.440 ;
        RECT 203.035 2985.340 203.295 2986.430 ;
        RECT 205.795 2986.200 206.645 2986.460 ;
        RECT 206.205 1761.865 206.465 1762.955 ;
        RECT 210.775 1762.360 211.035 1762.620 ;
        RECT 211.175 3045.430 211.435 3045.690 ;
        RECT 212.035 3044.165 212.295 3044.425 ;
        RECT 212.435 4445.680 212.695 4445.940 ;
        RECT 836.170 4974.785 836.430 4975.045 ;
        RECT 213.295 4444.535 213.555 4444.795 ;
        RECT 835.550 4974.505 835.810 4974.765 ;
        RECT 3326.455 4974.435 3326.715 4974.695 ;
        RECT 3327.075 4974.155 3327.335 4974.415 ;
        RECT 3332.435 4973.315 3332.695 4973.575 ;
        RECT 3333.055 4973.035 3333.315 4973.295 ;
        RECT 213.575 4443.565 213.835 4443.825 ;
        RECT 212.315 3043.315 212.575 3043.575 ;
        RECT 213.275 4440.320 213.535 4440.580 ;
        RECT 202.845 1761.325 203.695 1761.585 ;
        RECT 211.055 1761.390 211.315 1761.650 ;
        RECT 212.015 3040.070 212.275 3040.330 ;
        RECT 203.145 1757.235 203.405 1758.325 ;
        RECT 205.905 1758.095 206.755 1758.355 ;
        RECT 210.755 1758.145 211.015 1758.405 ;
        RECT 206.205 1755.885 206.465 1756.975 ;
        RECT 202.845 1755.345 203.695 1755.605 ;
        RECT 203.145 1751.255 203.405 1752.345 ;
        RECT 205.855 1752.115 206.705 1752.375 ;
        RECT 206.205 1749.905 206.465 1750.995 ;
        RECT 202.845 1749.365 203.695 1749.625 ;
        RECT 203.145 1745.275 203.405 1746.365 ;
        RECT 205.905 1746.135 206.755 1746.395 ;
        RECT 206.205 1743.925 206.465 1745.015 ;
        RECT 202.845 1743.385 203.695 1743.645 ;
        RECT 203.145 1739.295 203.405 1740.385 ;
        RECT 205.905 1740.155 206.755 1740.415 ;
        RECT 206.205 1737.945 206.465 1739.035 ;
        RECT 202.845 1737.405 203.695 1737.665 ;
        RECT 203.145 1733.315 203.405 1734.405 ;
        RECT 205.905 1734.175 206.755 1734.435 ;
        RECT 206.205 1731.965 206.465 1733.055 ;
        RECT 202.845 1731.425 203.695 1731.685 ;
        RECT 203.145 1727.335 203.405 1728.425 ;
        RECT 205.905 1728.195 206.755 1728.455 ;
        RECT 206.205 1725.985 206.465 1727.075 ;
        RECT 202.845 1725.445 203.695 1725.705 ;
        RECT 203.145 1721.355 203.405 1722.445 ;
        RECT 205.905 1722.215 206.755 1722.475 ;
        RECT 206.205 1720.005 206.465 1721.095 ;
        RECT 202.845 1719.465 203.695 1719.725 ;
        RECT 203.145 1715.805 203.405 1716.465 ;
        RECT 205.905 1716.235 206.755 1716.495 ;
        RECT 203.145 1715.375 203.405 1715.665 ;
        RECT 206.205 1714.025 206.465 1715.115 ;
        RECT 202.845 1713.485 203.695 1713.745 ;
        RECT 203.145 1709.395 203.405 1710.485 ;
        RECT 205.905 1710.255 206.755 1710.515 ;
        RECT 206.205 1708.045 206.465 1709.135 ;
        RECT 202.845 1707.505 203.695 1707.765 ;
        RECT 203.145 1703.415 203.405 1704.505 ;
        RECT 205.905 1704.275 206.755 1704.535 ;
        RECT 206.205 1702.065 206.465 1703.155 ;
        RECT 202.845 1701.525 203.695 1701.785 ;
        RECT 203.145 1697.435 203.405 1698.525 ;
        RECT 205.905 1698.295 206.755 1698.555 ;
        RECT 203.145 1691.455 203.405 1692.545 ;
        RECT 205.905 1692.315 206.755 1692.575 ;
        RECT 203.145 1685.475 203.405 1686.565 ;
        RECT 205.905 1686.335 206.755 1686.595 ;
        RECT 203.145 1679.495 203.405 1680.585 ;
        RECT 205.905 1680.355 206.755 1680.615 ;
        RECT 203.145 1673.515 203.405 1674.605 ;
        RECT 205.905 1674.375 206.755 1674.635 ;
        RECT 211.035 1757.525 211.295 1757.785 ;
        RECT 211.895 1756.260 212.155 1756.520 ;
        RECT 212.295 3039.450 212.555 3039.710 ;
        RECT 213.155 3038.305 213.415 3038.565 ;
        RECT 213.555 4439.700 213.815 4439.960 ;
        RECT 213.435 3037.335 213.695 3037.595 ;
        RECT 214.395 4434.340 214.655 4434.600 ;
        RECT 212.175 1755.410 212.435 1755.670 ;
        RECT 213.135 3034.090 213.395 3034.350 ;
        RECT 211.875 1752.165 212.135 1752.425 ;
        RECT 212.155 1751.545 212.415 1751.805 ;
        RECT 213.015 1750.400 213.275 1750.660 ;
        RECT 213.415 3033.470 213.675 3033.730 ;
        RECT 214.275 3032.205 214.535 3032.465 ;
        RECT 214.675 4433.720 214.935 4433.980 ;
        RECT 214.555 3031.355 214.815 3031.615 ;
        RECT 215.515 4428.360 215.775 4428.620 ;
        RECT 213.295 1749.430 213.555 1749.690 ;
        RECT 214.255 3028.110 214.515 3028.370 ;
        RECT 212.995 1746.185 213.255 1746.445 ;
        RECT 213.275 1745.565 213.535 1745.825 ;
        RECT 214.135 1744.300 214.395 1744.560 ;
        RECT 214.535 3027.490 214.795 3027.750 ;
        RECT 215.395 3026.345 215.655 3026.605 ;
        RECT 215.795 4427.740 216.055 4428.000 ;
        RECT 3376.520 3637.575 3376.780 3637.835 ;
        RECT 3381.640 3637.200 3381.900 3638.290 ;
        RECT 3376.240 3636.725 3376.500 3636.985 ;
        RECT 3384.410 3636.660 3385.260 3636.920 ;
        RECT 3376.540 3633.480 3376.800 3633.740 ;
        RECT 3376.260 3632.860 3376.520 3633.120 ;
        RECT 3375.260 3631.715 3375.520 3631.975 ;
        RECT 3374.980 3630.745 3375.240 3631.005 ;
        RECT 3375.280 3627.500 3375.540 3627.760 ;
        RECT 3375.000 3626.880 3375.260 3627.140 ;
        RECT 3374.140 3625.735 3374.400 3625.995 ;
        RECT 3373.860 3624.765 3374.120 3625.025 ;
        RECT 3374.160 3621.520 3374.420 3621.780 ;
        RECT 3373.880 3620.900 3374.140 3621.160 ;
        RECT 3373.020 3619.755 3373.280 3620.015 ;
        RECT 3372.740 3618.785 3373.000 3619.045 ;
        RECT 3373.040 3615.540 3373.300 3615.800 ;
        RECT 3372.760 3614.920 3373.020 3615.180 ;
        RECT 3371.920 3609.560 3372.180 3609.820 ;
        RECT 3371.640 3608.940 3371.900 3609.200 ;
        RECT 3370.800 3603.580 3371.060 3603.840 ;
        RECT 3370.520 3602.960 3370.780 3603.220 ;
        RECT 215.675 3025.375 215.935 3025.635 ;
        RECT 214.415 1743.450 214.675 1743.710 ;
        RECT 215.375 3022.130 215.635 3022.390 ;
        RECT 214.115 1740.205 214.375 1740.465 ;
        RECT 214.395 1739.585 214.655 1739.845 ;
        RECT 215.255 1738.440 215.515 1738.700 ;
        RECT 215.655 3021.510 215.915 3021.770 ;
        RECT 215.535 1737.470 215.795 1737.730 ;
        RECT 216.495 3016.150 216.755 3016.410 ;
        RECT 215.235 1734.225 215.495 1734.485 ;
        RECT 215.515 1733.605 215.775 1733.865 ;
        RECT 216.375 1732.460 216.635 1732.720 ;
        RECT 216.775 3015.530 217.035 3015.790 ;
        RECT 216.655 1731.490 216.915 1731.750 ;
        RECT 217.615 3010.170 217.875 3010.430 ;
        RECT 216.355 1728.245 216.615 1728.505 ;
        RECT 216.635 1727.625 216.895 1727.885 ;
        RECT 217.495 1726.480 217.755 1726.740 ;
        RECT 217.895 3009.550 218.155 3009.810 ;
        RECT 217.775 1725.510 218.035 1725.770 ;
        RECT 218.735 3004.190 218.995 3004.450 ;
        RECT 217.475 1722.265 217.735 1722.525 ;
        RECT 217.755 1721.645 218.015 1721.905 ;
        RECT 218.615 1720.500 218.875 1720.760 ;
        RECT 219.015 3003.570 219.275 3003.830 ;
        RECT 218.895 1719.530 219.155 1719.790 ;
        RECT 219.855 2998.210 220.115 2998.470 ;
        RECT 218.595 1716.285 218.855 1716.545 ;
        RECT 218.875 1715.665 219.135 1715.925 ;
        RECT 219.735 1714.520 219.995 1714.780 ;
        RECT 220.135 2997.590 220.395 2997.850 ;
        RECT 220.015 1713.550 220.275 1713.810 ;
        RECT 220.975 2992.230 221.235 2992.490 ;
        RECT 219.715 1710.305 219.975 1710.565 ;
        RECT 219.995 1709.685 220.255 1709.945 ;
        RECT 220.855 1708.540 221.115 1708.800 ;
        RECT 221.255 2991.610 221.515 2991.870 ;
        RECT 221.135 1707.570 221.395 1707.830 ;
        RECT 222.095 2986.250 222.355 2986.510 ;
        RECT 220.835 1704.325 221.095 1704.585 ;
        RECT 221.115 1703.705 221.375 1703.965 ;
        RECT 221.975 1702.560 222.235 1702.820 ;
        RECT 222.375 2985.630 222.635 2985.890 ;
        RECT 3381.350 3633.430 3382.200 3633.690 ;
        RECT 3384.700 3632.570 3384.960 3633.660 ;
        RECT 3381.640 3631.220 3381.900 3632.310 ;
        RECT 3384.410 3630.680 3385.260 3630.940 ;
        RECT 3381.350 3627.450 3382.200 3627.710 ;
        RECT 3384.700 3626.590 3384.960 3627.680 ;
        RECT 3381.640 3625.240 3381.900 3626.330 ;
        RECT 3384.410 3624.700 3385.260 3624.960 ;
        RECT 3381.350 3621.470 3382.200 3621.730 ;
        RECT 3384.700 3620.610 3384.960 3621.700 ;
        RECT 3381.640 3619.260 3381.900 3620.350 ;
        RECT 3384.410 3618.720 3385.260 3618.980 ;
        RECT 3381.350 3615.490 3382.200 3615.750 ;
        RECT 3384.700 3614.630 3384.960 3615.720 ;
        RECT 3381.350 3609.510 3382.200 3609.770 ;
        RECT 3384.700 3608.650 3384.960 3609.740 ;
        RECT 3381.350 3603.530 3382.200 3603.790 ;
        RECT 3384.700 3602.670 3384.960 3603.760 ;
        RECT 3376.660 2267.575 3376.920 2267.835 ;
        RECT 3381.640 2267.080 3381.900 2268.170 ;
        RECT 3376.380 2266.605 3376.640 2266.865 ;
        RECT 3384.410 2266.540 3385.260 2266.800 ;
        RECT 3375.400 2261.475 3375.660 2261.735 ;
        RECT 3381.640 2261.100 3381.900 2262.190 ;
        RECT 3375.120 2260.625 3375.380 2260.885 ;
        RECT 3384.410 2260.560 3385.260 2260.820 ;
        RECT 3374.280 2255.615 3374.540 2255.875 ;
        RECT 3381.640 2255.120 3381.900 2256.210 ;
        RECT 3374.000 2254.645 3374.260 2254.905 ;
        RECT 3384.410 2254.580 3385.260 2254.840 ;
        RECT 3373.160 2249.515 3373.420 2249.775 ;
        RECT 3381.640 2249.140 3381.900 2250.230 ;
        RECT 3372.880 2248.665 3373.140 2248.925 ;
        RECT 3384.410 2248.600 3385.260 2248.860 ;
        RECT 3372.040 2243.655 3372.300 2243.915 ;
        RECT 3381.640 2243.160 3381.900 2244.250 ;
        RECT 3371.760 2242.685 3372.020 2242.945 ;
        RECT 3384.410 2242.620 3385.260 2242.880 ;
        RECT 3370.920 2237.675 3371.180 2237.935 ;
        RECT 3381.640 2237.180 3381.900 2238.270 ;
        RECT 3370.640 2236.705 3370.900 2236.965 ;
        RECT 3384.410 2236.640 3385.260 2236.900 ;
        RECT 222.255 1701.590 222.515 1701.850 ;
        RECT 221.955 1698.345 222.215 1698.605 ;
        RECT 222.235 1697.725 222.495 1697.985 ;
        RECT 223.075 1692.365 223.335 1692.625 ;
        RECT 223.355 1691.745 223.615 1692.005 ;
        RECT 224.195 1686.385 224.455 1686.645 ;
        RECT 224.475 1685.765 224.735 1686.025 ;
        RECT 225.315 1680.405 225.575 1680.665 ;
        RECT 225.595 1679.785 225.855 1680.045 ;
        RECT 226.435 1674.425 226.695 1674.685 ;
        RECT 226.715 1673.805 226.975 1674.065 ;
        RECT 670.520 237.840 670.780 238.100 ;
        RECT 674.735 237.860 674.995 238.120 ;
        RECT 675.880 237.560 676.140 237.820 ;
        RECT 679.745 237.580 680.005 237.840 ;
        RECT 676.500 237.000 676.760 237.260 ;
        RECT 680.715 237.020 680.975 237.280 ;
        RECT 681.860 236.720 682.120 236.980 ;
        RECT 685.725 236.740 685.985 237.000 ;
        RECT 682.480 236.160 682.740 236.420 ;
        RECT 686.695 236.180 686.955 236.440 ;
        RECT 687.840 235.880 688.100 236.140 ;
        RECT 691.705 235.900 691.965 236.160 ;
        RECT 688.460 235.320 688.720 235.580 ;
        RECT 692.675 235.340 692.935 235.600 ;
        RECT 693.820 235.040 694.080 235.300 ;
        RECT 697.685 235.060 697.945 235.320 ;
        RECT 694.440 234.480 694.700 234.740 ;
        RECT 698.655 234.500 698.915 234.760 ;
        RECT 699.800 234.200 700.060 234.460 ;
        RECT 700.420 233.640 700.680 233.900 ;
        RECT 2147.520 237.980 2147.780 238.240 ;
        RECT 2152.880 237.700 2153.140 237.960 ;
        RECT 2153.500 237.140 2153.760 237.400 ;
        RECT 2158.860 236.860 2159.120 237.120 ;
        RECT 2159.480 236.300 2159.740 236.560 ;
        RECT 2164.840 236.020 2165.100 236.280 ;
        RECT 2165.460 235.460 2165.720 235.720 ;
        RECT 2170.820 235.180 2171.080 235.440 ;
        RECT 2171.440 234.620 2171.700 234.880 ;
        RECT 2176.800 234.340 2177.060 234.600 ;
        RECT 703.665 232.540 703.925 232.800 ;
        RECT 2177.420 233.780 2177.680 234.040 ;
        RECT 704.515 232.260 704.775 232.520 ;
        RECT 2182.780 233.500 2183.040 233.760 ;
        RECT 705.780 231.960 706.040 232.220 ;
        RECT 709.645 231.980 709.905 232.240 ;
        RECT 2183.400 232.940 2183.660 233.200 ;
        RECT 706.400 231.680 706.660 231.940 ;
        RECT 710.615 231.700 710.875 231.960 ;
        RECT 2188.760 232.660 2189.020 232.920 ;
        RECT 711.760 231.400 712.020 231.660 ;
        RECT 715.625 231.420 715.885 231.680 ;
        RECT 2189.380 232.100 2189.640 232.360 ;
        RECT 712.380 231.120 712.640 231.380 ;
        RECT 716.475 231.140 716.735 231.400 ;
        RECT 2194.740 231.820 2195.000 232.080 ;
        RECT 717.740 230.840 718.000 231.100 ;
        RECT 721.605 230.860 721.865 231.120 ;
        RECT 2195.360 231.260 2195.620 231.520 ;
        RECT 718.360 230.560 718.620 230.820 ;
        RECT 722.575 230.580 722.835 230.840 ;
        RECT 2200.720 230.980 2200.980 231.240 ;
        RECT 723.720 230.280 723.980 230.540 ;
        RECT 727.585 230.300 727.845 230.560 ;
        RECT 2201.340 230.420 2201.600 230.680 ;
        RECT 724.340 230.000 724.600 230.260 ;
        RECT 728.555 230.020 728.815 230.280 ;
        RECT 2206.700 230.140 2206.960 230.400 ;
        RECT 729.700 229.720 729.960 229.980 ;
        RECT 733.565 229.740 733.825 230.000 ;
        RECT 730.320 229.440 730.580 229.700 ;
        RECT 734.535 229.460 734.795 229.720 ;
        RECT 2207.320 229.580 2207.580 229.840 ;
        RECT 735.680 229.160 735.940 229.420 ;
        RECT 739.545 229.180 739.805 229.440 ;
        RECT 2212.680 229.300 2212.940 229.560 ;
        RECT 736.300 228.600 736.560 228.860 ;
        RECT 740.515 228.620 740.775 228.880 ;
        RECT 2213.300 228.740 2213.560 229.000 ;
        RECT 741.660 228.320 741.920 228.580 ;
        RECT 745.525 228.340 745.785 228.600 ;
        RECT 2218.660 228.460 2218.920 228.720 ;
        RECT 742.280 227.760 742.540 228.020 ;
        RECT 746.495 227.780 746.755 228.040 ;
        RECT 2219.280 227.900 2219.540 228.160 ;
        RECT 747.640 227.480 747.900 227.740 ;
        RECT 751.505 227.500 751.765 227.760 ;
        RECT 2224.640 227.620 2224.900 227.880 ;
        RECT 748.260 226.920 748.520 227.180 ;
        RECT 752.475 226.940 752.735 227.200 ;
        RECT 2225.260 227.060 2225.520 227.320 ;
        RECT 753.620 226.640 753.880 226.900 ;
        RECT 757.485 226.660 757.745 226.920 ;
        RECT 2230.620 226.780 2230.880 227.040 ;
        RECT 754.240 226.080 754.500 226.340 ;
        RECT 758.455 226.100 758.715 226.360 ;
        RECT 2231.240 226.220 2231.500 226.480 ;
        RECT 759.600 225.800 759.860 226.060 ;
        RECT 763.465 225.820 763.725 226.080 ;
        RECT 2236.600 225.940 2236.860 226.200 ;
        RECT 764.435 225.260 764.695 225.520 ;
        RECT 2237.220 225.380 2237.480 225.640 ;
        RECT 769.445 224.980 769.705 225.240 ;
        RECT 2242.580 225.100 2242.840 225.360 ;
        RECT 770.415 224.420 770.675 224.680 ;
        RECT 2243.200 224.540 2243.460 224.800 ;
        RECT 775.425 224.140 775.685 224.400 ;
        RECT 2248.560 224.260 2248.820 224.520 ;
        RECT 776.275 223.580 776.535 223.840 ;
        RECT 2249.180 223.700 2249.440 223.960 ;
        RECT 781.405 223.300 781.665 223.560 ;
        RECT 2254.540 223.420 2254.800 223.680 ;
        RECT 782.375 222.740 782.635 223.000 ;
        RECT 2255.160 222.860 2255.420 223.120 ;
        RECT 787.385 222.460 787.645 222.720 ;
        RECT 2260.520 222.580 2260.780 222.840 ;
        RECT 788.235 221.900 788.495 222.160 ;
        RECT 2261.140 222.020 2261.400 222.280 ;
        RECT 793.365 221.340 793.625 221.600 ;
        RECT 2266.500 221.460 2266.760 221.720 ;
        RECT 794.335 220.780 794.595 221.040 ;
        RECT 2267.120 220.900 2267.380 221.160 ;
        RECT 670.470 215.510 670.730 216.360 ;
        RECT 674.240 215.810 675.330 216.070 ;
        RECT 676.450 215.510 676.710 216.360 ;
        RECT 680.220 215.810 681.310 216.070 ;
        RECT 682.430 215.510 682.690 216.360 ;
        RECT 686.200 215.810 687.290 216.070 ;
        RECT 688.410 215.510 688.670 216.360 ;
        RECT 692.180 215.810 693.270 216.070 ;
        RECT 694.390 215.510 694.650 216.360 ;
        RECT 698.160 215.810 699.250 216.070 ;
        RECT 700.370 215.510 700.630 216.360 ;
        RECT 704.140 215.810 705.230 216.070 ;
        RECT 706.350 215.510 706.610 216.360 ;
        RECT 710.120 215.810 711.210 216.070 ;
        RECT 712.330 215.510 712.590 216.360 ;
        RECT 716.100 215.810 717.190 216.070 ;
        RECT 718.310 215.510 718.570 216.360 ;
        RECT 722.080 215.810 723.170 216.070 ;
        RECT 724.290 215.510 724.550 216.360 ;
        RECT 728.060 215.810 729.150 216.070 ;
        RECT 730.270 215.510 730.530 216.360 ;
        RECT 734.040 215.810 735.130 216.070 ;
        RECT 736.250 215.510 736.510 216.360 ;
        RECT 740.020 215.810 741.110 216.070 ;
        RECT 742.230 215.510 742.490 216.360 ;
        RECT 746.000 215.810 747.090 216.070 ;
        RECT 748.210 215.510 748.470 216.360 ;
        RECT 751.980 215.810 753.070 216.070 ;
        RECT 754.190 215.510 754.450 216.360 ;
        RECT 757.960 215.810 759.050 216.070 ;
        RECT 763.940 215.810 765.030 216.070 ;
        RECT 769.920 215.810 771.010 216.070 ;
        RECT 775.900 215.810 776.990 216.070 ;
        RECT 781.880 215.810 782.970 216.070 ;
        RECT 787.860 215.810 788.950 216.070 ;
        RECT 793.840 215.810 794.930 216.070 ;
        RECT 2147.470 215.510 2147.730 216.360 ;
        RECT 2153.450 215.510 2153.710 216.360 ;
        RECT 2159.430 215.510 2159.690 216.360 ;
        RECT 2165.410 215.510 2165.670 216.360 ;
        RECT 2171.390 215.510 2171.650 216.360 ;
        RECT 2177.370 215.510 2177.630 216.360 ;
        RECT 2183.350 215.510 2183.610 216.360 ;
        RECT 2189.330 215.510 2189.590 216.360 ;
        RECT 2195.310 215.510 2195.570 216.360 ;
        RECT 2201.290 215.510 2201.550 216.360 ;
        RECT 2207.270 215.510 2207.530 216.360 ;
        RECT 2213.250 215.510 2213.510 216.360 ;
        RECT 2219.230 215.510 2219.490 216.360 ;
        RECT 2225.210 215.510 2225.470 216.360 ;
        RECT 2231.190 215.510 2231.450 216.360 ;
        RECT 2237.170 215.510 2237.430 216.360 ;
        RECT 2243.150 215.510 2243.410 216.360 ;
        RECT 2249.130 215.510 2249.390 216.360 ;
        RECT 2255.110 215.510 2255.370 216.360 ;
        RECT 2261.090 215.510 2261.350 216.360 ;
        RECT 2267.070 215.510 2267.330 216.360 ;
        RECT 675.590 212.750 676.680 213.010 ;
        RECT 679.680 212.450 679.940 213.300 ;
        RECT 681.570 212.750 682.660 213.010 ;
        RECT 685.660 212.450 685.920 213.300 ;
        RECT 687.550 212.750 688.640 213.010 ;
        RECT 691.640 212.450 691.900 213.300 ;
        RECT 693.530 212.750 694.620 213.010 ;
        RECT 697.620 212.450 697.880 213.300 ;
        RECT 699.510 212.750 700.600 213.010 ;
        RECT 703.600 212.450 703.860 213.300 ;
        RECT 705.490 212.750 706.580 213.010 ;
        RECT 709.580 212.450 709.840 213.300 ;
        RECT 711.470 212.750 712.560 213.010 ;
        RECT 715.560 212.450 715.820 213.300 ;
        RECT 717.450 212.750 718.540 213.010 ;
        RECT 721.540 212.450 721.800 213.300 ;
        RECT 723.430 212.750 724.520 213.010 ;
        RECT 727.520 212.450 727.780 213.300 ;
        RECT 729.410 212.750 730.500 213.010 ;
        RECT 733.500 212.450 733.760 213.300 ;
        RECT 735.390 212.750 736.480 213.010 ;
        RECT 739.480 212.450 739.740 213.300 ;
        RECT 741.370 212.750 742.460 213.010 ;
        RECT 745.460 212.450 745.720 213.300 ;
        RECT 747.350 212.750 748.440 213.010 ;
        RECT 751.440 212.450 751.700 213.300 ;
        RECT 753.330 212.750 754.420 213.010 ;
        RECT 757.420 212.450 757.680 213.300 ;
        RECT 759.310 212.750 760.400 213.010 ;
        RECT 763.400 212.450 763.660 213.300 ;
        RECT 769.380 212.450 769.640 213.300 ;
        RECT 775.360 212.450 775.620 213.300 ;
        RECT 781.340 212.450 781.600 213.300 ;
        RECT 787.320 212.450 787.580 213.300 ;
        RECT 793.340 212.750 794.430 213.010 ;
        RECT 2152.590 212.750 2153.680 213.010 ;
        RECT 2158.570 212.750 2159.660 213.010 ;
        RECT 2164.550 212.750 2165.640 213.010 ;
        RECT 2170.530 212.750 2171.620 213.010 ;
        RECT 2176.510 212.750 2177.600 213.010 ;
        RECT 2182.490 212.750 2183.580 213.010 ;
        RECT 2188.470 212.750 2189.560 213.010 ;
        RECT 2194.450 212.750 2195.540 213.010 ;
        RECT 2200.430 212.750 2201.520 213.010 ;
        RECT 2206.410 212.750 2207.500 213.010 ;
        RECT 2212.390 212.750 2213.480 213.010 ;
        RECT 2218.370 212.750 2219.460 213.010 ;
        RECT 2224.350 212.750 2225.440 213.010 ;
        RECT 2230.330 212.750 2231.420 213.010 ;
        RECT 2236.310 212.750 2237.400 213.010 ;
        RECT 2242.290 212.750 2243.380 213.010 ;
        RECT 2248.270 212.750 2249.360 213.010 ;
        RECT 2254.250 212.750 2255.340 213.010 ;
        RECT 2260.230 212.750 2261.320 213.010 ;
        RECT 2267.080 212.450 2267.340 213.300 ;
      LAYER met2 ;
        RECT 2087.570 4986.345 2088.660 4986.665 ;
        RECT 835.260 4984.720 836.350 4985.040 ;
        RECT 841.240 4984.720 842.330 4985.040 ;
        RECT 847.220 4984.720 848.310 4985.040 ;
        RECT 835.550 4974.795 835.690 4984.720 ;
        RECT 836.090 4981.400 836.410 4982.250 ;
        RECT 836.170 4975.075 836.310 4981.400 ;
        RECT 841.530 4975.915 841.670 4984.720 ;
        RECT 842.070 4981.400 842.390 4982.250 ;
        RECT 842.150 4976.195 842.290 4981.400 ;
        RECT 847.510 4977.035 847.650 4984.720 ;
        RECT 2087.510 4983.025 2087.830 4983.875 ;
        RECT 848.050 4981.400 848.370 4982.250 ;
        RECT 848.130 4977.315 848.270 4981.400 ;
        RECT 847.510 4976.715 847.770 4977.035 ;
        RECT 848.130 4976.995 848.390 4977.315 ;
        RECT 841.530 4975.595 841.790 4975.915 ;
        RECT 842.150 4975.875 842.410 4976.195 ;
        RECT 835.550 4974.475 835.810 4974.795 ;
        RECT 836.170 4974.755 836.430 4975.075 ;
        RECT 835.550 4974.400 835.690 4974.475 ;
        RECT 836.170 4974.400 836.310 4974.755 ;
        RECT 841.530 4974.400 841.670 4975.595 ;
        RECT 842.150 4974.400 842.290 4975.875 ;
        RECT 847.510 4975.275 847.650 4976.715 ;
        RECT 848.130 4975.275 848.270 4976.995 ;
        RECT 2087.610 4976.825 2087.750 4983.025 ;
        RECT 2087.490 4976.505 2087.750 4976.825 ;
        RECT 2088.230 4976.545 2088.370 4986.345 ;
        RECT 3311.285 4985.675 3311.605 4986.525 ;
        RECT 3314.575 4985.935 3315.665 4986.255 ;
        RECT 3320.555 4985.935 3321.645 4986.255 ;
        RECT 3326.535 4985.935 3327.625 4986.255 ;
        RECT 3332.515 4985.935 3333.605 4986.255 ;
        RECT 3309.945 4982.875 3311.035 4983.195 ;
        RECT 3310.400 4976.945 3310.540 4982.875 ;
        RECT 3310.280 4976.625 3310.540 4976.945 ;
        RECT 3311.370 4976.665 3311.510 4985.675 ;
        RECT 3314.515 4982.615 3314.835 4983.465 ;
        RECT 3314.615 4976.965 3314.755 4982.615 ;
        RECT 2087.610 4976.430 2087.750 4976.505 ;
        RECT 2088.110 4976.225 2088.370 4976.545 ;
        RECT 2088.230 4976.065 2088.370 4976.225 ;
        RECT 3310.400 4972.845 3310.540 4976.625 ;
        RECT 3311.250 4976.345 3311.510 4976.665 ;
        RECT 3314.495 4976.645 3314.755 4976.965 ;
        RECT 3315.235 4976.685 3315.375 4985.935 ;
        RECT 3320.495 4982.615 3320.815 4983.465 ;
        RECT 3311.370 4972.845 3311.510 4976.345 ;
        RECT 3314.615 4972.845 3314.755 4976.645 ;
        RECT 3315.115 4976.365 3315.375 4976.685 ;
        RECT 3315.235 4972.845 3315.375 4976.365 ;
        RECT 3320.595 4975.845 3320.735 4982.615 ;
        RECT 3320.475 4975.525 3320.735 4975.845 ;
        RECT 3321.215 4975.565 3321.355 4985.935 ;
        RECT 3326.475 4982.615 3326.795 4983.465 ;
        RECT 3320.595 4972.845 3320.735 4975.525 ;
        RECT 3321.095 4975.245 3321.355 4975.565 ;
        RECT 3321.215 4972.845 3321.355 4975.245 ;
        RECT 3326.575 4974.725 3326.715 4982.615 ;
        RECT 3326.455 4974.405 3326.715 4974.725 ;
        RECT 3327.195 4974.445 3327.335 4985.935 ;
        RECT 3332.455 4982.615 3332.775 4983.465 ;
        RECT 3326.575 4972.845 3326.715 4974.405 ;
        RECT 3327.075 4974.125 3327.335 4974.445 ;
        RECT 3327.195 4972.845 3327.335 4974.125 ;
        RECT 3332.555 4973.605 3332.695 4982.615 ;
        RECT 3332.435 4973.285 3332.695 4973.605 ;
        RECT 3333.175 4973.325 3333.315 4985.935 ;
        RECT 3332.555 4972.845 3332.695 4973.285 ;
        RECT 3333.055 4973.005 3333.315 4973.325 ;
        RECT 3333.175 4972.845 3333.315 4973.005 ;
        RECT 205.940 4456.635 206.260 4457.090 ;
        RECT 211.025 4456.635 211.345 4456.755 ;
        RECT 205.940 4456.495 216.135 4456.635 ;
        RECT 205.940 4456.000 206.260 4456.495 ;
        RECT 202.610 4455.665 203.460 4455.750 ;
        RECT 211.305 4455.665 211.625 4455.785 ;
        RECT 202.610 4455.525 216.135 4455.665 ;
        RECT 202.610 4455.430 203.460 4455.525 ;
        RECT 202.880 4451.800 203.200 4452.460 ;
        RECT 205.670 4452.420 206.520 4452.520 ;
        RECT 211.005 4452.420 211.325 4452.540 ;
        RECT 205.670 4452.280 216.135 4452.420 ;
        RECT 205.670 4452.200 206.520 4452.280 ;
        RECT 211.285 4451.800 211.605 4451.920 ;
        RECT 202.880 4451.660 216.135 4451.800 ;
        RECT 202.880 4451.370 203.200 4451.660 ;
        RECT 205.940 4450.655 206.260 4451.110 ;
        RECT 205.940 4450.515 216.135 4450.655 ;
        RECT 205.940 4450.020 206.260 4450.515 ;
        RECT 212.145 4450.395 212.465 4450.515 ;
        RECT 202.610 4449.685 203.460 4449.770 ;
        RECT 212.425 4449.685 212.745 4449.805 ;
        RECT 202.610 4449.545 216.135 4449.685 ;
        RECT 202.610 4449.450 203.460 4449.545 ;
        RECT 202.880 4445.820 203.200 4446.480 ;
        RECT 205.670 4446.440 206.520 4446.540 ;
        RECT 212.125 4446.440 212.445 4446.560 ;
        RECT 205.670 4446.300 216.135 4446.440 ;
        RECT 205.670 4446.220 206.520 4446.300 ;
        RECT 212.405 4445.820 212.725 4445.940 ;
        RECT 202.880 4445.680 216.135 4445.820 ;
        RECT 202.880 4445.390 203.200 4445.680 ;
        RECT 205.940 4444.675 206.260 4445.130 ;
        RECT 213.265 4444.675 213.585 4444.795 ;
        RECT 205.940 4444.535 216.135 4444.675 ;
        RECT 205.940 4444.040 206.260 4444.535 ;
        RECT 202.610 4443.705 203.460 4443.790 ;
        RECT 213.545 4443.705 213.865 4443.825 ;
        RECT 202.610 4443.565 216.135 4443.705 ;
        RECT 202.610 4443.470 203.460 4443.565 ;
        RECT 202.880 4439.840 203.200 4440.500 ;
        RECT 205.670 4440.460 206.520 4440.560 ;
        RECT 213.245 4440.460 213.565 4440.580 ;
        RECT 205.670 4440.320 216.135 4440.460 ;
        RECT 205.670 4440.240 206.520 4440.320 ;
        RECT 213.525 4439.840 213.845 4439.960 ;
        RECT 202.880 4439.700 216.135 4439.840 ;
        RECT 202.880 4439.410 203.200 4439.700 ;
        RECT 202.880 4433.860 203.200 4434.520 ;
        RECT 205.670 4434.480 206.520 4434.580 ;
        RECT 214.365 4434.480 214.685 4434.600 ;
        RECT 205.670 4434.340 216.135 4434.480 ;
        RECT 205.670 4434.260 206.520 4434.340 ;
        RECT 214.645 4433.860 214.965 4433.980 ;
        RECT 202.880 4433.720 216.135 4433.860 ;
        RECT 202.880 4433.430 203.200 4433.720 ;
        RECT 202.880 4427.880 203.200 4428.540 ;
        RECT 205.670 4428.500 206.520 4428.600 ;
        RECT 215.485 4428.500 215.805 4428.620 ;
        RECT 205.670 4428.360 216.135 4428.500 ;
        RECT 205.670 4428.280 206.520 4428.360 ;
        RECT 215.765 4427.880 216.085 4428.000 ;
        RECT 202.880 4427.740 216.135 4427.880 ;
        RECT 202.880 4427.450 203.200 4427.740 ;
        RECT 3381.610 3637.835 3381.930 3638.290 ;
        RECT 3376.150 3637.695 3381.930 3637.835 ;
        RECT 3376.490 3637.575 3376.810 3637.695 ;
        RECT 3381.610 3637.200 3381.930 3637.695 ;
        RECT 3376.210 3636.865 3376.530 3636.985 ;
        RECT 3384.410 3636.865 3385.260 3636.950 ;
        RECT 3376.150 3636.725 3385.260 3636.865 ;
        RECT 3384.410 3636.630 3385.260 3636.725 ;
        RECT 3376.510 3633.620 3376.830 3633.740 ;
        RECT 3381.350 3633.620 3382.200 3633.720 ;
        RECT 3376.265 3633.480 3382.200 3633.620 ;
        RECT 3381.350 3633.400 3382.200 3633.480 ;
        RECT 3376.230 3633.000 3376.550 3633.120 ;
        RECT 3384.670 3633.000 3384.990 3633.660 ;
        RECT 3376.230 3632.860 3384.990 3633.000 ;
        RECT 3384.670 3632.570 3384.990 3632.860 ;
        RECT 3375.230 3631.855 3375.550 3631.975 ;
        RECT 3381.610 3631.855 3381.930 3632.310 ;
        RECT 3369.210 3631.715 3381.930 3631.855 ;
        RECT 3381.610 3631.220 3381.930 3631.715 ;
        RECT 3374.950 3630.885 3375.270 3631.005 ;
        RECT 3384.410 3630.885 3385.260 3630.970 ;
        RECT 3369.210 3630.745 3385.260 3630.885 ;
        RECT 3384.410 3630.650 3385.260 3630.745 ;
        RECT 3375.250 3627.640 3375.570 3627.760 ;
        RECT 3381.350 3627.640 3382.200 3627.740 ;
        RECT 3369.210 3627.500 3382.200 3627.640 ;
        RECT 3381.350 3627.420 3382.200 3627.500 ;
        RECT 3374.970 3627.020 3375.290 3627.140 ;
        RECT 3384.670 3627.020 3384.990 3627.680 ;
        RECT 3369.210 3626.880 3384.990 3627.020 ;
        RECT 3384.670 3626.590 3384.990 3626.880 ;
        RECT 3374.110 3625.875 3374.430 3625.995 ;
        RECT 3381.610 3625.875 3381.930 3626.330 ;
        RECT 3369.210 3625.735 3381.930 3625.875 ;
        RECT 3381.610 3625.240 3381.930 3625.735 ;
        RECT 3373.830 3624.905 3374.150 3625.025 ;
        RECT 3384.410 3624.905 3385.260 3624.990 ;
        RECT 3369.210 3624.765 3385.260 3624.905 ;
        RECT 3384.410 3624.670 3385.260 3624.765 ;
        RECT 3374.130 3621.660 3374.450 3621.780 ;
        RECT 3381.350 3621.660 3382.200 3621.760 ;
        RECT 3369.210 3621.520 3382.200 3621.660 ;
        RECT 3381.350 3621.440 3382.200 3621.520 ;
        RECT 3373.850 3621.040 3374.170 3621.160 ;
        RECT 3384.670 3621.040 3384.990 3621.700 ;
        RECT 3369.210 3620.900 3384.990 3621.040 ;
        RECT 3384.670 3620.610 3384.990 3620.900 ;
        RECT 3372.990 3619.895 3373.310 3620.015 ;
        RECT 3381.610 3619.895 3381.930 3620.350 ;
        RECT 3369.210 3619.755 3381.930 3619.895 ;
        RECT 3381.610 3619.260 3381.930 3619.755 ;
        RECT 3372.710 3618.925 3373.030 3619.045 ;
        RECT 3384.410 3618.925 3385.260 3619.010 ;
        RECT 3369.210 3618.785 3385.260 3618.925 ;
        RECT 3384.410 3618.690 3385.260 3618.785 ;
        RECT 3373.010 3615.680 3373.330 3615.800 ;
        RECT 3381.350 3615.680 3382.200 3615.780 ;
        RECT 3369.210 3615.540 3382.200 3615.680 ;
        RECT 3381.350 3615.460 3382.200 3615.540 ;
        RECT 3372.730 3615.060 3373.050 3615.180 ;
        RECT 3384.670 3615.060 3384.990 3615.720 ;
        RECT 3369.210 3614.920 3384.990 3615.060 ;
        RECT 3384.670 3614.630 3384.990 3614.920 ;
        RECT 3371.890 3609.700 3372.210 3609.820 ;
        RECT 3381.350 3609.700 3382.200 3609.800 ;
        RECT 3369.210 3609.560 3382.200 3609.700 ;
        RECT 3381.350 3609.480 3382.200 3609.560 ;
        RECT 3371.610 3609.080 3371.930 3609.200 ;
        RECT 3384.670 3609.080 3384.990 3609.740 ;
        RECT 3369.210 3608.940 3384.990 3609.080 ;
        RECT 3384.670 3608.650 3384.990 3608.940 ;
        RECT 3370.770 3603.720 3371.090 3603.840 ;
        RECT 3381.350 3603.720 3382.200 3603.820 ;
        RECT 3370.330 3603.580 3382.200 3603.720 ;
        RECT 3381.350 3603.500 3382.200 3603.580 ;
        RECT 3370.490 3603.100 3370.810 3603.220 ;
        RECT 3384.670 3603.100 3384.990 3603.760 ;
        RECT 3370.330 3602.960 3384.990 3603.100 ;
        RECT 3384.670 3602.670 3384.990 3602.960 ;
        RECT 206.065 3050.405 206.385 3050.860 ;
        RECT 210.885 3050.405 211.205 3050.525 ;
        RECT 206.065 3050.265 221.600 3050.405 ;
        RECT 206.065 3049.770 206.385 3050.265 ;
        RECT 202.735 3049.435 203.585 3049.520 ;
        RECT 211.165 3049.435 211.485 3049.555 ;
        RECT 202.735 3049.295 221.600 3049.435 ;
        RECT 202.735 3049.200 203.585 3049.295 ;
        RECT 203.005 3045.570 203.325 3046.230 ;
        RECT 205.795 3046.190 206.645 3046.290 ;
        RECT 210.865 3046.190 211.185 3046.310 ;
        RECT 205.795 3046.050 221.600 3046.190 ;
        RECT 205.795 3045.970 206.645 3046.050 ;
        RECT 211.145 3045.570 211.465 3045.690 ;
        RECT 203.005 3045.430 221.600 3045.570 ;
        RECT 203.005 3045.140 203.325 3045.430 ;
        RECT 206.065 3044.425 206.385 3044.880 ;
        RECT 206.065 3044.285 221.600 3044.425 ;
        RECT 206.065 3043.790 206.385 3044.285 ;
        RECT 212.005 3044.165 212.325 3044.285 ;
        RECT 202.735 3043.455 203.585 3043.540 ;
        RECT 212.285 3043.455 212.605 3043.575 ;
        RECT 202.735 3043.315 221.600 3043.455 ;
        RECT 202.735 3043.220 203.585 3043.315 ;
        RECT 203.005 3039.590 203.325 3040.250 ;
        RECT 205.795 3040.210 206.645 3040.310 ;
        RECT 211.985 3040.210 212.305 3040.330 ;
        RECT 205.795 3040.070 221.600 3040.210 ;
        RECT 205.795 3039.990 206.645 3040.070 ;
        RECT 212.265 3039.590 212.585 3039.710 ;
        RECT 203.005 3039.450 221.600 3039.590 ;
        RECT 203.005 3039.160 203.325 3039.450 ;
        RECT 206.065 3038.445 206.385 3038.900 ;
        RECT 213.125 3038.445 213.445 3038.565 ;
        RECT 206.065 3038.305 221.600 3038.445 ;
        RECT 206.065 3037.810 206.385 3038.305 ;
        RECT 202.735 3037.475 203.585 3037.560 ;
        RECT 213.405 3037.475 213.725 3037.595 ;
        RECT 202.735 3037.335 221.600 3037.475 ;
        RECT 202.735 3037.240 203.585 3037.335 ;
        RECT 203.005 3033.610 203.325 3034.270 ;
        RECT 205.795 3034.230 206.645 3034.330 ;
        RECT 213.105 3034.230 213.425 3034.350 ;
        RECT 205.795 3034.090 221.600 3034.230 ;
        RECT 205.795 3034.010 206.645 3034.090 ;
        RECT 213.385 3033.610 213.705 3033.730 ;
        RECT 203.005 3033.470 221.600 3033.610 ;
        RECT 203.005 3033.180 203.325 3033.470 ;
        RECT 206.065 3032.465 206.385 3032.920 ;
        RECT 206.065 3032.325 221.600 3032.465 ;
        RECT 206.065 3031.830 206.385 3032.325 ;
        RECT 214.245 3032.205 214.565 3032.325 ;
        RECT 202.735 3031.495 203.585 3031.580 ;
        RECT 214.525 3031.495 214.845 3031.615 ;
        RECT 202.735 3031.355 221.600 3031.495 ;
        RECT 202.735 3031.260 203.585 3031.355 ;
        RECT 203.005 3027.630 203.325 3028.290 ;
        RECT 205.795 3028.250 206.645 3028.350 ;
        RECT 214.225 3028.250 214.545 3028.370 ;
        RECT 205.795 3028.110 221.600 3028.250 ;
        RECT 205.795 3028.030 206.645 3028.110 ;
        RECT 214.505 3027.630 214.825 3027.750 ;
        RECT 203.005 3027.490 221.600 3027.630 ;
        RECT 203.005 3027.200 203.325 3027.490 ;
        RECT 206.065 3026.485 206.385 3026.940 ;
        RECT 215.365 3026.485 215.685 3026.605 ;
        RECT 206.065 3026.345 221.600 3026.485 ;
        RECT 206.065 3025.850 206.385 3026.345 ;
        RECT 202.735 3025.515 203.585 3025.600 ;
        RECT 215.645 3025.515 215.965 3025.635 ;
        RECT 202.735 3025.375 221.600 3025.515 ;
        RECT 202.735 3025.280 203.585 3025.375 ;
        RECT 203.005 3021.650 203.325 3022.310 ;
        RECT 205.795 3022.270 206.645 3022.370 ;
        RECT 215.345 3022.270 215.665 3022.390 ;
        RECT 205.795 3022.130 221.600 3022.270 ;
        RECT 205.795 3022.050 206.645 3022.130 ;
        RECT 215.625 3021.650 215.945 3021.770 ;
        RECT 203.005 3021.510 221.600 3021.650 ;
        RECT 203.005 3021.220 203.325 3021.510 ;
        RECT 203.005 3015.670 203.325 3016.330 ;
        RECT 205.795 3016.290 206.645 3016.390 ;
        RECT 216.465 3016.290 216.785 3016.410 ;
        RECT 205.795 3016.150 221.600 3016.290 ;
        RECT 205.795 3016.070 206.645 3016.150 ;
        RECT 216.745 3015.670 217.065 3015.790 ;
        RECT 203.005 3015.530 221.600 3015.670 ;
        RECT 203.005 3015.240 203.325 3015.530 ;
        RECT 203.005 3009.690 203.325 3010.350 ;
        RECT 205.795 3010.310 206.645 3010.410 ;
        RECT 217.585 3010.310 217.905 3010.430 ;
        RECT 205.795 3010.170 221.600 3010.310 ;
        RECT 205.795 3010.090 206.645 3010.170 ;
        RECT 217.865 3009.690 218.185 3009.810 ;
        RECT 203.005 3009.550 221.600 3009.690 ;
        RECT 203.005 3009.260 203.325 3009.550 ;
        RECT 203.005 3003.710 203.325 3004.370 ;
        RECT 205.795 3004.330 206.645 3004.430 ;
        RECT 218.705 3004.330 219.025 3004.450 ;
        RECT 205.795 3004.190 221.600 3004.330 ;
        RECT 205.795 3004.110 206.645 3004.190 ;
        RECT 218.985 3003.710 219.305 3003.830 ;
        RECT 203.005 3003.570 221.600 3003.710 ;
        RECT 203.005 3003.280 203.325 3003.570 ;
        RECT 203.005 2997.730 203.325 2998.390 ;
        RECT 205.795 2998.350 206.645 2998.450 ;
        RECT 219.825 2998.350 220.145 2998.470 ;
        RECT 205.795 2998.210 221.600 2998.350 ;
        RECT 205.795 2998.130 206.645 2998.210 ;
        RECT 220.105 2997.730 220.425 2997.850 ;
        RECT 203.005 2997.590 221.600 2997.730 ;
        RECT 203.005 2997.300 203.325 2997.590 ;
        RECT 203.005 2991.750 203.325 2992.410 ;
        RECT 205.795 2992.370 206.645 2992.470 ;
        RECT 220.945 2992.370 221.265 2992.490 ;
        RECT 205.795 2992.230 221.675 2992.370 ;
        RECT 205.795 2992.150 206.645 2992.230 ;
        RECT 221.225 2991.750 221.545 2991.870 ;
        RECT 203.005 2991.610 221.675 2991.750 ;
        RECT 203.005 2991.320 203.325 2991.610 ;
        RECT 203.005 2985.770 203.325 2986.430 ;
        RECT 205.795 2986.390 206.645 2986.490 ;
        RECT 222.065 2986.390 222.385 2986.510 ;
        RECT 205.795 2986.250 222.720 2986.390 ;
        RECT 205.795 2986.170 206.645 2986.250 ;
        RECT 222.345 2985.770 222.665 2985.890 ;
        RECT 203.005 2985.630 222.720 2985.770 ;
        RECT 203.005 2985.340 203.325 2985.630 ;
        RECT 3376.630 2267.715 3376.950 2267.835 ;
        RECT 3381.610 2267.715 3381.930 2268.170 ;
        RECT 3365.990 2267.575 3381.930 2267.715 ;
        RECT 3381.610 2267.080 3381.930 2267.575 ;
        RECT 3376.350 2266.745 3376.670 2266.865 ;
        RECT 3384.410 2266.745 3385.260 2266.830 ;
        RECT 3365.990 2266.605 3385.260 2266.745 ;
        RECT 3384.410 2266.510 3385.260 2266.605 ;
        RECT 3365.990 2262.740 3375.745 2262.880 ;
        RECT 3381.610 2261.735 3381.930 2262.190 ;
        RECT 3365.990 2261.595 3381.930 2261.735 ;
        RECT 3375.370 2261.475 3375.690 2261.595 ;
        RECT 3381.610 2261.100 3381.930 2261.595 ;
        RECT 3375.090 2260.765 3375.410 2260.885 ;
        RECT 3384.410 2260.765 3385.260 2260.850 ;
        RECT 3365.990 2260.625 3385.260 2260.765 ;
        RECT 3384.410 2260.530 3385.260 2260.625 ;
        RECT 3374.250 2255.755 3374.570 2255.875 ;
        RECT 3381.610 2255.755 3381.930 2256.210 ;
        RECT 3365.990 2255.615 3381.930 2255.755 ;
        RECT 3381.610 2255.120 3381.930 2255.615 ;
        RECT 3373.970 2254.785 3374.290 2254.905 ;
        RECT 3384.410 2254.785 3385.260 2254.870 ;
        RECT 3365.990 2254.645 3385.260 2254.785 ;
        RECT 3384.410 2254.550 3385.260 2254.645 ;
        RECT 3381.610 2249.775 3381.930 2250.230 ;
        RECT 3365.990 2249.635 3381.930 2249.775 ;
        RECT 3373.130 2249.515 3373.450 2249.635 ;
        RECT 3381.610 2249.140 3381.930 2249.635 ;
        RECT 3372.850 2248.805 3373.170 2248.925 ;
        RECT 3384.410 2248.805 3385.260 2248.890 ;
        RECT 3365.990 2248.665 3385.260 2248.805 ;
        RECT 3384.410 2248.570 3385.260 2248.665 ;
        RECT 3372.010 2243.795 3372.330 2243.915 ;
        RECT 3381.610 2243.795 3381.930 2244.250 ;
        RECT 3365.990 2243.655 3381.930 2243.795 ;
        RECT 3381.610 2243.160 3381.930 2243.655 ;
        RECT 3371.730 2242.825 3372.050 2242.945 ;
        RECT 3384.410 2242.825 3385.260 2242.910 ;
        RECT 3365.990 2242.685 3385.260 2242.825 ;
        RECT 3384.410 2242.590 3385.260 2242.685 ;
        RECT 3370.890 2237.815 3371.210 2237.935 ;
        RECT 3381.610 2237.815 3381.930 2238.270 ;
        RECT 3365.990 2237.675 3381.930 2237.815 ;
        RECT 3381.610 2237.180 3381.930 2237.675 ;
        RECT 3370.610 2236.845 3370.930 2236.965 ;
        RECT 3384.410 2236.845 3385.260 2236.930 ;
        RECT 3365.990 2236.705 3385.260 2236.845 ;
        RECT 3384.410 2236.610 3385.260 2236.705 ;
        RECT 206.175 1762.500 206.495 1762.955 ;
        RECT 210.745 1762.500 211.065 1762.620 ;
        RECT 206.175 1762.360 223.740 1762.500 ;
        RECT 206.175 1761.865 206.495 1762.360 ;
        RECT 202.845 1761.530 203.695 1761.615 ;
        RECT 211.025 1761.530 211.345 1761.650 ;
        RECT 202.845 1761.390 223.740 1761.530 ;
        RECT 202.845 1761.295 203.695 1761.390 ;
        RECT 203.115 1757.665 203.435 1758.325 ;
        RECT 205.905 1758.285 206.755 1758.385 ;
        RECT 210.725 1758.285 211.045 1758.405 ;
        RECT 205.905 1758.145 223.740 1758.285 ;
        RECT 205.905 1758.065 206.755 1758.145 ;
        RECT 211.005 1757.665 211.330 1757.785 ;
        RECT 203.115 1757.525 223.740 1757.665 ;
        RECT 203.115 1757.235 203.435 1757.525 ;
        RECT 206.175 1756.520 206.495 1756.975 ;
        RECT 206.175 1756.380 223.740 1756.520 ;
        RECT 206.175 1755.885 206.495 1756.380 ;
        RECT 211.865 1756.260 212.185 1756.380 ;
        RECT 202.845 1755.550 203.695 1755.635 ;
        RECT 212.145 1755.550 212.465 1755.670 ;
        RECT 202.845 1755.410 223.740 1755.550 ;
        RECT 202.845 1755.315 203.695 1755.410 ;
        RECT 203.115 1751.685 203.435 1752.345 ;
        RECT 205.855 1752.305 206.705 1752.405 ;
        RECT 211.845 1752.305 212.165 1752.425 ;
        RECT 205.855 1752.165 223.740 1752.305 ;
        RECT 205.855 1752.085 206.705 1752.165 ;
        RECT 212.125 1751.685 212.445 1751.805 ;
        RECT 203.115 1751.545 223.740 1751.685 ;
        RECT 203.115 1751.255 203.435 1751.545 ;
        RECT 206.175 1750.540 206.495 1750.995 ;
        RECT 212.985 1750.540 213.305 1750.660 ;
        RECT 206.175 1750.400 223.740 1750.540 ;
        RECT 206.175 1749.905 206.495 1750.400 ;
        RECT 202.845 1749.570 203.695 1749.655 ;
        RECT 213.265 1749.570 213.585 1749.690 ;
        RECT 202.845 1749.430 223.740 1749.570 ;
        RECT 202.845 1749.335 203.695 1749.430 ;
        RECT 203.115 1745.705 203.435 1746.365 ;
        RECT 205.905 1746.325 206.755 1746.425 ;
        RECT 212.965 1746.325 213.285 1746.445 ;
        RECT 205.905 1746.185 223.740 1746.325 ;
        RECT 205.905 1746.105 206.755 1746.185 ;
        RECT 213.245 1745.705 213.565 1745.825 ;
        RECT 203.115 1745.565 223.740 1745.705 ;
        RECT 203.115 1745.275 203.435 1745.565 ;
        RECT 206.175 1744.560 206.495 1745.015 ;
        RECT 206.175 1744.420 223.740 1744.560 ;
        RECT 206.175 1743.925 206.495 1744.420 ;
        RECT 214.105 1744.300 214.425 1744.420 ;
        RECT 202.845 1743.590 203.695 1743.675 ;
        RECT 214.385 1743.590 214.705 1743.710 ;
        RECT 202.845 1743.450 223.740 1743.590 ;
        RECT 202.845 1743.355 203.695 1743.450 ;
        RECT 203.115 1739.725 203.435 1740.385 ;
        RECT 205.905 1740.345 206.755 1740.445 ;
        RECT 214.085 1740.345 214.405 1740.465 ;
        RECT 205.905 1740.205 223.740 1740.345 ;
        RECT 205.905 1740.125 206.755 1740.205 ;
        RECT 214.365 1739.725 214.685 1739.845 ;
        RECT 203.115 1739.585 223.740 1739.725 ;
        RECT 203.115 1739.295 203.435 1739.585 ;
        RECT 206.175 1738.580 206.495 1739.035 ;
        RECT 215.225 1738.580 215.545 1738.700 ;
        RECT 206.175 1738.440 223.740 1738.580 ;
        RECT 206.175 1737.945 206.495 1738.440 ;
        RECT 202.845 1737.610 203.695 1737.695 ;
        RECT 215.505 1737.610 215.825 1737.730 ;
        RECT 202.845 1737.470 223.740 1737.610 ;
        RECT 202.845 1737.375 203.695 1737.470 ;
        RECT 203.115 1733.745 203.435 1734.405 ;
        RECT 205.905 1734.365 206.755 1734.465 ;
        RECT 215.205 1734.365 215.525 1734.485 ;
        RECT 205.905 1734.225 223.740 1734.365 ;
        RECT 205.905 1734.145 206.755 1734.225 ;
        RECT 215.485 1733.745 215.805 1733.865 ;
        RECT 203.115 1733.605 223.740 1733.745 ;
        RECT 203.115 1733.315 203.435 1733.605 ;
        RECT 206.175 1732.600 206.495 1733.055 ;
        RECT 216.345 1732.600 216.665 1732.720 ;
        RECT 206.175 1732.460 223.740 1732.600 ;
        RECT 206.175 1731.965 206.495 1732.460 ;
        RECT 202.845 1731.630 203.695 1731.715 ;
        RECT 216.625 1731.630 216.945 1731.750 ;
        RECT 202.845 1731.490 223.740 1731.630 ;
        RECT 202.845 1731.395 203.695 1731.490 ;
        RECT 203.115 1727.765 203.435 1728.425 ;
        RECT 205.905 1728.385 206.755 1728.485 ;
        RECT 216.325 1728.385 216.645 1728.505 ;
        RECT 205.905 1728.245 223.740 1728.385 ;
        RECT 205.905 1728.165 206.755 1728.245 ;
        RECT 216.605 1727.765 216.925 1727.885 ;
        RECT 203.115 1727.625 223.740 1727.765 ;
        RECT 203.115 1727.335 203.435 1727.625 ;
        RECT 206.175 1726.620 206.495 1727.075 ;
        RECT 217.465 1726.620 217.785 1726.740 ;
        RECT 206.175 1726.480 223.740 1726.620 ;
        RECT 206.175 1725.985 206.495 1726.480 ;
        RECT 202.845 1725.650 203.695 1725.735 ;
        RECT 217.745 1725.650 218.065 1725.770 ;
        RECT 202.845 1725.510 223.740 1725.650 ;
        RECT 202.845 1725.415 203.695 1725.510 ;
        RECT 203.115 1721.785 203.435 1722.445 ;
        RECT 205.905 1722.405 206.755 1722.505 ;
        RECT 217.445 1722.405 217.765 1722.525 ;
        RECT 205.905 1722.265 223.740 1722.405 ;
        RECT 205.905 1722.185 206.755 1722.265 ;
        RECT 217.725 1721.785 218.045 1721.905 ;
        RECT 203.115 1721.645 223.740 1721.785 ;
        RECT 203.115 1721.355 203.435 1721.645 ;
        RECT 206.175 1720.640 206.495 1721.095 ;
        RECT 218.585 1720.640 218.905 1720.760 ;
        RECT 206.175 1720.500 223.740 1720.640 ;
        RECT 206.175 1720.005 206.495 1720.500 ;
        RECT 202.845 1719.670 203.695 1719.755 ;
        RECT 218.865 1719.670 219.185 1719.790 ;
        RECT 202.845 1719.530 223.740 1719.670 ;
        RECT 202.845 1719.435 203.695 1719.530 ;
        RECT 203.115 1715.805 203.435 1716.465 ;
        RECT 205.905 1716.425 206.755 1716.525 ;
        RECT 218.565 1716.425 218.885 1716.545 ;
        RECT 205.905 1716.285 223.740 1716.425 ;
        RECT 205.905 1716.205 206.755 1716.285 ;
        RECT 218.845 1715.805 219.165 1715.925 ;
        RECT 202.845 1715.665 223.740 1715.805 ;
        RECT 203.115 1715.375 203.435 1715.665 ;
        RECT 206.175 1714.660 206.495 1715.115 ;
        RECT 219.705 1714.660 220.025 1714.780 ;
        RECT 206.175 1714.520 223.740 1714.660 ;
        RECT 206.175 1714.025 206.495 1714.520 ;
        RECT 202.845 1713.690 203.695 1713.775 ;
        RECT 219.985 1713.690 220.305 1713.810 ;
        RECT 202.845 1713.550 223.740 1713.690 ;
        RECT 202.845 1713.455 203.695 1713.550 ;
        RECT 203.115 1709.825 203.435 1710.485 ;
        RECT 205.905 1710.445 206.755 1710.545 ;
        RECT 219.685 1710.445 220.005 1710.565 ;
        RECT 205.905 1710.305 223.740 1710.445 ;
        RECT 205.905 1710.225 206.755 1710.305 ;
        RECT 219.965 1709.825 220.285 1709.945 ;
        RECT 203.115 1709.685 223.740 1709.825 ;
        RECT 203.115 1709.395 203.435 1709.685 ;
        RECT 206.175 1708.680 206.495 1709.135 ;
        RECT 220.825 1708.680 221.145 1708.800 ;
        RECT 206.175 1708.540 223.740 1708.680 ;
        RECT 206.175 1708.045 206.495 1708.540 ;
        RECT 202.845 1707.710 203.695 1707.795 ;
        RECT 221.105 1707.710 221.425 1707.830 ;
        RECT 202.845 1707.570 223.740 1707.710 ;
        RECT 202.845 1707.475 203.695 1707.570 ;
        RECT 203.115 1703.845 203.435 1704.505 ;
        RECT 205.905 1704.465 206.755 1704.565 ;
        RECT 220.805 1704.465 221.125 1704.585 ;
        RECT 205.905 1704.325 223.740 1704.465 ;
        RECT 205.905 1704.245 206.755 1704.325 ;
        RECT 221.085 1703.845 221.405 1703.965 ;
        RECT 203.115 1703.705 223.740 1703.845 ;
        RECT 203.115 1703.415 203.435 1703.705 ;
        RECT 206.175 1702.700 206.495 1703.155 ;
        RECT 221.945 1702.700 222.265 1702.820 ;
        RECT 206.175 1702.560 223.740 1702.700 ;
        RECT 206.175 1702.065 206.495 1702.560 ;
        RECT 202.845 1701.730 203.695 1701.815 ;
        RECT 222.225 1701.730 222.545 1701.850 ;
        RECT 202.845 1701.590 223.740 1701.730 ;
        RECT 202.845 1701.495 203.695 1701.590 ;
        RECT 203.115 1697.865 203.435 1698.525 ;
        RECT 205.905 1698.485 206.755 1698.585 ;
        RECT 221.925 1698.485 222.245 1698.605 ;
        RECT 205.905 1698.345 223.740 1698.485 ;
        RECT 205.905 1698.265 206.755 1698.345 ;
        RECT 222.205 1697.865 222.525 1697.985 ;
        RECT 203.115 1697.725 223.740 1697.865 ;
        RECT 203.115 1697.435 203.435 1697.725 ;
        RECT 203.115 1691.885 203.435 1692.545 ;
        RECT 205.905 1692.505 206.755 1692.605 ;
        RECT 223.045 1692.505 223.365 1692.625 ;
        RECT 205.905 1692.365 223.745 1692.505 ;
        RECT 205.905 1692.285 206.755 1692.365 ;
        RECT 223.325 1691.885 223.645 1692.005 ;
        RECT 203.115 1691.745 223.745 1691.885 ;
        RECT 203.115 1691.455 203.435 1691.745 ;
        RECT 203.115 1685.905 203.435 1686.565 ;
        RECT 205.905 1686.525 206.755 1686.625 ;
        RECT 224.165 1686.525 224.485 1686.645 ;
        RECT 205.905 1686.385 224.805 1686.525 ;
        RECT 205.905 1686.305 206.755 1686.385 ;
        RECT 224.445 1685.905 224.765 1686.025 ;
        RECT 203.115 1685.765 224.805 1685.905 ;
        RECT 203.115 1685.475 203.435 1685.765 ;
        RECT 203.115 1679.925 203.435 1680.585 ;
        RECT 205.905 1680.545 206.755 1680.645 ;
        RECT 225.285 1680.545 225.605 1680.665 ;
        RECT 205.905 1680.405 226.030 1680.545 ;
        RECT 205.905 1680.325 206.755 1680.405 ;
        RECT 225.565 1679.925 225.885 1680.045 ;
        RECT 203.115 1679.785 226.030 1679.925 ;
        RECT 203.115 1679.495 203.435 1679.785 ;
        RECT 203.115 1673.945 203.435 1674.605 ;
        RECT 205.905 1674.565 206.755 1674.665 ;
        RECT 226.405 1674.565 226.725 1674.685 ;
        RECT 205.905 1674.425 227.100 1674.565 ;
        RECT 205.905 1674.345 206.755 1674.425 ;
        RECT 226.685 1673.945 227.005 1674.065 ;
        RECT 203.115 1673.805 227.100 1673.945 ;
        RECT 203.115 1673.515 203.435 1673.805 ;
        RECT 2147.520 238.270 2147.660 238.365 ;
        RECT 670.520 238.130 670.660 238.225 ;
        RECT 674.735 238.150 674.875 238.225 ;
        RECT 670.520 237.810 670.780 238.130 ;
        RECT 674.735 237.830 674.995 238.150 ;
        RECT 2147.520 237.950 2147.780 238.270 ;
        RECT 2152.880 237.990 2153.020 238.050 ;
        RECT 675.880 237.850 676.020 237.900 ;
        RECT 679.745 237.870 679.885 237.925 ;
        RECT 670.520 216.360 670.660 237.810 ;
        RECT 670.440 215.510 670.760 216.360 ;
        RECT 674.735 216.100 674.875 237.830 ;
        RECT 675.880 237.530 676.140 237.850 ;
        RECT 679.745 237.550 680.005 237.870 ;
        RECT 674.240 215.780 675.330 216.100 ;
        RECT 675.880 213.040 676.020 237.530 ;
        RECT 676.500 237.290 676.640 237.400 ;
        RECT 676.500 236.970 676.760 237.290 ;
        RECT 676.500 216.360 676.640 236.970 ;
        RECT 676.420 215.510 676.740 216.360 ;
        RECT 679.745 213.300 679.885 237.550 ;
        RECT 680.715 237.310 680.855 237.400 ;
        RECT 680.715 236.990 680.975 237.310 ;
        RECT 681.860 237.010 682.000 237.050 ;
        RECT 685.725 237.030 685.865 237.085 ;
        RECT 680.715 216.100 680.855 236.990 ;
        RECT 681.860 236.690 682.120 237.010 ;
        RECT 685.725 236.710 685.985 237.030 ;
        RECT 680.220 215.780 681.310 216.100 ;
        RECT 675.590 212.720 676.680 213.040 ;
        RECT 679.650 212.450 679.970 213.300 ;
        RECT 681.860 213.040 682.000 236.690 ;
        RECT 682.480 236.450 682.620 236.545 ;
        RECT 682.480 236.130 682.740 236.450 ;
        RECT 682.480 216.360 682.620 236.130 ;
        RECT 682.400 215.510 682.720 216.360 ;
        RECT 685.725 213.300 685.865 236.710 ;
        RECT 686.695 236.470 686.835 236.520 ;
        RECT 686.695 236.150 686.955 236.470 ;
        RECT 687.840 236.170 687.980 236.235 ;
        RECT 691.705 236.190 691.845 236.260 ;
        RECT 686.695 216.100 686.835 236.150 ;
        RECT 687.840 235.850 688.100 236.170 ;
        RECT 691.705 235.870 691.965 236.190 ;
        RECT 686.200 215.780 687.290 216.100 ;
        RECT 681.570 212.720 682.660 213.040 ;
        RECT 685.630 212.450 685.950 213.300 ;
        RECT 687.840 213.040 687.980 235.850 ;
        RECT 688.460 235.610 688.600 235.815 ;
        RECT 688.460 235.290 688.720 235.610 ;
        RECT 688.460 216.360 688.600 235.290 ;
        RECT 688.380 215.510 688.700 216.360 ;
        RECT 691.705 213.300 691.845 235.870 ;
        RECT 692.675 235.630 692.815 235.695 ;
        RECT 692.675 235.310 692.935 235.630 ;
        RECT 693.820 235.330 693.960 235.450 ;
        RECT 697.685 235.350 697.825 235.470 ;
        RECT 692.675 216.100 692.815 235.310 ;
        RECT 693.820 235.010 694.080 235.330 ;
        RECT 697.685 235.030 697.945 235.350 ;
        RECT 692.180 215.780 693.270 216.100 ;
        RECT 687.550 212.720 688.640 213.040 ;
        RECT 691.610 212.450 691.930 213.300 ;
        RECT 693.820 213.040 693.960 235.010 ;
        RECT 694.440 234.770 694.580 234.870 ;
        RECT 694.440 234.450 694.700 234.770 ;
        RECT 694.440 216.360 694.580 234.450 ;
        RECT 694.360 215.510 694.680 216.360 ;
        RECT 697.685 213.300 697.825 235.030 ;
        RECT 698.655 234.790 698.795 234.905 ;
        RECT 698.655 234.470 698.915 234.790 ;
        RECT 699.800 234.490 699.940 234.515 ;
        RECT 698.655 216.100 698.795 234.470 ;
        RECT 699.800 234.170 700.060 234.490 ;
        RECT 698.160 215.780 699.250 216.100 ;
        RECT 693.530 212.720 694.620 213.040 ;
        RECT 697.590 212.450 697.910 213.300 ;
        RECT 699.800 213.040 699.940 234.170 ;
        RECT 700.420 233.930 700.560 234.060 ;
        RECT 700.420 233.610 700.680 233.930 ;
        RECT 700.420 216.360 700.560 233.610 ;
        RECT 703.665 232.830 703.805 232.890 ;
        RECT 703.665 232.510 703.925 232.830 ;
        RECT 704.635 232.550 704.775 232.680 ;
        RECT 700.340 215.510 700.660 216.360 ;
        RECT 703.665 213.300 703.805 232.510 ;
        RECT 704.515 232.230 704.775 232.550 ;
        RECT 704.635 216.100 704.775 232.230 ;
        RECT 705.780 232.250 705.920 232.315 ;
        RECT 709.645 232.270 709.785 232.310 ;
        RECT 705.780 231.930 706.040 232.250 ;
        RECT 706.400 231.970 706.540 232.150 ;
        RECT 704.140 215.780 705.230 216.100 ;
        RECT 699.510 212.720 700.600 213.040 ;
        RECT 703.570 212.450 703.890 213.300 ;
        RECT 705.780 213.040 705.920 231.930 ;
        RECT 706.400 231.650 706.660 231.970 ;
        RECT 709.645 231.950 709.905 232.270 ;
        RECT 710.615 231.990 710.755 232.190 ;
        RECT 706.400 216.360 706.540 231.650 ;
        RECT 706.320 215.510 706.640 216.360 ;
        RECT 709.645 213.300 709.785 231.950 ;
        RECT 710.615 231.670 710.875 231.990 ;
        RECT 711.760 231.690 711.900 231.750 ;
        RECT 715.625 231.710 715.765 231.780 ;
        RECT 710.615 216.100 710.755 231.670 ;
        RECT 711.760 231.370 712.020 231.690 ;
        RECT 712.380 231.410 712.520 231.505 ;
        RECT 710.120 215.780 711.210 216.100 ;
        RECT 705.490 212.720 706.580 213.040 ;
        RECT 709.550 212.450 709.870 213.300 ;
        RECT 711.760 213.040 711.900 231.370 ;
        RECT 712.380 231.090 712.640 231.410 ;
        RECT 715.625 231.390 715.885 231.710 ;
        RECT 716.595 231.430 716.735 231.525 ;
        RECT 712.380 216.360 712.520 231.090 ;
        RECT 712.300 215.510 712.620 216.360 ;
        RECT 715.625 213.300 715.765 231.390 ;
        RECT 716.475 231.110 716.735 231.430 ;
        RECT 716.595 216.100 716.735 231.110 ;
        RECT 717.740 231.130 717.880 232.345 ;
        RECT 717.740 230.810 718.000 231.130 ;
        RECT 718.360 230.850 718.500 232.345 ;
        RECT 721.605 231.150 721.745 232.345 ;
        RECT 716.100 215.780 717.190 216.100 ;
        RECT 711.470 212.720 712.560 213.040 ;
        RECT 715.530 212.450 715.850 213.300 ;
        RECT 717.740 213.040 717.880 230.810 ;
        RECT 718.360 230.530 718.620 230.850 ;
        RECT 721.605 230.830 721.865 231.150 ;
        RECT 722.575 230.870 722.715 232.345 ;
        RECT 718.360 216.360 718.500 230.530 ;
        RECT 718.280 215.510 718.600 216.360 ;
        RECT 721.605 213.300 721.745 230.830 ;
        RECT 722.575 230.550 722.835 230.870 ;
        RECT 723.720 230.570 723.860 232.345 ;
        RECT 722.575 216.100 722.715 230.550 ;
        RECT 723.720 230.250 723.980 230.570 ;
        RECT 724.340 230.290 724.480 232.345 ;
        RECT 727.585 230.590 727.725 232.345 ;
        RECT 722.080 215.780 723.170 216.100 ;
        RECT 717.450 212.720 718.540 213.040 ;
        RECT 721.510 212.450 721.830 213.300 ;
        RECT 723.720 213.040 723.860 230.250 ;
        RECT 724.340 229.970 724.600 230.290 ;
        RECT 727.585 230.270 727.845 230.590 ;
        RECT 728.555 230.310 728.695 232.345 ;
        RECT 724.340 216.360 724.480 229.970 ;
        RECT 724.260 215.510 724.580 216.360 ;
        RECT 727.585 213.300 727.725 230.270 ;
        RECT 728.555 229.990 728.815 230.310 ;
        RECT 729.700 230.010 729.840 232.345 ;
        RECT 728.555 216.100 728.695 229.990 ;
        RECT 729.700 229.690 729.960 230.010 ;
        RECT 730.320 229.730 730.460 232.345 ;
        RECT 733.565 230.030 733.705 232.345 ;
        RECT 728.060 215.780 729.150 216.100 ;
        RECT 723.430 212.720 724.520 213.040 ;
        RECT 727.490 212.450 727.810 213.300 ;
        RECT 729.700 213.040 729.840 229.690 ;
        RECT 730.320 229.410 730.580 229.730 ;
        RECT 733.565 229.710 733.825 230.030 ;
        RECT 734.535 229.750 734.675 232.345 ;
        RECT 730.320 216.360 730.460 229.410 ;
        RECT 730.240 215.510 730.560 216.360 ;
        RECT 733.565 213.300 733.705 229.710 ;
        RECT 734.535 229.430 734.795 229.750 ;
        RECT 735.680 229.450 735.820 232.345 ;
        RECT 734.535 216.100 734.675 229.430 ;
        RECT 735.680 229.130 735.940 229.450 ;
        RECT 734.040 215.780 735.130 216.100 ;
        RECT 729.410 212.720 730.500 213.040 ;
        RECT 733.470 212.450 733.790 213.300 ;
        RECT 735.680 213.040 735.820 229.130 ;
        RECT 736.300 228.890 736.440 232.345 ;
        RECT 739.545 229.470 739.685 232.345 ;
        RECT 739.545 229.150 739.805 229.470 ;
        RECT 736.300 228.570 736.560 228.890 ;
        RECT 736.300 216.360 736.440 228.570 ;
        RECT 736.220 215.510 736.540 216.360 ;
        RECT 739.545 213.300 739.685 229.150 ;
        RECT 740.515 228.910 740.655 232.345 ;
        RECT 740.515 228.590 740.775 228.910 ;
        RECT 741.660 228.610 741.800 232.345 ;
        RECT 740.515 216.100 740.655 228.590 ;
        RECT 741.660 228.290 741.920 228.610 ;
        RECT 740.020 215.780 741.110 216.100 ;
        RECT 735.390 212.720 736.480 213.040 ;
        RECT 739.450 212.450 739.770 213.300 ;
        RECT 741.660 213.040 741.800 228.290 ;
        RECT 742.280 228.050 742.420 232.345 ;
        RECT 745.525 228.630 745.665 232.345 ;
        RECT 745.525 228.310 745.785 228.630 ;
        RECT 742.280 227.730 742.540 228.050 ;
        RECT 742.280 216.360 742.420 227.730 ;
        RECT 742.200 215.510 742.520 216.360 ;
        RECT 745.525 213.300 745.665 228.310 ;
        RECT 746.495 228.070 746.635 232.345 ;
        RECT 746.495 227.750 746.755 228.070 ;
        RECT 747.640 227.770 747.780 232.345 ;
        RECT 746.495 216.100 746.635 227.750 ;
        RECT 747.640 227.450 747.900 227.770 ;
        RECT 746.000 215.780 747.090 216.100 ;
        RECT 741.370 212.720 742.460 213.040 ;
        RECT 745.430 212.450 745.750 213.300 ;
        RECT 747.640 213.040 747.780 227.450 ;
        RECT 748.260 227.210 748.400 232.345 ;
        RECT 751.505 227.790 751.645 232.345 ;
        RECT 751.505 227.470 751.765 227.790 ;
        RECT 748.260 226.890 748.520 227.210 ;
        RECT 748.260 216.360 748.400 226.890 ;
        RECT 748.180 215.510 748.500 216.360 ;
        RECT 751.505 213.300 751.645 227.470 ;
        RECT 752.475 227.230 752.615 232.345 ;
        RECT 752.475 226.910 752.735 227.230 ;
        RECT 753.620 226.930 753.760 232.345 ;
        RECT 752.475 216.100 752.615 226.910 ;
        RECT 753.620 226.610 753.880 226.930 ;
        RECT 751.980 215.780 753.070 216.100 ;
        RECT 747.350 212.720 748.440 213.040 ;
        RECT 751.410 212.450 751.730 213.300 ;
        RECT 753.620 213.040 753.760 226.610 ;
        RECT 754.240 226.370 754.380 232.345 ;
        RECT 757.485 226.950 757.625 232.345 ;
        RECT 757.485 226.630 757.745 226.950 ;
        RECT 754.240 226.050 754.500 226.370 ;
        RECT 754.240 216.360 754.380 226.050 ;
        RECT 754.160 215.510 754.480 216.360 ;
        RECT 757.485 213.300 757.625 226.630 ;
        RECT 758.455 226.390 758.595 232.345 ;
        RECT 758.455 226.070 758.715 226.390 ;
        RECT 759.600 226.090 759.740 232.345 ;
        RECT 763.465 226.110 763.605 232.345 ;
        RECT 758.455 216.100 758.595 226.070 ;
        RECT 759.600 225.770 759.860 226.090 ;
        RECT 763.465 225.790 763.725 226.110 ;
        RECT 757.960 215.780 759.050 216.100 ;
        RECT 753.330 212.720 754.420 213.040 ;
        RECT 757.390 212.450 757.710 213.300 ;
        RECT 759.600 213.040 759.740 225.770 ;
        RECT 763.465 213.300 763.605 225.790 ;
        RECT 764.435 225.550 764.575 232.345 ;
        RECT 764.435 225.230 764.695 225.550 ;
        RECT 769.445 225.270 769.585 232.345 ;
        RECT 764.435 216.100 764.575 225.230 ;
        RECT 769.445 224.950 769.705 225.270 ;
        RECT 763.940 215.780 765.030 216.100 ;
        RECT 769.445 213.300 769.585 224.950 ;
        RECT 770.415 224.710 770.555 232.345 ;
        RECT 770.415 224.390 770.675 224.710 ;
        RECT 775.425 224.430 775.565 232.345 ;
        RECT 770.415 216.100 770.555 224.390 ;
        RECT 775.425 224.110 775.685 224.430 ;
        RECT 769.920 215.780 771.010 216.100 ;
        RECT 775.425 213.300 775.565 224.110 ;
        RECT 776.395 223.870 776.535 232.345 ;
        RECT 776.275 223.550 776.535 223.870 ;
        RECT 776.395 216.100 776.535 223.550 ;
        RECT 781.405 223.590 781.545 232.345 ;
        RECT 781.405 223.270 781.665 223.590 ;
        RECT 775.900 215.780 776.990 216.100 ;
        RECT 781.405 213.300 781.545 223.270 ;
        RECT 782.375 223.030 782.515 232.345 ;
        RECT 782.375 222.710 782.635 223.030 ;
        RECT 787.385 222.750 787.525 232.345 ;
        RECT 782.375 216.100 782.515 222.710 ;
        RECT 787.385 222.430 787.645 222.750 ;
        RECT 781.880 215.780 782.970 216.100 ;
        RECT 787.385 213.300 787.525 222.430 ;
        RECT 788.355 222.190 788.495 232.345 ;
        RECT 788.235 221.870 788.495 222.190 ;
        RECT 788.355 216.100 788.495 221.870 ;
        RECT 793.365 221.630 793.505 232.345 ;
        RECT 793.365 221.310 793.625 221.630 ;
        RECT 787.860 215.780 788.950 216.100 ;
        RECT 793.365 214.240 793.505 221.310 ;
        RECT 794.335 221.070 794.475 232.345 ;
        RECT 794.335 220.750 794.595 221.070 ;
        RECT 794.335 216.100 794.475 220.750 ;
        RECT 2147.520 216.360 2147.660 237.950 ;
        RECT 2152.880 237.670 2153.140 237.990 ;
        RECT 793.840 215.780 794.930 216.100 ;
        RECT 2147.440 215.510 2147.760 216.360 ;
        RECT 793.365 214.100 794.140 214.240 ;
        RECT 759.310 212.720 760.400 213.040 ;
        RECT 763.370 212.450 763.690 213.300 ;
        RECT 769.350 212.450 769.670 213.300 ;
        RECT 775.330 212.450 775.650 213.300 ;
        RECT 781.310 212.450 781.630 213.300 ;
        RECT 787.290 212.450 787.610 213.300 ;
        RECT 794.000 213.040 794.140 214.100 ;
        RECT 2152.880 213.040 2153.020 237.670 ;
        RECT 2153.500 237.430 2153.640 237.525 ;
        RECT 2153.500 237.110 2153.760 237.430 ;
        RECT 2158.860 237.150 2159.000 237.235 ;
        RECT 2153.500 216.360 2153.640 237.110 ;
        RECT 2158.860 236.830 2159.120 237.150 ;
        RECT 2153.420 215.510 2153.740 216.360 ;
        RECT 2158.860 213.040 2159.000 236.830 ;
        RECT 2159.480 236.590 2159.620 236.705 ;
        RECT 2159.480 236.270 2159.740 236.590 ;
        RECT 2164.840 236.310 2164.980 236.395 ;
        RECT 2159.480 216.360 2159.620 236.270 ;
        RECT 2164.840 235.990 2165.100 236.310 ;
        RECT 2159.400 215.510 2159.720 216.360 ;
        RECT 2164.840 213.040 2164.980 235.990 ;
        RECT 2165.460 235.750 2165.600 235.815 ;
        RECT 2165.460 235.430 2165.720 235.750 ;
        RECT 2170.820 235.470 2170.960 235.540 ;
        RECT 2165.460 216.360 2165.600 235.430 ;
        RECT 2170.820 235.150 2171.080 235.470 ;
        RECT 2165.380 215.510 2165.700 216.360 ;
        RECT 2170.820 213.040 2170.960 235.150 ;
        RECT 2171.440 234.910 2171.580 234.990 ;
        RECT 2171.440 234.590 2171.700 234.910 ;
        RECT 2176.800 234.630 2176.940 234.675 ;
        RECT 2171.440 216.360 2171.580 234.590 ;
        RECT 2176.800 234.310 2177.060 234.630 ;
        RECT 2171.360 215.510 2171.680 216.360 ;
        RECT 2176.800 213.040 2176.940 234.310 ;
        RECT 2177.420 234.070 2177.560 234.180 ;
        RECT 2177.420 233.750 2177.680 234.070 ;
        RECT 2182.780 233.790 2182.920 233.845 ;
        RECT 2177.420 216.360 2177.560 233.750 ;
        RECT 2182.780 233.470 2183.040 233.790 ;
        RECT 2177.340 215.510 2177.660 216.360 ;
        RECT 2182.780 213.040 2182.920 233.470 ;
        RECT 2183.400 233.230 2183.540 233.310 ;
        RECT 2183.400 232.910 2183.660 233.230 ;
        RECT 2188.760 232.950 2188.900 233.000 ;
        RECT 2183.400 216.360 2183.540 232.910 ;
        RECT 2188.760 232.630 2189.020 232.950 ;
        RECT 2183.320 215.510 2183.640 216.360 ;
        RECT 2188.760 213.040 2188.900 232.630 ;
        RECT 2189.380 232.390 2189.520 232.485 ;
        RECT 2189.380 232.070 2189.640 232.390 ;
        RECT 2194.740 232.110 2194.880 232.485 ;
        RECT 2189.380 216.360 2189.520 232.070 ;
        RECT 2194.740 231.790 2195.000 232.110 ;
        RECT 2189.300 215.510 2189.620 216.360 ;
        RECT 2194.740 213.040 2194.880 231.790 ;
        RECT 2195.360 231.550 2195.500 232.485 ;
        RECT 2195.360 231.230 2195.620 231.550 ;
        RECT 2200.720 231.270 2200.860 232.485 ;
        RECT 2195.360 216.360 2195.500 231.230 ;
        RECT 2200.720 230.950 2200.980 231.270 ;
        RECT 2195.280 215.510 2195.600 216.360 ;
        RECT 2200.720 213.040 2200.860 230.950 ;
        RECT 2201.340 230.710 2201.480 232.485 ;
        RECT 2201.340 230.390 2201.600 230.710 ;
        RECT 2206.700 230.430 2206.840 232.485 ;
        RECT 2201.340 216.360 2201.480 230.390 ;
        RECT 2206.700 230.110 2206.960 230.430 ;
        RECT 2201.260 215.510 2201.580 216.360 ;
        RECT 2206.700 213.040 2206.840 230.110 ;
        RECT 2207.320 229.870 2207.460 232.485 ;
        RECT 2207.320 229.550 2207.580 229.870 ;
        RECT 2212.680 229.590 2212.820 232.485 ;
        RECT 2207.320 216.360 2207.460 229.550 ;
        RECT 2212.680 229.270 2212.940 229.590 ;
        RECT 2207.240 215.510 2207.560 216.360 ;
        RECT 2212.680 213.040 2212.820 229.270 ;
        RECT 2213.300 229.030 2213.440 232.485 ;
        RECT 2213.300 228.710 2213.560 229.030 ;
        RECT 2218.660 228.750 2218.800 232.485 ;
        RECT 2213.300 216.360 2213.440 228.710 ;
        RECT 2218.660 228.430 2218.920 228.750 ;
        RECT 2213.220 215.510 2213.540 216.360 ;
        RECT 2218.660 213.040 2218.800 228.430 ;
        RECT 2219.280 228.190 2219.420 232.485 ;
        RECT 2219.280 227.870 2219.540 228.190 ;
        RECT 2224.640 227.910 2224.780 232.485 ;
        RECT 2219.280 216.360 2219.420 227.870 ;
        RECT 2224.640 227.590 2224.900 227.910 ;
        RECT 2219.200 215.510 2219.520 216.360 ;
        RECT 2224.640 213.040 2224.780 227.590 ;
        RECT 2225.260 227.350 2225.400 232.485 ;
        RECT 2225.260 227.030 2225.520 227.350 ;
        RECT 2230.620 227.070 2230.760 232.485 ;
        RECT 2225.260 216.360 2225.400 227.030 ;
        RECT 2230.620 226.750 2230.880 227.070 ;
        RECT 2225.180 215.510 2225.500 216.360 ;
        RECT 2230.620 213.040 2230.760 226.750 ;
        RECT 2231.240 226.510 2231.380 232.485 ;
        RECT 2231.240 226.190 2231.500 226.510 ;
        RECT 2236.600 226.230 2236.740 232.485 ;
        RECT 2231.240 216.360 2231.380 226.190 ;
        RECT 2236.600 225.910 2236.860 226.230 ;
        RECT 2231.160 215.510 2231.480 216.360 ;
        RECT 2236.600 213.040 2236.740 225.910 ;
        RECT 2237.220 225.670 2237.360 232.485 ;
        RECT 2237.220 225.350 2237.480 225.670 ;
        RECT 2242.580 225.390 2242.720 232.485 ;
        RECT 2237.220 216.360 2237.360 225.350 ;
        RECT 2242.580 225.070 2242.840 225.390 ;
        RECT 2237.140 215.510 2237.460 216.360 ;
        RECT 2242.580 213.040 2242.720 225.070 ;
        RECT 2243.200 224.830 2243.340 232.485 ;
        RECT 2243.200 224.510 2243.460 224.830 ;
        RECT 2248.560 224.550 2248.700 232.485 ;
        RECT 2243.200 216.360 2243.340 224.510 ;
        RECT 2248.560 224.230 2248.820 224.550 ;
        RECT 2243.120 215.510 2243.440 216.360 ;
        RECT 2248.560 213.040 2248.700 224.230 ;
        RECT 2249.180 223.990 2249.320 232.485 ;
        RECT 2249.180 223.670 2249.440 223.990 ;
        RECT 2254.540 223.710 2254.680 232.485 ;
        RECT 2249.180 216.360 2249.320 223.670 ;
        RECT 2254.540 223.390 2254.800 223.710 ;
        RECT 2249.100 215.510 2249.420 216.360 ;
        RECT 2254.540 213.040 2254.680 223.390 ;
        RECT 2255.160 223.150 2255.300 232.485 ;
        RECT 2255.160 222.830 2255.420 223.150 ;
        RECT 2260.520 222.870 2260.660 232.485 ;
        RECT 2255.160 216.360 2255.300 222.830 ;
        RECT 2260.520 222.550 2260.780 222.870 ;
        RECT 2255.080 215.510 2255.400 216.360 ;
        RECT 2260.520 213.040 2260.660 222.550 ;
        RECT 2261.140 222.310 2261.280 232.485 ;
        RECT 2261.140 221.990 2261.400 222.310 ;
        RECT 2261.140 216.360 2261.280 221.990 ;
        RECT 2266.500 221.750 2266.640 232.485 ;
        RECT 2266.500 221.430 2266.760 221.750 ;
        RECT 2261.060 215.510 2261.380 216.360 ;
        RECT 2266.500 214.170 2266.640 221.430 ;
        RECT 2267.120 221.190 2267.260 232.485 ;
        RECT 2267.120 220.870 2267.380 221.190 ;
        RECT 2267.120 216.360 2267.260 220.870 ;
        RECT 2267.040 215.510 2267.360 216.360 ;
        RECT 2266.500 214.030 2267.275 214.170 ;
        RECT 2267.135 213.300 2267.275 214.030 ;
        RECT 793.340 212.720 794.430 213.040 ;
        RECT 2152.590 212.720 2153.680 213.040 ;
        RECT 2158.570 212.720 2159.660 213.040 ;
        RECT 2164.550 212.720 2165.640 213.040 ;
        RECT 2170.530 212.720 2171.620 213.040 ;
        RECT 2176.510 212.720 2177.600 213.040 ;
        RECT 2182.490 212.720 2183.580 213.040 ;
        RECT 2188.470 212.720 2189.560 213.040 ;
        RECT 2194.450 212.720 2195.540 213.040 ;
        RECT 2200.430 212.720 2201.520 213.040 ;
        RECT 2206.410 212.720 2207.500 213.040 ;
        RECT 2212.390 212.720 2213.480 213.040 ;
        RECT 2218.370 212.720 2219.460 213.040 ;
        RECT 2224.350 212.720 2225.440 213.040 ;
        RECT 2230.330 212.720 2231.420 213.040 ;
        RECT 2236.310 212.720 2237.400 213.040 ;
        RECT 2242.290 212.720 2243.380 213.040 ;
        RECT 2248.270 212.720 2249.360 213.040 ;
        RECT 2254.250 212.720 2255.340 213.040 ;
        RECT 2260.230 212.720 2261.320 213.040 ;
        RECT 2267.050 212.450 2267.370 213.300 ;
  END
END gpio_signal_buffering
END LIBRARY

