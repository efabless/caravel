module mgmt_protect (caravel_clk,
    caravel_clk2,
    caravel_rstn,
    mprj_ack_i_core,
    mprj_ack_i_user,
    mprj_cyc_o_core,
    mprj_cyc_o_user,
    mprj_iena_wb,
    mprj_stb_o_core,
    mprj_stb_o_user,
    mprj_we_o_core,
    mprj_we_o_user,
    user1_vcc_powergood,
    user1_vdd_powergood,
    user2_vcc_powergood,
    user2_vdd_powergood,
    user_clock,
    user_clock2,
    user_reset,
    la_data_in_core,
    la_data_in_mprj,
    la_data_out_core,
    la_data_out_mprj,
    la_iena_mprj,
    la_oenb_core,
    la_oenb_mprj,
    mprj_adr_o_core,
    mprj_adr_o_user,
    mprj_dat_i_core,
    mprj_dat_i_user,
    mprj_dat_o_core,
    mprj_dat_o_user,
    mprj_sel_o_core,
    mprj_sel_o_user,
    user_irq,
    user_irq_core,
    user_irq_ena);
 input caravel_clk;
 input caravel_clk2;
 input caravel_rstn;
 output mprj_ack_i_core;
 input mprj_ack_i_user;
 input mprj_cyc_o_core;
 output mprj_cyc_o_user;
 input mprj_iena_wb;
 input mprj_stb_o_core;
 output mprj_stb_o_user;
 input mprj_we_o_core;
 output mprj_we_o_user;
 output user1_vcc_powergood;
 output user1_vdd_powergood;
 output user2_vcc_powergood;
 output user2_vdd_powergood;
 output user_clock;
 output user_clock2;
 output user_reset;
 output [127:0] la_data_in_core;
 output [127:0] la_data_in_mprj;
 input [127:0] la_data_out_core;
 input [127:0] la_data_out_mprj;
 input [127:0] la_iena_mprj;
 output [127:0] la_oenb_core;
 input [127:0] la_oenb_mprj;
 input [31:0] mprj_adr_o_core;
 output [31:0] mprj_adr_o_user;
 output [31:0] mprj_dat_i_core;
 input [31:0] mprj_dat_i_user;
 input [31:0] mprj_dat_o_core;
 output [31:0] mprj_dat_o_user;
 input [3:0] mprj_sel_o_core;
 output [3:0] mprj_sel_o_user;
 output [2:0] user_irq;
 input [2:0] user_irq_core;
 input [2:0] user_irq_ena;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire \la_data_in_enable[0] ;
 wire \la_data_in_enable[100] ;
 wire \la_data_in_enable[101] ;
 wire \la_data_in_enable[102] ;
 wire \la_data_in_enable[103] ;
 wire \la_data_in_enable[104] ;
 wire \la_data_in_enable[105] ;
 wire \la_data_in_enable[106] ;
 wire \la_data_in_enable[107] ;
 wire \la_data_in_enable[108] ;
 wire \la_data_in_enable[109] ;
 wire \la_data_in_enable[10] ;
 wire \la_data_in_enable[110] ;
 wire \la_data_in_enable[111] ;
 wire \la_data_in_enable[112] ;
 wire \la_data_in_enable[113] ;
 wire \la_data_in_enable[114] ;
 wire \la_data_in_enable[115] ;
 wire \la_data_in_enable[116] ;
 wire \la_data_in_enable[117] ;
 wire \la_data_in_enable[118] ;
 wire \la_data_in_enable[119] ;
 wire \la_data_in_enable[11] ;
 wire \la_data_in_enable[120] ;
 wire \la_data_in_enable[121] ;
 wire \la_data_in_enable[122] ;
 wire \la_data_in_enable[123] ;
 wire \la_data_in_enable[124] ;
 wire \la_data_in_enable[125] ;
 wire \la_data_in_enable[126] ;
 wire \la_data_in_enable[127] ;
 wire \la_data_in_enable[12] ;
 wire \la_data_in_enable[13] ;
 wire \la_data_in_enable[14] ;
 wire \la_data_in_enable[15] ;
 wire \la_data_in_enable[16] ;
 wire \la_data_in_enable[17] ;
 wire \la_data_in_enable[18] ;
 wire \la_data_in_enable[19] ;
 wire \la_data_in_enable[1] ;
 wire \la_data_in_enable[20] ;
 wire \la_data_in_enable[21] ;
 wire \la_data_in_enable[22] ;
 wire \la_data_in_enable[23] ;
 wire \la_data_in_enable[24] ;
 wire \la_data_in_enable[25] ;
 wire \la_data_in_enable[26] ;
 wire \la_data_in_enable[27] ;
 wire \la_data_in_enable[28] ;
 wire \la_data_in_enable[29] ;
 wire \la_data_in_enable[2] ;
 wire \la_data_in_enable[30] ;
 wire \la_data_in_enable[31] ;
 wire \la_data_in_enable[32] ;
 wire \la_data_in_enable[33] ;
 wire \la_data_in_enable[34] ;
 wire \la_data_in_enable[35] ;
 wire \la_data_in_enable[36] ;
 wire \la_data_in_enable[37] ;
 wire \la_data_in_enable[38] ;
 wire \la_data_in_enable[39] ;
 wire \la_data_in_enable[3] ;
 wire \la_data_in_enable[40] ;
 wire \la_data_in_enable[41] ;
 wire \la_data_in_enable[42] ;
 wire \la_data_in_enable[43] ;
 wire \la_data_in_enable[44] ;
 wire \la_data_in_enable[45] ;
 wire \la_data_in_enable[46] ;
 wire \la_data_in_enable[47] ;
 wire \la_data_in_enable[48] ;
 wire \la_data_in_enable[49] ;
 wire \la_data_in_enable[4] ;
 wire \la_data_in_enable[50] ;
 wire \la_data_in_enable[51] ;
 wire \la_data_in_enable[52] ;
 wire \la_data_in_enable[53] ;
 wire \la_data_in_enable[54] ;
 wire \la_data_in_enable[55] ;
 wire \la_data_in_enable[56] ;
 wire \la_data_in_enable[57] ;
 wire \la_data_in_enable[58] ;
 wire \la_data_in_enable[59] ;
 wire \la_data_in_enable[5] ;
 wire \la_data_in_enable[60] ;
 wire \la_data_in_enable[61] ;
 wire \la_data_in_enable[62] ;
 wire \la_data_in_enable[63] ;
 wire \la_data_in_enable[64] ;
 wire \la_data_in_enable[65] ;
 wire \la_data_in_enable[66] ;
 wire \la_data_in_enable[67] ;
 wire \la_data_in_enable[68] ;
 wire \la_data_in_enable[69] ;
 wire \la_data_in_enable[6] ;
 wire \la_data_in_enable[70] ;
 wire \la_data_in_enable[71] ;
 wire \la_data_in_enable[72] ;
 wire \la_data_in_enable[73] ;
 wire \la_data_in_enable[74] ;
 wire \la_data_in_enable[75] ;
 wire \la_data_in_enable[76] ;
 wire \la_data_in_enable[77] ;
 wire \la_data_in_enable[78] ;
 wire \la_data_in_enable[79] ;
 wire \la_data_in_enable[7] ;
 wire \la_data_in_enable[80] ;
 wire \la_data_in_enable[81] ;
 wire \la_data_in_enable[82] ;
 wire \la_data_in_enable[83] ;
 wire \la_data_in_enable[84] ;
 wire \la_data_in_enable[85] ;
 wire \la_data_in_enable[86] ;
 wire \la_data_in_enable[87] ;
 wire \la_data_in_enable[88] ;
 wire \la_data_in_enable[89] ;
 wire \la_data_in_enable[8] ;
 wire \la_data_in_enable[90] ;
 wire \la_data_in_enable[91] ;
 wire \la_data_in_enable[92] ;
 wire \la_data_in_enable[93] ;
 wire \la_data_in_enable[94] ;
 wire \la_data_in_enable[95] ;
 wire \la_data_in_enable[96] ;
 wire \la_data_in_enable[97] ;
 wire \la_data_in_enable[98] ;
 wire \la_data_in_enable[99] ;
 wire \la_data_in_enable[9] ;
 wire \la_data_in_mprj_bar[0] ;
 wire \la_data_in_mprj_bar[100] ;
 wire \la_data_in_mprj_bar[101] ;
 wire \la_data_in_mprj_bar[102] ;
 wire \la_data_in_mprj_bar[103] ;
 wire \la_data_in_mprj_bar[104] ;
 wire \la_data_in_mprj_bar[105] ;
 wire \la_data_in_mprj_bar[106] ;
 wire \la_data_in_mprj_bar[107] ;
 wire \la_data_in_mprj_bar[108] ;
 wire \la_data_in_mprj_bar[109] ;
 wire \la_data_in_mprj_bar[10] ;
 wire \la_data_in_mprj_bar[110] ;
 wire \la_data_in_mprj_bar[111] ;
 wire \la_data_in_mprj_bar[112] ;
 wire \la_data_in_mprj_bar[113] ;
 wire \la_data_in_mprj_bar[114] ;
 wire \la_data_in_mprj_bar[115] ;
 wire \la_data_in_mprj_bar[116] ;
 wire \la_data_in_mprj_bar[117] ;
 wire \la_data_in_mprj_bar[118] ;
 wire \la_data_in_mprj_bar[119] ;
 wire \la_data_in_mprj_bar[11] ;
 wire \la_data_in_mprj_bar[120] ;
 wire \la_data_in_mprj_bar[121] ;
 wire \la_data_in_mprj_bar[122] ;
 wire \la_data_in_mprj_bar[123] ;
 wire \la_data_in_mprj_bar[124] ;
 wire \la_data_in_mprj_bar[125] ;
 wire \la_data_in_mprj_bar[126] ;
 wire \la_data_in_mprj_bar[127] ;
 wire \la_data_in_mprj_bar[12] ;
 wire \la_data_in_mprj_bar[13] ;
 wire \la_data_in_mprj_bar[14] ;
 wire \la_data_in_mprj_bar[15] ;
 wire \la_data_in_mprj_bar[16] ;
 wire \la_data_in_mprj_bar[17] ;
 wire \la_data_in_mprj_bar[18] ;
 wire \la_data_in_mprj_bar[19] ;
 wire \la_data_in_mprj_bar[1] ;
 wire \la_data_in_mprj_bar[20] ;
 wire \la_data_in_mprj_bar[21] ;
 wire \la_data_in_mprj_bar[22] ;
 wire \la_data_in_mprj_bar[23] ;
 wire \la_data_in_mprj_bar[24] ;
 wire \la_data_in_mprj_bar[25] ;
 wire \la_data_in_mprj_bar[26] ;
 wire \la_data_in_mprj_bar[27] ;
 wire \la_data_in_mprj_bar[28] ;
 wire \la_data_in_mprj_bar[29] ;
 wire \la_data_in_mprj_bar[2] ;
 wire \la_data_in_mprj_bar[30] ;
 wire \la_data_in_mprj_bar[31] ;
 wire \la_data_in_mprj_bar[32] ;
 wire \la_data_in_mprj_bar[33] ;
 wire \la_data_in_mprj_bar[34] ;
 wire \la_data_in_mprj_bar[35] ;
 wire \la_data_in_mprj_bar[36] ;
 wire \la_data_in_mprj_bar[37] ;
 wire \la_data_in_mprj_bar[38] ;
 wire \la_data_in_mprj_bar[39] ;
 wire \la_data_in_mprj_bar[3] ;
 wire \la_data_in_mprj_bar[40] ;
 wire \la_data_in_mprj_bar[41] ;
 wire \la_data_in_mprj_bar[42] ;
 wire \la_data_in_mprj_bar[43] ;
 wire \la_data_in_mprj_bar[44] ;
 wire \la_data_in_mprj_bar[45] ;
 wire \la_data_in_mprj_bar[46] ;
 wire \la_data_in_mprj_bar[47] ;
 wire \la_data_in_mprj_bar[48] ;
 wire \la_data_in_mprj_bar[49] ;
 wire \la_data_in_mprj_bar[4] ;
 wire \la_data_in_mprj_bar[50] ;
 wire \la_data_in_mprj_bar[51] ;
 wire \la_data_in_mprj_bar[52] ;
 wire \la_data_in_mprj_bar[53] ;
 wire \la_data_in_mprj_bar[54] ;
 wire \la_data_in_mprj_bar[55] ;
 wire \la_data_in_mprj_bar[56] ;
 wire \la_data_in_mprj_bar[57] ;
 wire \la_data_in_mprj_bar[58] ;
 wire \la_data_in_mprj_bar[59] ;
 wire \la_data_in_mprj_bar[5] ;
 wire \la_data_in_mprj_bar[60] ;
 wire \la_data_in_mprj_bar[61] ;
 wire \la_data_in_mprj_bar[62] ;
 wire \la_data_in_mprj_bar[63] ;
 wire \la_data_in_mprj_bar[64] ;
 wire \la_data_in_mprj_bar[65] ;
 wire \la_data_in_mprj_bar[66] ;
 wire \la_data_in_mprj_bar[67] ;
 wire \la_data_in_mprj_bar[68] ;
 wire \la_data_in_mprj_bar[69] ;
 wire \la_data_in_mprj_bar[6] ;
 wire \la_data_in_mprj_bar[70] ;
 wire \la_data_in_mprj_bar[71] ;
 wire \la_data_in_mprj_bar[72] ;
 wire \la_data_in_mprj_bar[73] ;
 wire \la_data_in_mprj_bar[74] ;
 wire \la_data_in_mprj_bar[75] ;
 wire \la_data_in_mprj_bar[76] ;
 wire \la_data_in_mprj_bar[77] ;
 wire \la_data_in_mprj_bar[78] ;
 wire \la_data_in_mprj_bar[79] ;
 wire \la_data_in_mprj_bar[7] ;
 wire \la_data_in_mprj_bar[80] ;
 wire \la_data_in_mprj_bar[81] ;
 wire \la_data_in_mprj_bar[82] ;
 wire \la_data_in_mprj_bar[83] ;
 wire \la_data_in_mprj_bar[84] ;
 wire \la_data_in_mprj_bar[85] ;
 wire \la_data_in_mprj_bar[86] ;
 wire \la_data_in_mprj_bar[87] ;
 wire \la_data_in_mprj_bar[88] ;
 wire \la_data_in_mprj_bar[89] ;
 wire \la_data_in_mprj_bar[8] ;
 wire \la_data_in_mprj_bar[90] ;
 wire \la_data_in_mprj_bar[91] ;
 wire \la_data_in_mprj_bar[92] ;
 wire \la_data_in_mprj_bar[93] ;
 wire \la_data_in_mprj_bar[94] ;
 wire \la_data_in_mprj_bar[95] ;
 wire \la_data_in_mprj_bar[96] ;
 wire \la_data_in_mprj_bar[97] ;
 wire \la_data_in_mprj_bar[98] ;
 wire \la_data_in_mprj_bar[99] ;
 wire \la_data_in_mprj_bar[9] ;
 wire mprj_ack_i_core_bar;
 wire \mprj_dat_i_core_bar[0] ;
 wire \mprj_dat_i_core_bar[10] ;
 wire \mprj_dat_i_core_bar[11] ;
 wire \mprj_dat_i_core_bar[12] ;
 wire \mprj_dat_i_core_bar[13] ;
 wire \mprj_dat_i_core_bar[14] ;
 wire \mprj_dat_i_core_bar[15] ;
 wire \mprj_dat_i_core_bar[16] ;
 wire \mprj_dat_i_core_bar[17] ;
 wire \mprj_dat_i_core_bar[18] ;
 wire \mprj_dat_i_core_bar[19] ;
 wire \mprj_dat_i_core_bar[1] ;
 wire \mprj_dat_i_core_bar[20] ;
 wire \mprj_dat_i_core_bar[21] ;
 wire \mprj_dat_i_core_bar[22] ;
 wire \mprj_dat_i_core_bar[23] ;
 wire \mprj_dat_i_core_bar[24] ;
 wire \mprj_dat_i_core_bar[25] ;
 wire \mprj_dat_i_core_bar[26] ;
 wire \mprj_dat_i_core_bar[27] ;
 wire \mprj_dat_i_core_bar[28] ;
 wire \mprj_dat_i_core_bar[29] ;
 wire \mprj_dat_i_core_bar[2] ;
 wire \mprj_dat_i_core_bar[30] ;
 wire \mprj_dat_i_core_bar[31] ;
 wire \mprj_dat_i_core_bar[3] ;
 wire \mprj_dat_i_core_bar[4] ;
 wire \mprj_dat_i_core_bar[5] ;
 wire \mprj_dat_i_core_bar[6] ;
 wire \mprj_dat_i_core_bar[7] ;
 wire \mprj_dat_i_core_bar[8] ;
 wire \mprj_dat_i_core_bar[9] ;
 wire \mprj_logic1[0] ;
 wire \mprj_logic1[100] ;
 wire \mprj_logic1[101] ;
 wire \mprj_logic1[102] ;
 wire \mprj_logic1[103] ;
 wire \mprj_logic1[104] ;
 wire \mprj_logic1[105] ;
 wire \mprj_logic1[106] ;
 wire \mprj_logic1[107] ;
 wire \mprj_logic1[108] ;
 wire \mprj_logic1[109] ;
 wire \mprj_logic1[10] ;
 wire \mprj_logic1[110] ;
 wire \mprj_logic1[111] ;
 wire \mprj_logic1[112] ;
 wire \mprj_logic1[113] ;
 wire \mprj_logic1[114] ;
 wire \mprj_logic1[115] ;
 wire \mprj_logic1[116] ;
 wire \mprj_logic1[117] ;
 wire \mprj_logic1[118] ;
 wire \mprj_logic1[119] ;
 wire \mprj_logic1[11] ;
 wire \mprj_logic1[120] ;
 wire \mprj_logic1[121] ;
 wire \mprj_logic1[122] ;
 wire \mprj_logic1[123] ;
 wire \mprj_logic1[124] ;
 wire \mprj_logic1[125] ;
 wire \mprj_logic1[126] ;
 wire \mprj_logic1[127] ;
 wire \mprj_logic1[128] ;
 wire \mprj_logic1[129] ;
 wire \mprj_logic1[12] ;
 wire \mprj_logic1[130] ;
 wire \mprj_logic1[131] ;
 wire \mprj_logic1[132] ;
 wire \mprj_logic1[133] ;
 wire \mprj_logic1[134] ;
 wire \mprj_logic1[135] ;
 wire \mprj_logic1[136] ;
 wire \mprj_logic1[137] ;
 wire \mprj_logic1[138] ;
 wire \mprj_logic1[139] ;
 wire \mprj_logic1[13] ;
 wire \mprj_logic1[140] ;
 wire \mprj_logic1[141] ;
 wire \mprj_logic1[142] ;
 wire \mprj_logic1[143] ;
 wire \mprj_logic1[144] ;
 wire \mprj_logic1[145] ;
 wire \mprj_logic1[146] ;
 wire \mprj_logic1[147] ;
 wire \mprj_logic1[148] ;
 wire \mprj_logic1[149] ;
 wire \mprj_logic1[14] ;
 wire \mprj_logic1[150] ;
 wire \mprj_logic1[151] ;
 wire \mprj_logic1[152] ;
 wire \mprj_logic1[153] ;
 wire \mprj_logic1[154] ;
 wire \mprj_logic1[155] ;
 wire \mprj_logic1[156] ;
 wire \mprj_logic1[157] ;
 wire \mprj_logic1[158] ;
 wire \mprj_logic1[159] ;
 wire \mprj_logic1[15] ;
 wire \mprj_logic1[160] ;
 wire \mprj_logic1[161] ;
 wire \mprj_logic1[162] ;
 wire \mprj_logic1[163] ;
 wire \mprj_logic1[164] ;
 wire \mprj_logic1[165] ;
 wire \mprj_logic1[166] ;
 wire \mprj_logic1[167] ;
 wire \mprj_logic1[168] ;
 wire \mprj_logic1[169] ;
 wire \mprj_logic1[16] ;
 wire \mprj_logic1[170] ;
 wire \mprj_logic1[171] ;
 wire \mprj_logic1[172] ;
 wire \mprj_logic1[173] ;
 wire \mprj_logic1[174] ;
 wire \mprj_logic1[175] ;
 wire \mprj_logic1[176] ;
 wire \mprj_logic1[177] ;
 wire \mprj_logic1[178] ;
 wire \mprj_logic1[179] ;
 wire \mprj_logic1[17] ;
 wire \mprj_logic1[180] ;
 wire \mprj_logic1[181] ;
 wire \mprj_logic1[182] ;
 wire \mprj_logic1[183] ;
 wire \mprj_logic1[184] ;
 wire \mprj_logic1[185] ;
 wire \mprj_logic1[186] ;
 wire \mprj_logic1[187] ;
 wire \mprj_logic1[188] ;
 wire \mprj_logic1[189] ;
 wire \mprj_logic1[18] ;
 wire \mprj_logic1[190] ;
 wire \mprj_logic1[191] ;
 wire \mprj_logic1[192] ;
 wire \mprj_logic1[193] ;
 wire \mprj_logic1[194] ;
 wire \mprj_logic1[195] ;
 wire \mprj_logic1[196] ;
 wire \mprj_logic1[197] ;
 wire \mprj_logic1[198] ;
 wire \mprj_logic1[199] ;
 wire \mprj_logic1[19] ;
 wire \mprj_logic1[1] ;
 wire \mprj_logic1[200] ;
 wire \mprj_logic1[201] ;
 wire \mprj_logic1[202] ;
 wire \mprj_logic1[203] ;
 wire \mprj_logic1[204] ;
 wire \mprj_logic1[205] ;
 wire \mprj_logic1[206] ;
 wire \mprj_logic1[207] ;
 wire \mprj_logic1[208] ;
 wire \mprj_logic1[209] ;
 wire \mprj_logic1[20] ;
 wire \mprj_logic1[210] ;
 wire \mprj_logic1[211] ;
 wire \mprj_logic1[212] ;
 wire \mprj_logic1[213] ;
 wire \mprj_logic1[214] ;
 wire \mprj_logic1[215] ;
 wire \mprj_logic1[216] ;
 wire \mprj_logic1[217] ;
 wire \mprj_logic1[218] ;
 wire \mprj_logic1[219] ;
 wire \mprj_logic1[21] ;
 wire \mprj_logic1[220] ;
 wire \mprj_logic1[221] ;
 wire \mprj_logic1[222] ;
 wire \mprj_logic1[223] ;
 wire \mprj_logic1[224] ;
 wire \mprj_logic1[225] ;
 wire \mprj_logic1[226] ;
 wire \mprj_logic1[227] ;
 wire \mprj_logic1[228] ;
 wire \mprj_logic1[229] ;
 wire \mprj_logic1[22] ;
 wire \mprj_logic1[230] ;
 wire \mprj_logic1[231] ;
 wire \mprj_logic1[232] ;
 wire \mprj_logic1[233] ;
 wire \mprj_logic1[234] ;
 wire \mprj_logic1[235] ;
 wire \mprj_logic1[236] ;
 wire \mprj_logic1[237] ;
 wire \mprj_logic1[238] ;
 wire \mprj_logic1[239] ;
 wire \mprj_logic1[23] ;
 wire \mprj_logic1[240] ;
 wire \mprj_logic1[241] ;
 wire \mprj_logic1[242] ;
 wire \mprj_logic1[243] ;
 wire \mprj_logic1[244] ;
 wire \mprj_logic1[245] ;
 wire \mprj_logic1[246] ;
 wire \mprj_logic1[247] ;
 wire \mprj_logic1[248] ;
 wire \mprj_logic1[249] ;
 wire \mprj_logic1[24] ;
 wire \mprj_logic1[250] ;
 wire \mprj_logic1[251] ;
 wire \mprj_logic1[252] ;
 wire \mprj_logic1[253] ;
 wire \mprj_logic1[254] ;
 wire \mprj_logic1[255] ;
 wire \mprj_logic1[256] ;
 wire \mprj_logic1[257] ;
 wire \mprj_logic1[258] ;
 wire \mprj_logic1[259] ;
 wire \mprj_logic1[25] ;
 wire \mprj_logic1[260] ;
 wire \mprj_logic1[261] ;
 wire \mprj_logic1[262] ;
 wire \mprj_logic1[263] ;
 wire \mprj_logic1[264] ;
 wire \mprj_logic1[265] ;
 wire \mprj_logic1[266] ;
 wire \mprj_logic1[267] ;
 wire \mprj_logic1[268] ;
 wire \mprj_logic1[269] ;
 wire \mprj_logic1[26] ;
 wire \mprj_logic1[270] ;
 wire \mprj_logic1[271] ;
 wire \mprj_logic1[272] ;
 wire \mprj_logic1[273] ;
 wire \mprj_logic1[274] ;
 wire \mprj_logic1[275] ;
 wire \mprj_logic1[276] ;
 wire \mprj_logic1[277] ;
 wire \mprj_logic1[278] ;
 wire \mprj_logic1[279] ;
 wire \mprj_logic1[27] ;
 wire \mprj_logic1[280] ;
 wire \mprj_logic1[281] ;
 wire \mprj_logic1[282] ;
 wire \mprj_logic1[283] ;
 wire \mprj_logic1[284] ;
 wire \mprj_logic1[285] ;
 wire \mprj_logic1[286] ;
 wire \mprj_logic1[287] ;
 wire \mprj_logic1[288] ;
 wire \mprj_logic1[289] ;
 wire \mprj_logic1[28] ;
 wire \mprj_logic1[290] ;
 wire \mprj_logic1[291] ;
 wire \mprj_logic1[292] ;
 wire \mprj_logic1[293] ;
 wire \mprj_logic1[294] ;
 wire \mprj_logic1[295] ;
 wire \mprj_logic1[296] ;
 wire \mprj_logic1[297] ;
 wire \mprj_logic1[298] ;
 wire \mprj_logic1[299] ;
 wire \mprj_logic1[29] ;
 wire \mprj_logic1[2] ;
 wire \mprj_logic1[300] ;
 wire \mprj_logic1[301] ;
 wire \mprj_logic1[302] ;
 wire \mprj_logic1[303] ;
 wire \mprj_logic1[304] ;
 wire \mprj_logic1[305] ;
 wire \mprj_logic1[306] ;
 wire \mprj_logic1[307] ;
 wire \mprj_logic1[308] ;
 wire \mprj_logic1[309] ;
 wire \mprj_logic1[30] ;
 wire \mprj_logic1[310] ;
 wire \mprj_logic1[311] ;
 wire \mprj_logic1[312] ;
 wire \mprj_logic1[313] ;
 wire \mprj_logic1[314] ;
 wire \mprj_logic1[315] ;
 wire \mprj_logic1[316] ;
 wire \mprj_logic1[317] ;
 wire \mprj_logic1[318] ;
 wire \mprj_logic1[319] ;
 wire \mprj_logic1[31] ;
 wire \mprj_logic1[320] ;
 wire \mprj_logic1[321] ;
 wire \mprj_logic1[322] ;
 wire \mprj_logic1[323] ;
 wire \mprj_logic1[324] ;
 wire \mprj_logic1[325] ;
 wire \mprj_logic1[326] ;
 wire \mprj_logic1[327] ;
 wire \mprj_logic1[328] ;
 wire \mprj_logic1[329] ;
 wire \mprj_logic1[32] ;
 wire \mprj_logic1[330] ;
 wire \mprj_logic1[331] ;
 wire \mprj_logic1[332] ;
 wire \mprj_logic1[333] ;
 wire \mprj_logic1[334] ;
 wire \mprj_logic1[335] ;
 wire \mprj_logic1[336] ;
 wire \mprj_logic1[337] ;
 wire \mprj_logic1[338] ;
 wire \mprj_logic1[339] ;
 wire \mprj_logic1[33] ;
 wire \mprj_logic1[340] ;
 wire \mprj_logic1[341] ;
 wire \mprj_logic1[342] ;
 wire \mprj_logic1[343] ;
 wire \mprj_logic1[344] ;
 wire \mprj_logic1[345] ;
 wire \mprj_logic1[346] ;
 wire \mprj_logic1[347] ;
 wire \mprj_logic1[348] ;
 wire \mprj_logic1[349] ;
 wire \mprj_logic1[34] ;
 wire \mprj_logic1[350] ;
 wire \mprj_logic1[351] ;
 wire \mprj_logic1[352] ;
 wire \mprj_logic1[353] ;
 wire \mprj_logic1[354] ;
 wire \mprj_logic1[355] ;
 wire \mprj_logic1[356] ;
 wire \mprj_logic1[357] ;
 wire \mprj_logic1[358] ;
 wire \mprj_logic1[359] ;
 wire \mprj_logic1[35] ;
 wire \mprj_logic1[360] ;
 wire \mprj_logic1[361] ;
 wire \mprj_logic1[362] ;
 wire \mprj_logic1[363] ;
 wire \mprj_logic1[364] ;
 wire \mprj_logic1[365] ;
 wire \mprj_logic1[366] ;
 wire \mprj_logic1[367] ;
 wire \mprj_logic1[368] ;
 wire \mprj_logic1[369] ;
 wire \mprj_logic1[36] ;
 wire \mprj_logic1[370] ;
 wire \mprj_logic1[371] ;
 wire \mprj_logic1[372] ;
 wire \mprj_logic1[373] ;
 wire \mprj_logic1[374] ;
 wire \mprj_logic1[375] ;
 wire \mprj_logic1[376] ;
 wire \mprj_logic1[377] ;
 wire \mprj_logic1[378] ;
 wire \mprj_logic1[379] ;
 wire \mprj_logic1[37] ;
 wire \mprj_logic1[380] ;
 wire \mprj_logic1[381] ;
 wire \mprj_logic1[382] ;
 wire \mprj_logic1[383] ;
 wire \mprj_logic1[384] ;
 wire \mprj_logic1[385] ;
 wire \mprj_logic1[386] ;
 wire \mprj_logic1[387] ;
 wire \mprj_logic1[388] ;
 wire \mprj_logic1[389] ;
 wire \mprj_logic1[38] ;
 wire \mprj_logic1[390] ;
 wire \mprj_logic1[391] ;
 wire \mprj_logic1[392] ;
 wire \mprj_logic1[393] ;
 wire \mprj_logic1[394] ;
 wire \mprj_logic1[395] ;
 wire \mprj_logic1[396] ;
 wire \mprj_logic1[397] ;
 wire \mprj_logic1[398] ;
 wire \mprj_logic1[399] ;
 wire \mprj_logic1[39] ;
 wire \mprj_logic1[3] ;
 wire \mprj_logic1[400] ;
 wire \mprj_logic1[401] ;
 wire \mprj_logic1[402] ;
 wire \mprj_logic1[403] ;
 wire \mprj_logic1[404] ;
 wire \mprj_logic1[405] ;
 wire \mprj_logic1[406] ;
 wire \mprj_logic1[407] ;
 wire \mprj_logic1[408] ;
 wire \mprj_logic1[409] ;
 wire \mprj_logic1[40] ;
 wire \mprj_logic1[410] ;
 wire \mprj_logic1[411] ;
 wire \mprj_logic1[412] ;
 wire \mprj_logic1[413] ;
 wire \mprj_logic1[414] ;
 wire \mprj_logic1[415] ;
 wire \mprj_logic1[416] ;
 wire \mprj_logic1[417] ;
 wire \mprj_logic1[418] ;
 wire \mprj_logic1[419] ;
 wire \mprj_logic1[41] ;
 wire \mprj_logic1[420] ;
 wire \mprj_logic1[421] ;
 wire \mprj_logic1[422] ;
 wire \mprj_logic1[423] ;
 wire \mprj_logic1[424] ;
 wire \mprj_logic1[425] ;
 wire \mprj_logic1[426] ;
 wire \mprj_logic1[427] ;
 wire \mprj_logic1[428] ;
 wire \mprj_logic1[429] ;
 wire \mprj_logic1[42] ;
 wire \mprj_logic1[430] ;
 wire \mprj_logic1[431] ;
 wire \mprj_logic1[432] ;
 wire \mprj_logic1[433] ;
 wire \mprj_logic1[434] ;
 wire \mprj_logic1[435] ;
 wire \mprj_logic1[436] ;
 wire \mprj_logic1[437] ;
 wire \mprj_logic1[438] ;
 wire \mprj_logic1[439] ;
 wire \mprj_logic1[43] ;
 wire \mprj_logic1[440] ;
 wire \mprj_logic1[441] ;
 wire \mprj_logic1[442] ;
 wire \mprj_logic1[443] ;
 wire \mprj_logic1[444] ;
 wire \mprj_logic1[445] ;
 wire \mprj_logic1[446] ;
 wire \mprj_logic1[447] ;
 wire \mprj_logic1[448] ;
 wire \mprj_logic1[449] ;
 wire \mprj_logic1[44] ;
 wire \mprj_logic1[450] ;
 wire \mprj_logic1[451] ;
 wire \mprj_logic1[452] ;
 wire \mprj_logic1[453] ;
 wire \mprj_logic1[454] ;
 wire \mprj_logic1[455] ;
 wire \mprj_logic1[456] ;
 wire \mprj_logic1[457] ;
 wire \mprj_logic1[458] ;
 wire \mprj_logic1[459] ;
 wire \mprj_logic1[45] ;
 wire \mprj_logic1[460] ;
 wire \mprj_logic1[462] ;
 wire \mprj_logic1[46] ;
 wire \mprj_logic1[47] ;
 wire \mprj_logic1[48] ;
 wire \mprj_logic1[49] ;
 wire \mprj_logic1[4] ;
 wire \mprj_logic1[50] ;
 wire \mprj_logic1[51] ;
 wire \mprj_logic1[52] ;
 wire \mprj_logic1[53] ;
 wire \mprj_logic1[54] ;
 wire \mprj_logic1[55] ;
 wire \mprj_logic1[56] ;
 wire \mprj_logic1[57] ;
 wire \mprj_logic1[58] ;
 wire \mprj_logic1[59] ;
 wire \mprj_logic1[5] ;
 wire \mprj_logic1[60] ;
 wire \mprj_logic1[61] ;
 wire \mprj_logic1[62] ;
 wire \mprj_logic1[63] ;
 wire \mprj_logic1[64] ;
 wire \mprj_logic1[65] ;
 wire \mprj_logic1[66] ;
 wire \mprj_logic1[67] ;
 wire \mprj_logic1[68] ;
 wire \mprj_logic1[69] ;
 wire \mprj_logic1[6] ;
 wire \mprj_logic1[70] ;
 wire \mprj_logic1[71] ;
 wire \mprj_logic1[72] ;
 wire \mprj_logic1[73] ;
 wire \mprj_logic1[74] ;
 wire \mprj_logic1[75] ;
 wire \mprj_logic1[76] ;
 wire \mprj_logic1[77] ;
 wire \mprj_logic1[78] ;
 wire \mprj_logic1[79] ;
 wire \mprj_logic1[7] ;
 wire \mprj_logic1[80] ;
 wire \mprj_logic1[81] ;
 wire \mprj_logic1[82] ;
 wire \mprj_logic1[83] ;
 wire \mprj_logic1[84] ;
 wire \mprj_logic1[85] ;
 wire \mprj_logic1[86] ;
 wire \mprj_logic1[87] ;
 wire \mprj_logic1[88] ;
 wire \mprj_logic1[89] ;
 wire \mprj_logic1[8] ;
 wire \mprj_logic1[90] ;
 wire \mprj_logic1[91] ;
 wire \mprj_logic1[92] ;
 wire \mprj_logic1[93] ;
 wire \mprj_logic1[94] ;
 wire \mprj_logic1[95] ;
 wire \mprj_logic1[96] ;
 wire \mprj_logic1[97] ;
 wire \mprj_logic1[98] ;
 wire \mprj_logic1[99] ;
 wire \mprj_logic1[9] ;
 wire \user_irq_bar[0] ;
 wire \user_irq_bar[1] ;
 wire \user_irq_bar[2] ;
 wire \user_irq_enable[0] ;
 wire \user_irq_enable[1] ;
 wire \user_irq_enable[2] ;
 wire wb_in_enable;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;

 sky130_fd_sc_hd__inv_2 _0462_ (.A(\la_data_in_mprj_bar[17] ),
    .Y(net627));
 sky130_fd_sc_hd__clkinv_2 _0463_ (.A(\la_data_in_mprj_bar[18] ),
    .Y(net628));
 sky130_fd_sc_hd__inv_2 _0464_ (.A(\la_data_in_mprj_bar[19] ),
    .Y(net629));
 sky130_fd_sc_hd__inv_2 _0465_ (.A(\la_data_in_mprj_bar[20] ),
    .Y(net631));
 sky130_fd_sc_hd__inv_2 _0466_ (.A(\la_data_in_mprj_bar[21] ),
    .Y(net632));
 sky130_fd_sc_hd__clkinv_2 _0467_ (.A(\la_data_in_mprj_bar[22] ),
    .Y(net633));
 sky130_fd_sc_hd__inv_2 _0468_ (.A(\la_data_in_mprj_bar[23] ),
    .Y(net634));
 sky130_fd_sc_hd__clkinv_2 _0469_ (.A(\la_data_in_mprj_bar[24] ),
    .Y(net635));
 sky130_fd_sc_hd__inv_2 _0470_ (.A(\la_data_in_mprj_bar[25] ),
    .Y(net636));
 sky130_fd_sc_hd__inv_2 _0471_ (.A(\la_data_in_mprj_bar[26] ),
    .Y(net637));
 sky130_fd_sc_hd__clkinv_2 _0472_ (.A(\la_data_in_mprj_bar[27] ),
    .Y(net638));
 sky130_fd_sc_hd__inv_2 _0473_ (.A(\la_data_in_mprj_bar[28] ),
    .Y(net639));
 sky130_fd_sc_hd__inv_2 _0474_ (.A(\la_data_in_mprj_bar[29] ),
    .Y(net640));
 sky130_fd_sc_hd__inv_2 _0475_ (.A(\la_data_in_mprj_bar[30] ),
    .Y(net642));
 sky130_fd_sc_hd__inv_1 _0476_ (.A(\la_data_in_mprj_bar[31] ),
    .Y(net643));
 sky130_fd_sc_hd__clkinv_2 _0477_ (.A(\la_data_in_mprj_bar[32] ),
    .Y(net644));
 sky130_fd_sc_hd__inv_2 _0478_ (.A(\la_data_in_mprj_bar[33] ),
    .Y(net645));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\la_data_in_mprj_bar[34] ),
    .Y(net646));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(\la_data_in_mprj_bar[35] ),
    .Y(net647));
 sky130_fd_sc_hd__clkinv_2 _0481_ (.A(\la_data_in_mprj_bar[36] ),
    .Y(net648));
 sky130_fd_sc_hd__inv_2 _0482_ (.A(\la_data_in_mprj_bar[37] ),
    .Y(net649));
 sky130_fd_sc_hd__inv_2 _0483_ (.A(\la_data_in_mprj_bar[38] ),
    .Y(net650));
 sky130_fd_sc_hd__clkinv_2 _0484_ (.A(\la_data_in_mprj_bar[39] ),
    .Y(net651));
 sky130_fd_sc_hd__inv_2 _0485_ (.A(\la_data_in_mprj_bar[40] ),
    .Y(net653));
 sky130_fd_sc_hd__clkinv_2 _0486_ (.A(\la_data_in_mprj_bar[41] ),
    .Y(net654));
 sky130_fd_sc_hd__inv_2 _0487_ (.A(\la_data_in_mprj_bar[42] ),
    .Y(net655));
 sky130_fd_sc_hd__clkinv_2 _0488_ (.A(\la_data_in_mprj_bar[43] ),
    .Y(net656));
 sky130_fd_sc_hd__clkinv_2 _0489_ (.A(\la_data_in_mprj_bar[44] ),
    .Y(net657));
 sky130_fd_sc_hd__inv_2 _0490_ (.A(\la_data_in_mprj_bar[45] ),
    .Y(net658));
 sky130_fd_sc_hd__clkinv_2 _0491_ (.A(\la_data_in_mprj_bar[46] ),
    .Y(net659));
 sky130_fd_sc_hd__inv_2 _0492_ (.A(\la_data_in_mprj_bar[47] ),
    .Y(net660));
 sky130_fd_sc_hd__clkinv_2 _0493_ (.A(\la_data_in_mprj_bar[48] ),
    .Y(net661));
 sky130_fd_sc_hd__inv_2 _0494_ (.A(\la_data_in_mprj_bar[49] ),
    .Y(net662));
 sky130_fd_sc_hd__clkinv_2 _0495_ (.A(\la_data_in_mprj_bar[50] ),
    .Y(net664));
 sky130_fd_sc_hd__inv_2 _0496_ (.A(\la_data_in_mprj_bar[51] ),
    .Y(net665));
 sky130_fd_sc_hd__inv_1 _0497_ (.A(\la_data_in_mprj_bar[52] ),
    .Y(net666));
 sky130_fd_sc_hd__clkinv_2 _0498_ (.A(\la_data_in_mprj_bar[53] ),
    .Y(net667));
 sky130_fd_sc_hd__clkinv_2 _0499_ (.A(\la_data_in_mprj_bar[54] ),
    .Y(net668));
 sky130_fd_sc_hd__inv_2 _0500_ (.A(\la_data_in_mprj_bar[55] ),
    .Y(net669));
 sky130_fd_sc_hd__inv_2 _0501_ (.A(\la_data_in_mprj_bar[56] ),
    .Y(net670));
 sky130_fd_sc_hd__inv_2 _0502_ (.A(\la_data_in_mprj_bar[57] ),
    .Y(net671));
 sky130_fd_sc_hd__inv_2 _0503_ (.A(\la_data_in_mprj_bar[58] ),
    .Y(net672));
 sky130_fd_sc_hd__inv_2 _0504_ (.A(\la_data_in_mprj_bar[59] ),
    .Y(net673));
 sky130_fd_sc_hd__inv_2 _0505_ (.A(\la_data_in_mprj_bar[60] ),
    .Y(net675));
 sky130_fd_sc_hd__inv_2 _0506_ (.A(\la_data_in_mprj_bar[61] ),
    .Y(net676));
 sky130_fd_sc_hd__inv_2 _0507_ (.A(\la_data_in_mprj_bar[62] ),
    .Y(net677));
 sky130_fd_sc_hd__inv_2 _0508_ (.A(\la_data_in_mprj_bar[63] ),
    .Y(net678));
 sky130_fd_sc_hd__inv_2 _0509_ (.A(\la_data_in_mprj_bar[64] ),
    .Y(net679));
 sky130_fd_sc_hd__inv_2 _0510_ (.A(\la_data_in_mprj_bar[65] ),
    .Y(net680));
 sky130_fd_sc_hd__inv_2 _0511_ (.A(\la_data_in_mprj_bar[66] ),
    .Y(net681));
 sky130_fd_sc_hd__inv_2 _0512_ (.A(\la_data_in_mprj_bar[67] ),
    .Y(net682));
 sky130_fd_sc_hd__inv_2 _0513_ (.A(\la_data_in_mprj_bar[68] ),
    .Y(net683));
 sky130_fd_sc_hd__inv_2 _0514_ (.A(\la_data_in_mprj_bar[69] ),
    .Y(net684));
 sky130_fd_sc_hd__inv_2 _0515_ (.A(net1080),
    .Y(net686));
 sky130_fd_sc_hd__inv_2 _0516_ (.A(net1079),
    .Y(net687));
 sky130_fd_sc_hd__inv_2 _0517_ (.A(net1077),
    .Y(net688));
 sky130_fd_sc_hd__clkinv_2 _0518_ (.A(net1075),
    .Y(net689));
 sky130_fd_sc_hd__inv_2 _0519_ (.A(net1073),
    .Y(net690));
 sky130_fd_sc_hd__inv_2 _0520_ (.A(net1070),
    .Y(net691));
 sky130_fd_sc_hd__inv_2 _0521_ (.A(net1067),
    .Y(net692));
 sky130_fd_sc_hd__inv_2 _0522_ (.A(net1063),
    .Y(net693));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(net1061),
    .Y(net694));
 sky130_fd_sc_hd__inv_2 _0524_ (.A(net1059),
    .Y(net695));
 sky130_fd_sc_hd__inv_2 _0525_ (.A(net1056),
    .Y(net697));
 sky130_fd_sc_hd__inv_2 _0526_ (.A(net1053),
    .Y(net698));
 sky130_fd_sc_hd__inv_2 _0527_ (.A(net1051),
    .Y(net699));
 sky130_fd_sc_hd__inv_2 _0528_ (.A(net1049),
    .Y(net700));
 sky130_fd_sc_hd__inv_2 _0529_ (.A(net1046),
    .Y(net701));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(net1044),
    .Y(net702));
 sky130_fd_sc_hd__clkinv_2 _0531_ (.A(net1042),
    .Y(net703));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(net1039),
    .Y(net704));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(net1036),
    .Y(net705));
 sky130_fd_sc_hd__clkinv_2 _0534_ (.A(net1035),
    .Y(net706));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(net1032),
    .Y(net708));
 sky130_fd_sc_hd__clkinv_2 _0536_ (.A(net1030),
    .Y(net709));
 sky130_fd_sc_hd__inv_2 _0537_ (.A(net1028),
    .Y(net710));
 sky130_fd_sc_hd__inv_2 _0538_ (.A(net1026),
    .Y(net711));
 sky130_fd_sc_hd__inv_2 _0539_ (.A(net1024),
    .Y(net712));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(net1021),
    .Y(net713));
 sky130_fd_sc_hd__inv_2 _0541_ (.A(net1019),
    .Y(net714));
 sky130_fd_sc_hd__inv_2 _0542_ (.A(net1017),
    .Y(net715));
 sky130_fd_sc_hd__inv_2 _0543_ (.A(net1015),
    .Y(net716));
 sky130_fd_sc_hd__inv_2 _0544_ (.A(net1013),
    .Y(net717));
 sky130_fd_sc_hd__inv_2 _0545_ (.A(net1086),
    .Y(net592));
 sky130_fd_sc_hd__inv_2 _0546_ (.A(net1084),
    .Y(net593));
 sky130_fd_sc_hd__inv_2 _0547_ (.A(net1083),
    .Y(net594));
 sky130_fd_sc_hd__inv_2 _0548_ (.A(net1081),
    .Y(net595));
 sky130_fd_sc_hd__clkinv_4 _0549_ (.A(\la_data_in_mprj_bar[104] ),
    .Y(net596));
 sky130_fd_sc_hd__clkinv_2 _0550_ (.A(\la_data_in_mprj_bar[105] ),
    .Y(net597));
 sky130_fd_sc_hd__clkinv_4 _0551_ (.A(\la_data_in_mprj_bar[106] ),
    .Y(net598));
 sky130_fd_sc_hd__inv_2 _0552_ (.A(\la_data_in_mprj_bar[107] ),
    .Y(net599));
 sky130_fd_sc_hd__inv_2 _0553_ (.A(\la_data_in_mprj_bar[108] ),
    .Y(net600));
 sky130_fd_sc_hd__clkinv_4 _0554_ (.A(\la_data_in_mprj_bar[109] ),
    .Y(net601));
 sky130_fd_sc_hd__clkinv_4 _0555_ (.A(\la_data_in_mprj_bar[110] ),
    .Y(net603));
 sky130_fd_sc_hd__clkinv_4 _0556_ (.A(\la_data_in_mprj_bar[111] ),
    .Y(net604));
 sky130_fd_sc_hd__clkinv_4 _0557_ (.A(\la_data_in_mprj_bar[112] ),
    .Y(net605));
 sky130_fd_sc_hd__clkinv_4 _0558_ (.A(\la_data_in_mprj_bar[113] ),
    .Y(net606));
 sky130_fd_sc_hd__clkinv_4 _0559_ (.A(\la_data_in_mprj_bar[114] ),
    .Y(net607));
 sky130_fd_sc_hd__clkinv_4 _0560_ (.A(\la_data_in_mprj_bar[115] ),
    .Y(net608));
 sky130_fd_sc_hd__clkinv_4 _0561_ (.A(\la_data_in_mprj_bar[116] ),
    .Y(net609));
 sky130_fd_sc_hd__clkinv_4 _0562_ (.A(\la_data_in_mprj_bar[117] ),
    .Y(net610));
 sky130_fd_sc_hd__inv_2 _0563_ (.A(\la_data_in_mprj_bar[118] ),
    .Y(net611));
 sky130_fd_sc_hd__clkinv_2 _0564_ (.A(\la_data_in_mprj_bar[119] ),
    .Y(net612));
 sky130_fd_sc_hd__clkinv_4 _0565_ (.A(\la_data_in_mprj_bar[120] ),
    .Y(net614));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(\la_data_in_mprj_bar[121] ),
    .Y(net615));
 sky130_fd_sc_hd__inv_2 _0567_ (.A(\la_data_in_mprj_bar[122] ),
    .Y(net616));
 sky130_fd_sc_hd__inv_2 _0568_ (.A(\la_data_in_mprj_bar[123] ),
    .Y(net617));
 sky130_fd_sc_hd__clkinv_2 _0569_ (.A(\la_data_in_mprj_bar[124] ),
    .Y(net618));
 sky130_fd_sc_hd__inv_2 _0570_ (.A(\la_data_in_mprj_bar[125] ),
    .Y(net619));
 sky130_fd_sc_hd__clkinv_2 _0571_ (.A(\la_data_in_mprj_bar[126] ),
    .Y(net620));
 sky130_fd_sc_hd__clkinv_2 _0572_ (.A(\la_data_in_mprj_bar[127] ),
    .Y(net621));
 sky130_fd_sc_hd__inv_2 _0573_ (.A(\user_irq_bar[0] ),
    .Y(net957));
 sky130_fd_sc_hd__inv_2 _0574_ (.A(\user_irq_bar[1] ),
    .Y(net958));
 sky130_fd_sc_hd__inv_2 _0575_ (.A(\user_irq_bar[2] ),
    .Y(net959));
 sky130_fd_sc_hd__clkinv_2 _0576_ (.A(\mprj_dat_i_core_bar[0] ),
    .Y(net881));
 sky130_fd_sc_hd__clkinv_2 _0577_ (.A(\mprj_dat_i_core_bar[1] ),
    .Y(net892));
 sky130_fd_sc_hd__inv_2 _0578_ (.A(\mprj_dat_i_core_bar[2] ),
    .Y(net903));
 sky130_fd_sc_hd__inv_2 _0579_ (.A(\mprj_dat_i_core_bar[3] ),
    .Y(net906));
 sky130_fd_sc_hd__inv_2 _0580_ (.A(\mprj_dat_i_core_bar[4] ),
    .Y(net907));
 sky130_fd_sc_hd__clkinv_2 _0581_ (.A(\mprj_dat_i_core_bar[5] ),
    .Y(net908));
 sky130_fd_sc_hd__clkinv_2 _0582_ (.A(\mprj_dat_i_core_bar[6] ),
    .Y(net909));
 sky130_fd_sc_hd__inv_2 _0583_ (.A(\mprj_dat_i_core_bar[7] ),
    .Y(net910));
 sky130_fd_sc_hd__clkinv_2 _0584_ (.A(\mprj_dat_i_core_bar[8] ),
    .Y(net911));
 sky130_fd_sc_hd__inv_2 _0585_ (.A(\mprj_dat_i_core_bar[9] ),
    .Y(net912));
 sky130_fd_sc_hd__inv_2 _0586_ (.A(\mprj_dat_i_core_bar[10] ),
    .Y(net882));
 sky130_fd_sc_hd__inv_2 _0587_ (.A(\mprj_dat_i_core_bar[11] ),
    .Y(net883));
 sky130_fd_sc_hd__clkinv_2 _0588_ (.A(\mprj_dat_i_core_bar[12] ),
    .Y(net884));
 sky130_fd_sc_hd__inv_2 _0589_ (.A(\mprj_dat_i_core_bar[13] ),
    .Y(net885));
 sky130_fd_sc_hd__inv_2 _0590_ (.A(\mprj_dat_i_core_bar[14] ),
    .Y(net886));
 sky130_fd_sc_hd__inv_2 _0591_ (.A(\mprj_dat_i_core_bar[15] ),
    .Y(net887));
 sky130_fd_sc_hd__inv_2 _0592_ (.A(\mprj_dat_i_core_bar[16] ),
    .Y(net888));
 sky130_fd_sc_hd__inv_2 _0593_ (.A(\mprj_dat_i_core_bar[17] ),
    .Y(net889));
 sky130_fd_sc_hd__inv_2 _0594_ (.A(\mprj_dat_i_core_bar[18] ),
    .Y(net890));
 sky130_fd_sc_hd__inv_2 _0595_ (.A(\mprj_dat_i_core_bar[19] ),
    .Y(net891));
 sky130_fd_sc_hd__inv_2 _0596_ (.A(\mprj_dat_i_core_bar[20] ),
    .Y(net893));
 sky130_fd_sc_hd__inv_2 _0597_ (.A(\mprj_dat_i_core_bar[21] ),
    .Y(net894));
 sky130_fd_sc_hd__inv_2 _0598_ (.A(\mprj_dat_i_core_bar[22] ),
    .Y(net895));
 sky130_fd_sc_hd__inv_2 _0599_ (.A(\mprj_dat_i_core_bar[23] ),
    .Y(net896));
 sky130_fd_sc_hd__inv_2 _0600_ (.A(\mprj_dat_i_core_bar[24] ),
    .Y(net897));
 sky130_fd_sc_hd__inv_2 _0601_ (.A(\mprj_dat_i_core_bar[25] ),
    .Y(net898));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\mprj_dat_i_core_bar[26] ),
    .Y(net899));
 sky130_fd_sc_hd__inv_2 _0603_ (.A(\mprj_dat_i_core_bar[27] ),
    .Y(net900));
 sky130_fd_sc_hd__inv_2 _0604_ (.A(\mprj_dat_i_core_bar[28] ),
    .Y(net901));
 sky130_fd_sc_hd__inv_2 _0605_ (.A(\mprj_dat_i_core_bar[29] ),
    .Y(net902));
 sky130_fd_sc_hd__inv_2 _0606_ (.A(\mprj_dat_i_core_bar[30] ),
    .Y(net904));
 sky130_fd_sc_hd__inv_2 _0607_ (.A(\mprj_dat_i_core_bar[31] ),
    .Y(net905));
 sky130_fd_sc_hd__clkinv_2 _0608_ (.A(mprj_ack_i_core_bar),
    .Y(net847));
 sky130_fd_sc_hd__and2_1 _0609_ (.A(net2417),
    .B(net171),
    .X(_0000_));
 sky130_fd_sc_hd__clkbuf_1 _0610_ (.A(_0000_),
    .X(\la_data_in_enable[1] ));
 sky130_fd_sc_hd__and2_1 _0611_ (.A(net2415),
    .B(net182),
    .X(_0001_));
 sky130_fd_sc_hd__clkbuf_1 _0612_ (.A(_0001_),
    .X(\la_data_in_enable[2] ));
 sky130_fd_sc_hd__and2_1 _0613_ (.A(net2413),
    .B(net193),
    .X(_0002_));
 sky130_fd_sc_hd__clkbuf_1 _0614_ (.A(_0002_),
    .X(\la_data_in_enable[3] ));
 sky130_fd_sc_hd__and2_1 _0615_ (.A(net2410),
    .B(net204),
    .X(_0003_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0003_),
    .X(\la_data_in_enable[4] ));
 sky130_fd_sc_hd__and2_1 _0617_ (.A(net2408),
    .B(net215),
    .X(_0004_));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(_0004_),
    .X(\la_data_in_enable[5] ));
 sky130_fd_sc_hd__and2_1 _0619_ (.A(net2407),
    .B(net226),
    .X(_0005_));
 sky130_fd_sc_hd__clkbuf_1 _0620_ (.A(_0005_),
    .X(\la_data_in_enable[6] ));
 sky130_fd_sc_hd__and2_1 _0621_ (.A(net2405),
    .B(net237),
    .X(_0006_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0006_),
    .X(\la_data_in_enable[7] ));
 sky130_fd_sc_hd__and2_1 _0623_ (.A(net2404),
    .B(net248),
    .X(_0007_));
 sky130_fd_sc_hd__clkbuf_1 _0624_ (.A(_0007_),
    .X(\la_data_in_enable[8] ));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(net2403),
    .B(net1974),
    .X(_0008_));
 sky130_fd_sc_hd__clkbuf_1 _0626_ (.A(_0008_),
    .X(\la_data_in_enable[9] ));
 sky130_fd_sc_hd__and2_1 _0627_ (.A(net2402),
    .B(net2024),
    .X(_0009_));
 sky130_fd_sc_hd__clkbuf_1 _0628_ (.A(_0009_),
    .X(\la_data_in_enable[10] ));
 sky130_fd_sc_hd__and2_1 _0629_ (.A(net2399),
    .B(net154),
    .X(_0010_));
 sky130_fd_sc_hd__clkbuf_1 _0630_ (.A(_0010_),
    .X(\la_data_in_enable[11] ));
 sky130_fd_sc_hd__and2_1 _0631_ (.A(net2396),
    .B(net163),
    .X(_0011_));
 sky130_fd_sc_hd__clkbuf_1 _0632_ (.A(_0011_),
    .X(\la_data_in_enable[12] ));
 sky130_fd_sc_hd__and2_1 _0633_ (.A(net2392),
    .B(net164),
    .X(_0012_));
 sky130_fd_sc_hd__clkbuf_1 _0634_ (.A(_0012_),
    .X(\la_data_in_enable[13] ));
 sky130_fd_sc_hd__and2_1 _0635_ (.A(net2390),
    .B(net165),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_1 _0636_ (.A(_0013_),
    .X(\la_data_in_enable[14] ));
 sky130_fd_sc_hd__and2_1 _0637_ (.A(net2388),
    .B(net166),
    .X(_0014_));
 sky130_fd_sc_hd__clkbuf_1 _0638_ (.A(_0014_),
    .X(\la_data_in_enable[15] ));
 sky130_fd_sc_hd__and2_1 _0639_ (.A(net2386),
    .B(net167),
    .X(_0015_));
 sky130_fd_sc_hd__clkbuf_1 _0640_ (.A(_0015_),
    .X(\la_data_in_enable[16] ));
 sky130_fd_sc_hd__and2_1 _0641_ (.A(net2384),
    .B(net168),
    .X(_0016_));
 sky130_fd_sc_hd__clkbuf_1 _0642_ (.A(_0016_),
    .X(\la_data_in_enable[17] ));
 sky130_fd_sc_hd__and2_1 _0643_ (.A(net2382),
    .B(net169),
    .X(_0017_));
 sky130_fd_sc_hd__clkbuf_1 _0644_ (.A(_0017_),
    .X(\la_data_in_enable[18] ));
 sky130_fd_sc_hd__and2_1 _0645_ (.A(net2380),
    .B(net170),
    .X(_0018_));
 sky130_fd_sc_hd__clkbuf_1 _0646_ (.A(_0018_),
    .X(\la_data_in_enable[19] ));
 sky130_fd_sc_hd__and2_1 _0647_ (.A(net2378),
    .B(net172),
    .X(_0019_));
 sky130_fd_sc_hd__clkbuf_1 _0648_ (.A(_0019_),
    .X(\la_data_in_enable[20] ));
 sky130_fd_sc_hd__and2_1 _0649_ (.A(net2377),
    .B(net173),
    .X(_0020_));
 sky130_fd_sc_hd__clkbuf_1 _0650_ (.A(_0020_),
    .X(\la_data_in_enable[21] ));
 sky130_fd_sc_hd__and2_1 _0651_ (.A(net2375),
    .B(net174),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_1 _0652_ (.A(_0021_),
    .X(\la_data_in_enable[22] ));
 sky130_fd_sc_hd__and2_1 _0653_ (.A(net2372),
    .B(net2006),
    .X(_0022_));
 sky130_fd_sc_hd__clkbuf_1 _0654_ (.A(_0022_),
    .X(\la_data_in_enable[23] ));
 sky130_fd_sc_hd__and2_1 _0655_ (.A(net2370),
    .B(net176),
    .X(_0023_));
 sky130_fd_sc_hd__clkbuf_1 _0656_ (.A(_0023_),
    .X(\la_data_in_enable[24] ));
 sky130_fd_sc_hd__and2_1 _0657_ (.A(net2368),
    .B(net177),
    .X(_0024_));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(_0024_),
    .X(\la_data_in_enable[25] ));
 sky130_fd_sc_hd__and2_1 _0659_ (.A(net2366),
    .B(net178),
    .X(_0025_));
 sky130_fd_sc_hd__clkbuf_1 _0660_ (.A(_0025_),
    .X(\la_data_in_enable[26] ));
 sky130_fd_sc_hd__and2_1 _0661_ (.A(net2365),
    .B(net179),
    .X(_0026_));
 sky130_fd_sc_hd__clkbuf_1 _0662_ (.A(_0026_),
    .X(\la_data_in_enable[27] ));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(net2363),
    .B(net2005),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_1 _0664_ (.A(_0027_),
    .X(\la_data_in_enable[28] ));
 sky130_fd_sc_hd__and2_1 _0665_ (.A(net2361),
    .B(net181),
    .X(_0028_));
 sky130_fd_sc_hd__clkbuf_1 _0666_ (.A(_0028_),
    .X(\la_data_in_enable[29] ));
 sky130_fd_sc_hd__and2_1 _0667_ (.A(net2359),
    .B(net183),
    .X(_0029_));
 sky130_fd_sc_hd__clkbuf_1 _0668_ (.A(_0029_),
    .X(\la_data_in_enable[30] ));
 sky130_fd_sc_hd__and2_1 _0669_ (.A(net2358),
    .B(net184),
    .X(_0030_));
 sky130_fd_sc_hd__clkbuf_1 _0670_ (.A(_0030_),
    .X(\la_data_in_enable[31] ));
 sky130_fd_sc_hd__and2_1 _0671_ (.A(net2357),
    .B(net185),
    .X(_0031_));
 sky130_fd_sc_hd__clkbuf_1 _0672_ (.A(net1632),
    .X(\la_data_in_enable[32] ));
 sky130_fd_sc_hd__and2_1 _0673_ (.A(net2355),
    .B(net186),
    .X(_0032_));
 sky130_fd_sc_hd__clkbuf_1 _0674_ (.A(_0032_),
    .X(\la_data_in_enable[33] ));
 sky130_fd_sc_hd__and2_1 _0675_ (.A(net2354),
    .B(net187),
    .X(_0033_));
 sky130_fd_sc_hd__clkbuf_1 _0676_ (.A(_0033_),
    .X(\la_data_in_enable[34] ));
 sky130_fd_sc_hd__and2_1 _0677_ (.A(net2352),
    .B(net2004),
    .X(_0034_));
 sky130_fd_sc_hd__clkbuf_1 _0678_ (.A(_0034_),
    .X(\la_data_in_enable[35] ));
 sky130_fd_sc_hd__and2_1 _0679_ (.A(net2351),
    .B(net189),
    .X(_0035_));
 sky130_fd_sc_hd__clkbuf_1 _0680_ (.A(_0035_),
    .X(\la_data_in_enable[36] ));
 sky130_fd_sc_hd__and2_1 _0681_ (.A(\mprj_logic1[367] ),
    .B(net190),
    .X(_0036_));
 sky130_fd_sc_hd__clkbuf_1 _0682_ (.A(net1631),
    .X(\la_data_in_enable[37] ));
 sky130_fd_sc_hd__and2_1 _0683_ (.A(net2349),
    .B(net2003),
    .X(_0037_));
 sky130_fd_sc_hd__clkbuf_1 _0684_ (.A(_0037_),
    .X(\la_data_in_enable[38] ));
 sky130_fd_sc_hd__and2_1 _0685_ (.A(net2348),
    .B(net192),
    .X(_0038_));
 sky130_fd_sc_hd__clkbuf_1 _0686_ (.A(_0038_),
    .X(\la_data_in_enable[39] ));
 sky130_fd_sc_hd__and2_1 _0687_ (.A(net2347),
    .B(net194),
    .X(_0039_));
 sky130_fd_sc_hd__clkbuf_1 _0688_ (.A(_0039_),
    .X(\la_data_in_enable[40] ));
 sky130_fd_sc_hd__and2_1 _0689_ (.A(net2346),
    .B(net2002),
    .X(_0040_));
 sky130_fd_sc_hd__clkbuf_1 _0690_ (.A(_0040_),
    .X(\la_data_in_enable[41] ));
 sky130_fd_sc_hd__and2_1 _0691_ (.A(net2345),
    .B(net196),
    .X(_0041_));
 sky130_fd_sc_hd__clkbuf_1 _0692_ (.A(_0041_),
    .X(\la_data_in_enable[42] ));
 sky130_fd_sc_hd__and2_1 _0693_ (.A(net2344),
    .B(net2001),
    .X(_0042_));
 sky130_fd_sc_hd__clkbuf_1 _0694_ (.A(_0042_),
    .X(\la_data_in_enable[43] ));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(net2343),
    .B(net198),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_1 _0696_ (.A(_0043_),
    .X(\la_data_in_enable[44] ));
 sky130_fd_sc_hd__and2_1 _0697_ (.A(net2342),
    .B(net2000),
    .X(_0044_));
 sky130_fd_sc_hd__clkbuf_1 _0698_ (.A(_0044_),
    .X(\la_data_in_enable[45] ));
 sky130_fd_sc_hd__and2_1 _0699_ (.A(net2341),
    .B(net200),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_1 _0700_ (.A(_0045_),
    .X(\la_data_in_enable[46] ));
 sky130_fd_sc_hd__and2_1 _0701_ (.A(net2340),
    .B(net1999),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_1 _0702_ (.A(_0046_),
    .X(\la_data_in_enable[47] ));
 sky130_fd_sc_hd__and2_1 _0703_ (.A(net2339),
    .B(net1998),
    .X(_0047_));
 sky130_fd_sc_hd__clkbuf_1 _0704_ (.A(_0047_),
    .X(\la_data_in_enable[48] ));
 sky130_fd_sc_hd__and2_1 _0705_ (.A(\mprj_logic1[379] ),
    .B(net203),
    .X(_0048_));
 sky130_fd_sc_hd__clkbuf_1 _0706_ (.A(_0048_),
    .X(\la_data_in_enable[49] ));
 sky130_fd_sc_hd__and2_1 _0707_ (.A(net2338),
    .B(net1997),
    .X(_0049_));
 sky130_fd_sc_hd__clkbuf_1 _0708_ (.A(_0049_),
    .X(\la_data_in_enable[50] ));
 sky130_fd_sc_hd__and2_1 _0709_ (.A(net2337),
    .B(net1996),
    .X(_0050_));
 sky130_fd_sc_hd__clkbuf_1 _0710_ (.A(_0050_),
    .X(\la_data_in_enable[51] ));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(net2336),
    .B(net207),
    .X(_0051_));
 sky130_fd_sc_hd__clkbuf_1 _0712_ (.A(_0051_),
    .X(\la_data_in_enable[52] ));
 sky130_fd_sc_hd__and2_1 _0713_ (.A(net2335),
    .B(net1995),
    .X(_0052_));
 sky130_fd_sc_hd__clkbuf_1 _0714_ (.A(_0052_),
    .X(\la_data_in_enable[53] ));
 sky130_fd_sc_hd__and2_1 _0715_ (.A(net2334),
    .B(net1994),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_1 _0716_ (.A(_0053_),
    .X(\la_data_in_enable[54] ));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(\mprj_logic1[385] ),
    .B(net210),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_1 _0718_ (.A(_0054_),
    .X(\la_data_in_enable[55] ));
 sky130_fd_sc_hd__and2_1 _0719_ (.A(net2333),
    .B(net211),
    .X(_0055_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0720_ (.A(_0055_),
    .X(\la_data_in_enable[56] ));
 sky130_fd_sc_hd__and2_1 _0721_ (.A(net2332),
    .B(net1993),
    .X(_0056_));
 sky130_fd_sc_hd__clkbuf_1 _0722_ (.A(_0056_),
    .X(\la_data_in_enable[57] ));
 sky130_fd_sc_hd__and2_1 _0723_ (.A(\mprj_logic1[388] ),
    .B(net213),
    .X(_0057_));
 sky130_fd_sc_hd__clkbuf_1 _0724_ (.A(_0057_),
    .X(\la_data_in_enable[58] ));
 sky130_fd_sc_hd__and2_1 _0725_ (.A(\mprj_logic1[389] ),
    .B(net214),
    .X(_0058_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0726_ (.A(_0058_),
    .X(\la_data_in_enable[59] ));
 sky130_fd_sc_hd__and2_1 _0727_ (.A(net2331),
    .B(net1992),
    .X(_0059_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0728_ (.A(_0059_),
    .X(\la_data_in_enable[60] ));
 sky130_fd_sc_hd__and2_1 _0729_ (.A(net2330),
    .B(net1991),
    .X(_0060_));
 sky130_fd_sc_hd__clkbuf_1 _0730_ (.A(_0060_),
    .X(\la_data_in_enable[61] ));
 sky130_fd_sc_hd__and2_1 _0731_ (.A(\mprj_logic1[392] ),
    .B(net218),
    .X(_0061_));
 sky130_fd_sc_hd__clkbuf_1 _0732_ (.A(_0061_),
    .X(\la_data_in_enable[62] ));
 sky130_fd_sc_hd__and2_1 _0733_ (.A(\mprj_logic1[393] ),
    .B(net219),
    .X(_0062_));
 sky130_fd_sc_hd__clkbuf_1 _0734_ (.A(_0062_),
    .X(\la_data_in_enable[63] ));
 sky130_fd_sc_hd__and2_1 _0735_ (.A(\mprj_logic1[394] ),
    .B(net220),
    .X(_0063_));
 sky130_fd_sc_hd__clkbuf_1 _0736_ (.A(_0063_),
    .X(\la_data_in_enable[64] ));
 sky130_fd_sc_hd__and2_1 _0737_ (.A(\mprj_logic1[395] ),
    .B(net221),
    .X(_0064_));
 sky130_fd_sc_hd__clkbuf_1 _0738_ (.A(_0064_),
    .X(\la_data_in_enable[65] ));
 sky130_fd_sc_hd__and2_1 _0739_ (.A(\mprj_logic1[396] ),
    .B(net222),
    .X(_0065_));
 sky130_fd_sc_hd__clkbuf_1 _0740_ (.A(_0065_),
    .X(\la_data_in_enable[66] ));
 sky130_fd_sc_hd__and2_1 _0741_ (.A(\mprj_logic1[397] ),
    .B(net223),
    .X(_0066_));
 sky130_fd_sc_hd__clkbuf_1 _0742_ (.A(_0066_),
    .X(\la_data_in_enable[67] ));
 sky130_fd_sc_hd__and2_1 _0743_ (.A(\mprj_logic1[398] ),
    .B(net224),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_1 _0744_ (.A(_0067_),
    .X(\la_data_in_enable[68] ));
 sky130_fd_sc_hd__and2_1 _0745_ (.A(\mprj_logic1[399] ),
    .B(net1990),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_1 _0746_ (.A(_0068_),
    .X(\la_data_in_enable[69] ));
 sky130_fd_sc_hd__and2_1 _0747_ (.A(net2329),
    .B(net1989),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_1 _0748_ (.A(_0069_),
    .X(\la_data_in_enable[70] ));
 sky130_fd_sc_hd__and2_1 _0749_ (.A(net2328),
    .B(net1988),
    .X(_0070_));
 sky130_fd_sc_hd__clkbuf_1 _0750_ (.A(_0070_),
    .X(\la_data_in_enable[71] ));
 sky130_fd_sc_hd__and2_1 _0751_ (.A(net2327),
    .B(net1987),
    .X(_0071_));
 sky130_fd_sc_hd__clkbuf_1 _0752_ (.A(net1630),
    .X(\la_data_in_enable[72] ));
 sky130_fd_sc_hd__and2_1 _0753_ (.A(net2325),
    .B(net1985),
    .X(_0072_));
 sky130_fd_sc_hd__clkbuf_1 _0754_ (.A(_0072_),
    .X(\la_data_in_enable[73] ));
 sky130_fd_sc_hd__and2_1 _0755_ (.A(net2323),
    .B(net1983),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_1 _0756_ (.A(_0073_),
    .X(\la_data_in_enable[74] ));
 sky130_fd_sc_hd__and2_1 _0757_ (.A(net2321),
    .B(net1981),
    .X(_0074_));
 sky130_fd_sc_hd__clkbuf_1 _0758_ (.A(net1629),
    .X(\la_data_in_enable[75] ));
 sky130_fd_sc_hd__and2_4 _0759_ (.A(net2320),
    .B(net1980),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_1 _0760_ (.A(net1627),
    .X(\la_data_in_enable[76] ));
 sky130_fd_sc_hd__and2_4 _0761_ (.A(net2319),
    .B(net1979),
    .X(_0076_));
 sky130_fd_sc_hd__clkbuf_1 _0762_ (.A(net1625),
    .X(\la_data_in_enable[77] ));
 sky130_fd_sc_hd__and2_1 _0763_ (.A(net2318),
    .B(net235),
    .X(_0077_));
 sky130_fd_sc_hd__clkbuf_1 _0764_ (.A(net1623),
    .X(\la_data_in_enable[78] ));
 sky130_fd_sc_hd__and2_1 _0765_ (.A(net2317),
    .B(net236),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_1 _0766_ (.A(net1621),
    .X(\la_data_in_enable[79] ));
 sky130_fd_sc_hd__and2_1 _0767_ (.A(net2314),
    .B(net1977),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0768_ (.A(net1620),
    .X(\la_data_in_enable[80] ));
 sky130_fd_sc_hd__and2_1 _0769_ (.A(\mprj_logic1[411] ),
    .B(net239),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0770_ (.A(net1617),
    .X(\la_data_in_enable[81] ));
 sky130_fd_sc_hd__and2_2 _0771_ (.A(\mprj_logic1[412] ),
    .B(net240),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_1 _0772_ (.A(net1615),
    .X(\la_data_in_enable[82] ));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(net2313),
    .B(net241),
    .X(_0082_));
 sky130_fd_sc_hd__clkbuf_1 _0774_ (.A(net1612),
    .X(\la_data_in_enable[83] ));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(net2312),
    .B(net242),
    .X(_0083_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0776_ (.A(net1609),
    .X(\la_data_in_enable[84] ));
 sky130_fd_sc_hd__and2_1 _0777_ (.A(net2311),
    .B(net243),
    .X(_0084_));
 sky130_fd_sc_hd__clkbuf_1 _0778_ (.A(net1607),
    .X(\la_data_in_enable[85] ));
 sky130_fd_sc_hd__and2_1 _0779_ (.A(net2310),
    .B(net244),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0780_ (.A(net1605),
    .X(\la_data_in_enable[86] ));
 sky130_fd_sc_hd__and2_1 _0781_ (.A(net2307),
    .B(net1975),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0782_ (.A(_0086_),
    .X(\la_data_in_enable[87] ));
 sky130_fd_sc_hd__and2_1 _0783_ (.A(net2306),
    .B(net246),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_1 _0784_ (.A(net1602),
    .X(\la_data_in_enable[88] ));
 sky130_fd_sc_hd__and2_1 _0785_ (.A(net2305),
    .B(net247),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_1 _0786_ (.A(net1600),
    .X(\la_data_in_enable[89] ));
 sky130_fd_sc_hd__and2_1 _0787_ (.A(\mprj_logic1[420] ),
    .B(net249),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_1 _0788_ (.A(net1597),
    .X(\la_data_in_enable[90] ));
 sky130_fd_sc_hd__and2_1 _0789_ (.A(net2304),
    .B(net250),
    .X(_0090_));
 sky130_fd_sc_hd__clkbuf_1 _0790_ (.A(net1594),
    .X(\la_data_in_enable[91] ));
 sky130_fd_sc_hd__and2_1 _0791_ (.A(net2303),
    .B(net251),
    .X(_0091_));
 sky130_fd_sc_hd__clkbuf_1 _0792_ (.A(net1591),
    .X(\la_data_in_enable[92] ));
 sky130_fd_sc_hd__and2_1 _0793_ (.A(net2302),
    .B(net252),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_2 _0794_ (.A(net1588),
    .X(\la_data_in_enable[93] ));
 sky130_fd_sc_hd__and2_1 _0795_ (.A(net2301),
    .B(net253),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_1 _0796_ (.A(net1585),
    .X(\la_data_in_enable[94] ));
 sky130_fd_sc_hd__and2_1 _0797_ (.A(net2300),
    .B(net254),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_1 _0798_ (.A(net1582),
    .X(\la_data_in_enable[95] ));
 sky130_fd_sc_hd__and2_1 _0799_ (.A(net2299),
    .B(net255),
    .X(_0095_));
 sky130_fd_sc_hd__clkbuf_1 _0800_ (.A(net1580),
    .X(\la_data_in_enable[96] ));
 sky130_fd_sc_hd__and2_1 _0801_ (.A(net2298),
    .B(net256),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_1 _0802_ (.A(net1577),
    .X(\la_data_in_enable[97] ));
 sky130_fd_sc_hd__and2_1 _0803_ (.A(net2297),
    .B(net257),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_1 _0804_ (.A(net1575),
    .X(\la_data_in_enable[98] ));
 sky130_fd_sc_hd__and2_1 _0805_ (.A(net2296),
    .B(net258),
    .X(_0098_));
 sky130_fd_sc_hd__clkbuf_1 _0806_ (.A(net1572),
    .X(\la_data_in_enable[99] ));
 sky130_fd_sc_hd__and2_1 _0807_ (.A(net2295),
    .B(net133),
    .X(_0099_));
 sky130_fd_sc_hd__clkbuf_1 _0808_ (.A(net1570),
    .X(\la_data_in_enable[100] ));
 sky130_fd_sc_hd__and2_4 _0809_ (.A(\mprj_logic1[431] ),
    .B(net134),
    .X(_0100_));
 sky130_fd_sc_hd__clkbuf_1 _0810_ (.A(net1567),
    .X(\la_data_in_enable[101] ));
 sky130_fd_sc_hd__and2_1 _0811_ (.A(net2294),
    .B(net135),
    .X(_0101_));
 sky130_fd_sc_hd__clkbuf_1 _0812_ (.A(net1564),
    .X(\la_data_in_enable[102] ));
 sky130_fd_sc_hd__and2_1 _0813_ (.A(\mprj_logic1[433] ),
    .B(net136),
    .X(_0102_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0814_ (.A(net1561),
    .X(\la_data_in_enable[103] ));
 sky130_fd_sc_hd__and2_1 _0815_ (.A(net2293),
    .B(net137),
    .X(_0103_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0816_ (.A(net1558),
    .X(\la_data_in_enable[104] ));
 sky130_fd_sc_hd__and2_1 _0817_ (.A(net2292),
    .B(net138),
    .X(_0104_));
 sky130_fd_sc_hd__clkbuf_1 _0818_ (.A(net1556),
    .X(\la_data_in_enable[105] ));
 sky130_fd_sc_hd__and2_1 _0819_ (.A(net2290),
    .B(net139),
    .X(_0105_));
 sky130_fd_sc_hd__clkbuf_1 _0820_ (.A(net1555),
    .X(\la_data_in_enable[106] ));
 sky130_fd_sc_hd__and2_1 _0821_ (.A(net2287),
    .B(net2027),
    .X(_0106_));
 sky130_fd_sc_hd__clkbuf_1 _0822_ (.A(_0106_),
    .X(\la_data_in_enable[107] ));
 sky130_fd_sc_hd__and2_1 _0823_ (.A(net2284),
    .B(net2026),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _0824_ (.A(net1554),
    .X(\la_data_in_enable[108] ));
 sky130_fd_sc_hd__and2_1 _0825_ (.A(net2281),
    .B(net2025),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_1 _0826_ (.A(_0108_),
    .X(\la_data_in_enable[109] ));
 sky130_fd_sc_hd__and2_2 _0827_ (.A(net2279),
    .B(net2023),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0828_ (.A(_0109_),
    .X(\la_data_in_enable[110] ));
 sky130_fd_sc_hd__and2_1 _0829_ (.A(net2276),
    .B(net2022),
    .X(_0110_));
 sky130_fd_sc_hd__clkbuf_1 _0830_ (.A(_0110_),
    .X(\la_data_in_enable[111] ));
 sky130_fd_sc_hd__and2_1 _0831_ (.A(net2273),
    .B(net2020),
    .X(_0111_));
 sky130_fd_sc_hd__clkbuf_1 _0832_ (.A(_0111_),
    .X(\la_data_in_enable[112] ));
 sky130_fd_sc_hd__and2_1 _0833_ (.A(net2270),
    .B(net2019),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0834_ (.A(_0112_),
    .X(\la_data_in_enable[113] ));
 sky130_fd_sc_hd__and2_1 _0835_ (.A(net2268),
    .B(net148),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _0836_ (.A(net1553),
    .X(\la_data_in_enable[114] ));
 sky130_fd_sc_hd__and2_1 _0837_ (.A(net2264),
    .B(net2017),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_1 _0838_ (.A(_0114_),
    .X(\la_data_in_enable[115] ));
 sky130_fd_sc_hd__and2_1 _0839_ (.A(net2262),
    .B(net150),
    .X(_0115_));
 sky130_fd_sc_hd__clkbuf_1 _0840_ (.A(net1552),
    .X(\la_data_in_enable[116] ));
 sky130_fd_sc_hd__and2_1 _0841_ (.A(net2259),
    .B(net2016),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0842_ (.A(_0116_),
    .X(\la_data_in_enable[117] ));
 sky130_fd_sc_hd__and2_1 _0843_ (.A(net2256),
    .B(net2015),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_1 _0844_ (.A(_0117_),
    .X(\la_data_in_enable[118] ));
 sky130_fd_sc_hd__and2_1 _0845_ (.A(net2254),
    .B(net153),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_1 _0846_ (.A(_0118_),
    .X(\la_data_in_enable[119] ));
 sky130_fd_sc_hd__and2_1 _0847_ (.A(net2249),
    .B(net2013),
    .X(_0119_));
 sky130_fd_sc_hd__clkbuf_1 _0848_ (.A(_0119_),
    .X(\la_data_in_enable[120] ));
 sky130_fd_sc_hd__and2_1 _0849_ (.A(net2246),
    .B(net2012),
    .X(_0120_));
 sky130_fd_sc_hd__clkbuf_1 _0850_ (.A(_0120_),
    .X(\la_data_in_enable[121] ));
 sky130_fd_sc_hd__and2_1 _0851_ (.A(net2243),
    .B(net2011),
    .X(_0121_));
 sky130_fd_sc_hd__clkbuf_1 _0852_ (.A(_0121_),
    .X(\la_data_in_enable[122] ));
 sky130_fd_sc_hd__and2_1 _0853_ (.A(net2240),
    .B(net2010),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_1 _0854_ (.A(_0122_),
    .X(\la_data_in_enable[123] ));
 sky130_fd_sc_hd__and2_1 _0855_ (.A(net2237),
    .B(net2009),
    .X(_0123_));
 sky130_fd_sc_hd__clkbuf_1 _0856_ (.A(_0123_),
    .X(\la_data_in_enable[124] ));
 sky130_fd_sc_hd__and2_1 _0857_ (.A(net2234),
    .B(net160),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0858_ (.A(_0124_),
    .X(\la_data_in_enable[125] ));
 sky130_fd_sc_hd__and2_1 _0859_ (.A(net2231),
    .B(net2008),
    .X(_0125_));
 sky130_fd_sc_hd__clkbuf_1 _0860_ (.A(_0125_),
    .X(\la_data_in_enable[126] ));
 sky130_fd_sc_hd__and2_2 _0861_ (.A(net2229),
    .B(net162),
    .X(_0126_));
 sky130_fd_sc_hd__clkbuf_1 _0862_ (.A(_0126_),
    .X(\la_data_in_enable[127] ));
 sky130_fd_sc_hd__and2_1 _0863_ (.A(net2225),
    .B(net460),
    .X(_0127_));
 sky130_fd_sc_hd__clkbuf_1 _0864_ (.A(_0127_),
    .X(\user_irq_enable[0] ));
 sky130_fd_sc_hd__and2_1 _0865_ (.A(net2221),
    .B(net461),
    .X(_0128_));
 sky130_fd_sc_hd__clkbuf_1 _0866_ (.A(_0128_),
    .X(\user_irq_enable[1] ));
 sky130_fd_sc_hd__and2_1 _0867_ (.A(net2218),
    .B(net462),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_1 _0868_ (.A(_0129_),
    .X(\user_irq_enable[2] ));
 sky130_fd_sc_hd__and2_1 _0869_ (.A(net2210),
    .B(net453),
    .X(_0130_));
 sky130_fd_sc_hd__buf_6 _0870_ (.A(_0130_),
    .X(wb_in_enable));
 sky130_fd_sc_hd__and2b_1 _0871_ (.A_N(net1930),
    .B(net2848),
    .X(_0131_));
 sky130_fd_sc_hd__buf_2 _0872_ (.A(_0131_),
    .X(net960));
 sky130_fd_sc_hd__and2_2 _0873_ (.A(\mprj_logic1[1] ),
    .B(net2066),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0874_ (.A(_0132_),
    .X(net955));
 sky130_fd_sc_hd__and2_1 _0875_ (.A(net2524),
    .B(net2),
    .X(_0133_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0876_ (.A(_0133_),
    .X(net956));
 sky130_fd_sc_hd__and2_1 _0877_ (.A(\mprj_logic1[3] ),
    .B(net1697),
    .X(_0134_));
 sky130_fd_sc_hd__buf_6 _0878_ (.A(_0134_),
    .X(net880));
 sky130_fd_sc_hd__and2_1 _0879_ (.A(net2208),
    .B(net1650),
    .X(_0135_));
 sky130_fd_sc_hd__buf_6 _0880_ (.A(net1551),
    .X(net949));
 sky130_fd_sc_hd__and2_1 _0881_ (.A(net2195),
    .B(net1649),
    .X(_0136_));
 sky130_fd_sc_hd__buf_6 _0882_ (.A(net1550),
    .X(net950));
 sky130_fd_sc_hd__and2_1 _0883_ (.A(net2174),
    .B(net454),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0884_ (.A(net1549),
    .X(net945));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(net2148),
    .B(net455),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0886_ (.A(net1548),
    .X(net946));
 sky130_fd_sc_hd__and2_1 _0887_ (.A(net2109),
    .B(net456),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0888_ (.A(net1546),
    .X(net947));
 sky130_fd_sc_hd__and2_1 _0889_ (.A(net2075),
    .B(net457),
    .X(_0140_));
 sky130_fd_sc_hd__buf_6 _0890_ (.A(net1543),
    .X(net948));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(net2837),
    .B(net1826),
    .X(_0141_));
 sky130_fd_sc_hd__clkbuf_1 _0892_ (.A(_0141_),
    .X(net848));
 sky130_fd_sc_hd__and2_2 _0893_ (.A(\mprj_logic1[11] ),
    .B(net1786),
    .X(_0142_));
 sky130_fd_sc_hd__clkbuf_2 _0894_ (.A(_0142_),
    .X(net859));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(net2829),
    .B(net1738),
    .X(_0143_));
 sky130_fd_sc_hd__buf_2 _0896_ (.A(_0143_),
    .X(net870));
 sky130_fd_sc_hd__and2_1 _0897_ (.A(\mprj_logic1[13] ),
    .B(net1726),
    .X(_0144_));
 sky130_fd_sc_hd__clkbuf_2 _0898_ (.A(_0144_),
    .X(net873));
 sky130_fd_sc_hd__and2_2 _0899_ (.A(net2810),
    .B(net1721),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_2 _0900_ (.A(_0145_),
    .X(net874));
 sky130_fd_sc_hd__and2_1 _0901_ (.A(\mprj_logic1[15] ),
    .B(net1717),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0902_ (.A(_0146_),
    .X(net875));
 sky130_fd_sc_hd__and2_1 _0903_ (.A(\mprj_logic1[16] ),
    .B(net1714),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0904_ (.A(_0147_),
    .X(net876));
 sky130_fd_sc_hd__and2_1 _0905_ (.A(net2742),
    .B(net1708),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_2 _0906_ (.A(net1542),
    .X(net877));
 sky130_fd_sc_hd__and2_1 _0907_ (.A(\mprj_logic1[18] ),
    .B(net1703),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_2 _0908_ (.A(net1541),
    .X(net878));
 sky130_fd_sc_hd__and2_1 _0909_ (.A(\mprj_logic1[19] ),
    .B(net1700),
    .X(_0150_));
 sky130_fd_sc_hd__buf_6 _0910_ (.A(_0150_),
    .X(net879));
 sky130_fd_sc_hd__and2_1 _0911_ (.A(\mprj_logic1[20] ),
    .B(net1824),
    .X(_0151_));
 sky130_fd_sc_hd__clkbuf_1 _0912_ (.A(_0151_),
    .X(net849));
 sky130_fd_sc_hd__and2_2 _0913_ (.A(net2635),
    .B(net1822),
    .X(_0152_));
 sky130_fd_sc_hd__buf_6 _0914_ (.A(_0152_),
    .X(net850));
 sky130_fd_sc_hd__and2_1 _0915_ (.A(\mprj_logic1[22] ),
    .B(net1818),
    .X(_0153_));
 sky130_fd_sc_hd__clkbuf_2 _0916_ (.A(_0153_),
    .X(net851));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(\mprj_logic1[23] ),
    .B(net1815),
    .X(_0154_));
 sky130_fd_sc_hd__clkbuf_2 _0918_ (.A(_0154_),
    .X(net852));
 sky130_fd_sc_hd__and2_1 _0919_ (.A(\mprj_logic1[24] ),
    .B(net1812),
    .X(_0155_));
 sky130_fd_sc_hd__clkbuf_1 _0920_ (.A(_0155_),
    .X(net853));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(\mprj_logic1[25] ),
    .B(net1807),
    .X(_0156_));
 sky130_fd_sc_hd__clkbuf_1 _0922_ (.A(_0156_),
    .X(net854));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(net2597),
    .B(net1802),
    .X(_0157_));
 sky130_fd_sc_hd__buf_2 _0924_ (.A(_0157_),
    .X(net855));
 sky130_fd_sc_hd__and2_1 _0925_ (.A(\mprj_logic1[27] ),
    .B(net1799),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0926_ (.A(_0158_),
    .X(net856));
 sky130_fd_sc_hd__and2_1 _0927_ (.A(net2547),
    .B(net1794),
    .X(_0159_));
 sky130_fd_sc_hd__clkbuf_2 _0928_ (.A(_0159_),
    .X(net857));
 sky130_fd_sc_hd__and2_1 _0929_ (.A(\mprj_logic1[29] ),
    .B(net1790),
    .X(_0160_));
 sky130_fd_sc_hd__clkbuf_2 _0930_ (.A(_0160_),
    .X(net858));
 sky130_fd_sc_hd__and2_1 _0931_ (.A(\mprj_logic1[30] ),
    .B(net1783),
    .X(_0161_));
 sky130_fd_sc_hd__clkbuf_2 _0932_ (.A(_0161_),
    .X(net860));
 sky130_fd_sc_hd__and2_1 _0933_ (.A(net2462),
    .B(net1778),
    .X(_0162_));
 sky130_fd_sc_hd__clkbuf_2 _0934_ (.A(_0162_),
    .X(net861));
 sky130_fd_sc_hd__and2_1 _0935_ (.A(\mprj_logic1[32] ),
    .B(net1775),
    .X(_0163_));
 sky130_fd_sc_hd__buf_6 _0936_ (.A(_0163_),
    .X(net862));
 sky130_fd_sc_hd__and2_1 _0937_ (.A(\mprj_logic1[33] ),
    .B(net1771),
    .X(_0164_));
 sky130_fd_sc_hd__clkbuf_1 _0938_ (.A(_0164_),
    .X(net863));
 sky130_fd_sc_hd__and2_2 _0939_ (.A(\mprj_logic1[34] ),
    .B(net1766),
    .X(_0165_));
 sky130_fd_sc_hd__clkbuf_2 _0940_ (.A(_0165_),
    .X(net864));
 sky130_fd_sc_hd__and2_1 _0941_ (.A(\mprj_logic1[35] ),
    .B(net1761),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_2 _0942_ (.A(_0166_),
    .X(net865));
 sky130_fd_sc_hd__and2_1 _0943_ (.A(\mprj_logic1[36] ),
    .B(net1757),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_2 _0944_ (.A(_0167_),
    .X(net866));
 sky130_fd_sc_hd__and2_1 _0945_ (.A(\mprj_logic1[37] ),
    .B(net1752),
    .X(_0168_));
 sky130_fd_sc_hd__clkbuf_2 _0946_ (.A(_0168_),
    .X(net867));
 sky130_fd_sc_hd__and2_1 _0947_ (.A(\mprj_logic1[38] ),
    .B(net1748),
    .X(_0169_));
 sky130_fd_sc_hd__buf_4 _0948_ (.A(_0169_),
    .X(net868));
 sky130_fd_sc_hd__and2_1 _0949_ (.A(\mprj_logic1[39] ),
    .B(net1744),
    .X(_0170_));
 sky130_fd_sc_hd__clkbuf_2 _0950_ (.A(_0170_),
    .X(net869));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(\mprj_logic1[40] ),
    .B(net1734),
    .X(_0171_));
 sky130_fd_sc_hd__clkbuf_1 _0952_ (.A(_0171_),
    .X(net871));
 sky130_fd_sc_hd__and2_1 _0953_ (.A(\mprj_logic1[41] ),
    .B(net1730),
    .X(_0172_));
 sky130_fd_sc_hd__clkbuf_1 _0954_ (.A(_0172_),
    .X(net872));
 sky130_fd_sc_hd__and2_1 _0955_ (.A(\mprj_logic1[42] ),
    .B(net1694),
    .X(_0173_));
 sky130_fd_sc_hd__buf_6 _0956_ (.A(_0173_),
    .X(net913));
 sky130_fd_sc_hd__and2_1 _0957_ (.A(\mprj_logic1[43] ),
    .B(net1679),
    .X(_0174_));
 sky130_fd_sc_hd__buf_6 _0958_ (.A(_0174_),
    .X(net924));
 sky130_fd_sc_hd__and2_2 _0959_ (.A(net2253),
    .B(net1669),
    .X(_0175_));
 sky130_fd_sc_hd__buf_6 _0960_ (.A(net1540),
    .X(net935));
 sky130_fd_sc_hd__and2_1 _0961_ (.A(\mprj_logic1[45] ),
    .B(net1662),
    .X(_0176_));
 sky130_fd_sc_hd__buf_6 _0962_ (.A(_0176_),
    .X(net938));
 sky130_fd_sc_hd__and2_1 _0963_ (.A(\mprj_logic1[46] ),
    .B(net1660),
    .X(_0177_));
 sky130_fd_sc_hd__buf_6 _0964_ (.A(_0177_),
    .X(net939));
 sky130_fd_sc_hd__and2_1 _0965_ (.A(\mprj_logic1[47] ),
    .B(net1658),
    .X(_0178_));
 sky130_fd_sc_hd__clkbuf_1 _0966_ (.A(_0178_),
    .X(net940));
 sky130_fd_sc_hd__and2_1 _0967_ (.A(\mprj_logic1[48] ),
    .B(net1656),
    .X(_0179_));
 sky130_fd_sc_hd__clkbuf_1 _0968_ (.A(_0179_),
    .X(net941));
 sky130_fd_sc_hd__and2_1 _0969_ (.A(net2209),
    .B(net1654),
    .X(_0180_));
 sky130_fd_sc_hd__buf_6 _0970_ (.A(net1539),
    .X(net942));
 sky130_fd_sc_hd__and2_1 _0971_ (.A(\mprj_logic1[50] ),
    .B(net1652),
    .X(_0181_));
 sky130_fd_sc_hd__clkbuf_1 _0972_ (.A(_0181_),
    .X(net943));
 sky130_fd_sc_hd__and2_1 _0973_ (.A(net2207),
    .B(net1651),
    .X(_0182_));
 sky130_fd_sc_hd__buf_6 _0974_ (.A(net1538),
    .X(net944));
 sky130_fd_sc_hd__and2_1 _0975_ (.A(net2206),
    .B(net1693),
    .X(_0183_));
 sky130_fd_sc_hd__buf_6 _0976_ (.A(net1537),
    .X(net914));
 sky130_fd_sc_hd__and2_2 _0977_ (.A(net2204),
    .B(net1692),
    .X(_0184_));
 sky130_fd_sc_hd__buf_6 _0978_ (.A(net1536),
    .X(net915));
 sky130_fd_sc_hd__and2_1 _0979_ (.A(net2202),
    .B(net1691),
    .X(_0185_));
 sky130_fd_sc_hd__clkbuf_1 _0980_ (.A(net1535),
    .X(net916));
 sky130_fd_sc_hd__and2_1 _0981_ (.A(net2200),
    .B(net425),
    .X(_0186_));
 sky130_fd_sc_hd__clkbuf_1 _0982_ (.A(net1533),
    .X(net917));
 sky130_fd_sc_hd__and2_1 _0983_ (.A(net2199),
    .B(net1689),
    .X(_0187_));
 sky130_fd_sc_hd__buf_6 _0984_ (.A(net1532),
    .X(net918));
 sky130_fd_sc_hd__and2_1 _0985_ (.A(\mprj_logic1[57] ),
    .B(net1687),
    .X(_0188_));
 sky130_fd_sc_hd__buf_6 _0986_ (.A(net1531),
    .X(net919));
 sky130_fd_sc_hd__and2_2 _0987_ (.A(net2198),
    .B(net1685),
    .X(_0189_));
 sky130_fd_sc_hd__buf_6 _0988_ (.A(_0189_),
    .X(net920));
 sky130_fd_sc_hd__and2_1 _0989_ (.A(net2196),
    .B(net1684),
    .X(_0190_));
 sky130_fd_sc_hd__buf_6 _0990_ (.A(net1530),
    .X(net921));
 sky130_fd_sc_hd__and2_1 _0991_ (.A(net2194),
    .B(net1683),
    .X(_0191_));
 sky130_fd_sc_hd__buf_4 _0992_ (.A(net1528),
    .X(net922));
 sky130_fd_sc_hd__and2_1 _0993_ (.A(net2193),
    .B(net1682),
    .X(_0192_));
 sky130_fd_sc_hd__clkbuf_1 _0994_ (.A(net1526),
    .X(net923));
 sky130_fd_sc_hd__and2_2 _0995_ (.A(net2191),
    .B(net1678),
    .X(_0193_));
 sky130_fd_sc_hd__buf_6 _0996_ (.A(net1525),
    .X(net925));
 sky130_fd_sc_hd__and2_1 _0997_ (.A(net2190),
    .B(net1676),
    .X(_0194_));
 sky130_fd_sc_hd__clkbuf_1 _0998_ (.A(net1524),
    .X(net926));
 sky130_fd_sc_hd__and2_1 _0999_ (.A(net2189),
    .B(net1674),
    .X(_0195_));
 sky130_fd_sc_hd__clkbuf_1 _1000_ (.A(net1523),
    .X(net927));
 sky130_fd_sc_hd__and2_1 _1001_ (.A(net2188),
    .B(net1673),
    .X(_0196_));
 sky130_fd_sc_hd__buf_6 _1002_ (.A(net1522),
    .X(net928));
 sky130_fd_sc_hd__and2_1 _1003_ (.A(net2185),
    .B(net437),
    .X(_0197_));
 sky130_fd_sc_hd__buf_6 _1004_ (.A(net1520),
    .X(net929));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(net2182),
    .B(net438),
    .X(_0198_));
 sky130_fd_sc_hd__buf_6 _1006_ (.A(net1518),
    .X(net930));
 sky130_fd_sc_hd__and2_1 _1007_ (.A(net2180),
    .B(net439),
    .X(_0199_));
 sky130_fd_sc_hd__buf_6 _1008_ (.A(net1516),
    .X(net931));
 sky130_fd_sc_hd__and2_1 _1009_ (.A(net2176),
    .B(net440),
    .X(_0200_));
 sky130_fd_sc_hd__buf_6 _1010_ (.A(net1513),
    .X(net932));
 sky130_fd_sc_hd__and2_1 _1011_ (.A(net2172),
    .B(net1671),
    .X(_0201_));
 sky130_fd_sc_hd__buf_6 _1012_ (.A(net1512),
    .X(net933));
 sky130_fd_sc_hd__and2_1 _1013_ (.A(net2170),
    .B(net1670),
    .X(_0202_));
 sky130_fd_sc_hd__buf_6 _1014_ (.A(net1511),
    .X(net934));
 sky130_fd_sc_hd__and2_1 _1015_ (.A(net2169),
    .B(net1667),
    .X(_0203_));
 sky130_fd_sc_hd__buf_2 _1016_ (.A(net1510),
    .X(net936));
 sky130_fd_sc_hd__and2_1 _1017_ (.A(net2168),
    .B(net1665),
    .X(_0204_));
 sky130_fd_sc_hd__buf_4 _1018_ (.A(net1509),
    .X(net937));
 sky130_fd_sc_hd__and3b_1 _1019_ (.A_N(net260),
    .B(net2165),
    .C(net4),
    .X(_0205_));
 sky130_fd_sc_hd__clkbuf_2 _1020_ (.A(_0205_),
    .X(net463));
 sky130_fd_sc_hd__and3b_2 _1021_ (.A_N(net299),
    .B(net2162),
    .C(net43),
    .X(_0206_));
 sky130_fd_sc_hd__clkbuf_1 _1022_ (.A(_0206_),
    .X(net502));
 sky130_fd_sc_hd__and3b_1 _1023_ (.A_N(net310),
    .B(net2159),
    .C(net54),
    .X(_0207_));
 sky130_fd_sc_hd__clkbuf_1 _1024_ (.A(_0207_),
    .X(net513));
 sky130_fd_sc_hd__and3b_1 _1025_ (.A_N(net321),
    .B(net2156),
    .C(net65),
    .X(_0208_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1026_ (.A(_0208_),
    .X(net524));
 sky130_fd_sc_hd__and3b_1 _1027_ (.A_N(net332),
    .B(net2153),
    .C(net76),
    .X(_0209_));
 sky130_fd_sc_hd__clkbuf_2 _1028_ (.A(_0209_),
    .X(net535));
 sky130_fd_sc_hd__and3b_1 _1029_ (.A_N(net343),
    .B(net2150),
    .C(net87),
    .X(_0210_));
 sky130_fd_sc_hd__clkbuf_2 _1030_ (.A(_0210_),
    .X(net546));
 sky130_fd_sc_hd__and3b_1 _1031_ (.A_N(net354),
    .B(net2144),
    .C(net98),
    .X(_0211_));
 sky130_fd_sc_hd__clkbuf_2 _1032_ (.A(_0211_),
    .X(net557));
 sky130_fd_sc_hd__and3b_1 _1033_ (.A_N(net365),
    .B(net2140),
    .C(net109),
    .X(_0212_));
 sky130_fd_sc_hd__clkbuf_1 _1034_ (.A(net1508),
    .X(net568));
 sky130_fd_sc_hd__and3b_1 _1035_ (.A_N(net376),
    .B(net2137),
    .C(net120),
    .X(_0213_));
 sky130_fd_sc_hd__buf_2 _1036_ (.A(net1507),
    .X(net579));
 sky130_fd_sc_hd__and3b_1 _1037_ (.A_N(net387),
    .B(net2133),
    .C(net131),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_1 _1038_ (.A(net1506),
    .X(net590));
 sky130_fd_sc_hd__and3b_1 _1039_ (.A_N(net271),
    .B(net2129),
    .C(net15),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_2 _1040_ (.A(net1505),
    .X(net474));
 sky130_fd_sc_hd__and3b_1 _1041_ (.A_N(net282),
    .B(net2125),
    .C(net26),
    .X(_0216_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1042_ (.A(net1503),
    .X(net485));
 sky130_fd_sc_hd__and3b_1 _1043_ (.A_N(net291),
    .B(net2122),
    .C(net35),
    .X(_0217_));
 sky130_fd_sc_hd__clkbuf_2 _1044_ (.A(_0217_),
    .X(net494));
 sky130_fd_sc_hd__and3b_1 _1045_ (.A_N(net292),
    .B(net2119),
    .C(net36),
    .X(_0218_));
 sky130_fd_sc_hd__clkbuf_1 _1046_ (.A(net1502),
    .X(net495));
 sky130_fd_sc_hd__and3b_2 _1047_ (.A_N(net293),
    .B(net2115),
    .C(net37),
    .X(_0219_));
 sky130_fd_sc_hd__clkbuf_2 _1048_ (.A(net1501),
    .X(net496));
 sky130_fd_sc_hd__and3b_1 _1049_ (.A_N(net294),
    .B(net2111),
    .C(net38),
    .X(_0220_));
 sky130_fd_sc_hd__clkbuf_1 _1050_ (.A(net1499),
    .X(net497));
 sky130_fd_sc_hd__and3b_1 _1051_ (.A_N(net295),
    .B(net2106),
    .C(net39),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_1 _1052_ (.A(_0221_),
    .X(net498));
 sky130_fd_sc_hd__and3b_2 _1053_ (.A_N(net296),
    .B(net2103),
    .C(net40),
    .X(_0222_));
 sky130_fd_sc_hd__clkbuf_1 _1054_ (.A(net1498),
    .X(net499));
 sky130_fd_sc_hd__and3b_1 _1055_ (.A_N(net1937),
    .B(net2099),
    .C(net1743),
    .X(_0223_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1056_ (.A(net1496),
    .X(net500));
 sky130_fd_sc_hd__and3b_1 _1057_ (.A_N(net298),
    .B(net2096),
    .C(net42),
    .X(_0224_));
 sky130_fd_sc_hd__clkbuf_1 _1058_ (.A(_0224_),
    .X(net501));
 sky130_fd_sc_hd__and3b_1 _1059_ (.A_N(net1929),
    .B(net2092),
    .C(net1672),
    .X(_0225_));
 sky130_fd_sc_hd__clkbuf_1 _1060_ (.A(net1495),
    .X(net503));
 sky130_fd_sc_hd__and3b_1 _1061_ (.A_N(net301),
    .B(net2089),
    .C(net45),
    .X(_0226_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1062_ (.A(net1493),
    .X(net504));
 sky130_fd_sc_hd__and3b_1 _1063_ (.A_N(net302),
    .B(net2086),
    .C(net46),
    .X(_0227_));
 sky130_fd_sc_hd__clkbuf_2 _1064_ (.A(net1492),
    .X(net505));
 sky130_fd_sc_hd__and3b_1 _1065_ (.A_N(net303),
    .B(net2084),
    .C(net47),
    .X(_0228_));
 sky130_fd_sc_hd__clkbuf_2 _1066_ (.A(net1491),
    .X(net506));
 sky130_fd_sc_hd__and3b_1 _1067_ (.A_N(net304),
    .B(net2081),
    .C(net48),
    .X(_0229_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1068_ (.A(net1490),
    .X(net507));
 sky130_fd_sc_hd__and3b_1 _1069_ (.A_N(net305),
    .B(net2078),
    .C(net49),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_2 _1070_ (.A(net1489),
    .X(net508));
 sky130_fd_sc_hd__and3b_1 _1071_ (.A_N(net1928),
    .B(net2847),
    .C(net50),
    .X(_0231_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1072_ (.A(_0231_),
    .X(net509));
 sky130_fd_sc_hd__and3b_1 _1073_ (.A_N(net1926),
    .B(net2845),
    .C(net1648),
    .X(_0232_));
 sky130_fd_sc_hd__clkbuf_1 _1074_ (.A(_0232_),
    .X(net510));
 sky130_fd_sc_hd__and3b_1 _1075_ (.A_N(net308),
    .B(net2844),
    .C(net52),
    .X(_0233_));
 sky130_fd_sc_hd__clkbuf_2 _1076_ (.A(_0233_),
    .X(net511));
 sky130_fd_sc_hd__and3b_2 _1077_ (.A_N(net1924),
    .B(net2842),
    .C(net1647),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_1 _1078_ (.A(net1488),
    .X(net512));
 sky130_fd_sc_hd__and3b_2 _1079_ (.A_N(net311),
    .B(net2841),
    .C(net55),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_2 _1080_ (.A(_0235_),
    .X(net514));
 sky130_fd_sc_hd__and3b_1 _1081_ (.A_N(net312),
    .B(net2840),
    .C(net56),
    .X(_0236_));
 sky130_fd_sc_hd__clkbuf_1 _1082_ (.A(_0236_),
    .X(net515));
 sky130_fd_sc_hd__and3b_1 _1083_ (.A_N(net313),
    .B(net2839),
    .C(net57),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_1 _1084_ (.A(_0237_),
    .X(net516));
 sky130_fd_sc_hd__and3b_1 _1085_ (.A_N(net314),
    .B(net2838),
    .C(net58),
    .X(_0238_));
 sky130_fd_sc_hd__clkbuf_1 _1086_ (.A(_0238_),
    .X(net517));
 sky130_fd_sc_hd__and3b_1 _1087_ (.A_N(net315),
    .B(\mprj_logic1[108] ),
    .C(net59),
    .X(_0239_));
 sky130_fd_sc_hd__clkbuf_2 _1088_ (.A(_0239_),
    .X(net518));
 sky130_fd_sc_hd__and3b_1 _1089_ (.A_N(net1922),
    .B(\mprj_logic1[109] ),
    .C(net60),
    .X(_0240_));
 sky130_fd_sc_hd__clkbuf_2 _1090_ (.A(_0240_),
    .X(net519));
 sky130_fd_sc_hd__and3b_1 _1091_ (.A_N(net317),
    .B(\mprj_logic1[110] ),
    .C(net61),
    .X(_0241_));
 sky130_fd_sc_hd__clkbuf_2 _1092_ (.A(net1487),
    .X(net520));
 sky130_fd_sc_hd__and3b_1 _1093_ (.A_N(net318),
    .B(\mprj_logic1[111] ),
    .C(net62),
    .X(_0242_));
 sky130_fd_sc_hd__clkbuf_2 _1094_ (.A(_0242_),
    .X(net521));
 sky130_fd_sc_hd__and3b_1 _1095_ (.A_N(net319),
    .B(\mprj_logic1[112] ),
    .C(net63),
    .X(_0243_));
 sky130_fd_sc_hd__clkbuf_2 _1096_ (.A(net1486),
    .X(net522));
 sky130_fd_sc_hd__and3b_1 _1097_ (.A_N(net320),
    .B(\mprj_logic1[113] ),
    .C(net64),
    .X(_0244_));
 sky130_fd_sc_hd__clkbuf_2 _1098_ (.A(net1485),
    .X(net523));
 sky130_fd_sc_hd__and3b_1 _1099_ (.A_N(net1918),
    .B(net2836),
    .C(net66),
    .X(_0245_));
 sky130_fd_sc_hd__buf_4 _1100_ (.A(_0245_),
    .X(net525));
 sky130_fd_sc_hd__and3b_1 _1101_ (.A_N(net1916),
    .B(net2835),
    .C(net1646),
    .X(_0246_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1102_ (.A(net1483),
    .X(net526));
 sky130_fd_sc_hd__and3b_1 _1103_ (.A_N(net324),
    .B(\mprj_logic1[116] ),
    .C(net68),
    .X(_0247_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1104_ (.A(net1482),
    .X(net527));
 sky130_fd_sc_hd__and3b_1 _1105_ (.A_N(net1913),
    .B(net2834),
    .C(net1645),
    .X(_0248_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1106_ (.A(net1480),
    .X(net528));
 sky130_fd_sc_hd__and3b_1 _1107_ (.A_N(net326),
    .B(\mprj_logic1[118] ),
    .C(net70),
    .X(_0249_));
 sky130_fd_sc_hd__clkbuf_2 _1108_ (.A(net1479),
    .X(net529));
 sky130_fd_sc_hd__and3b_2 _1109_ (.A_N(net327),
    .B(\mprj_logic1[119] ),
    .C(net71),
    .X(_0250_));
 sky130_fd_sc_hd__clkbuf_2 _1110_ (.A(_0250_),
    .X(net530));
 sky130_fd_sc_hd__and3b_1 _1111_ (.A_N(net328),
    .B(\mprj_logic1[120] ),
    .C(net72),
    .X(_0251_));
 sky130_fd_sc_hd__clkbuf_2 _1112_ (.A(net1478),
    .X(net531));
 sky130_fd_sc_hd__and3b_2 _1113_ (.A_N(net1910),
    .B(net2833),
    .C(net73),
    .X(_0252_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1114_ (.A(net1477),
    .X(net532));
 sky130_fd_sc_hd__and3b_2 _1115_ (.A_N(net330),
    .B(\mprj_logic1[122] ),
    .C(net74),
    .X(_0253_));
 sky130_fd_sc_hd__clkbuf_1 _1116_ (.A(_0253_),
    .X(net533));
 sky130_fd_sc_hd__and3b_1 _1117_ (.A_N(net331),
    .B(\mprj_logic1[123] ),
    .C(net75),
    .X(_0254_));
 sky130_fd_sc_hd__clkbuf_2 _1118_ (.A(net1476),
    .X(net534));
 sky130_fd_sc_hd__and3b_1 _1119_ (.A_N(net333),
    .B(\mprj_logic1[124] ),
    .C(net77),
    .X(_0255_));
 sky130_fd_sc_hd__clkbuf_2 _1120_ (.A(net1475),
    .X(net536));
 sky130_fd_sc_hd__and3b_1 _1121_ (.A_N(net1902),
    .B(\mprj_logic1[125] ),
    .C(net78),
    .X(_0256_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1122_ (.A(net1473),
    .X(net537));
 sky130_fd_sc_hd__and3b_1 _1123_ (.A_N(net1900),
    .B(net2832),
    .C(net1644),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_2 _1124_ (.A(net1471),
    .X(net538));
 sky130_fd_sc_hd__and3b_1 _1125_ (.A_N(net1899),
    .B(net2831),
    .C(net1643),
    .X(_0258_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1126_ (.A(net1469),
    .X(net539));
 sky130_fd_sc_hd__and3b_1 _1127_ (.A_N(net1896),
    .B(net2830),
    .C(net1642),
    .X(_0259_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1128_ (.A(net1466),
    .X(net540));
 sky130_fd_sc_hd__and3b_1 _1129_ (.A_N(net1895),
    .B(\mprj_logic1[129] ),
    .C(net1641),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_2 _1130_ (.A(net1464),
    .X(net541));
 sky130_fd_sc_hd__and3b_1 _1131_ (.A_N(net339),
    .B(\mprj_logic1[130] ),
    .C(net83),
    .X(_0261_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1132_ (.A(net1462),
    .X(net542));
 sky130_fd_sc_hd__and3b_1 _1133_ (.A_N(net1891),
    .B(\mprj_logic1[131] ),
    .C(net84),
    .X(_0262_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1134_ (.A(net1460),
    .X(net543));
 sky130_fd_sc_hd__and3b_1 _1135_ (.A_N(net1890),
    .B(\mprj_logic1[132] ),
    .C(net1640),
    .X(_0263_));
 sky130_fd_sc_hd__clkbuf_2 _1136_ (.A(net1458),
    .X(net544));
 sky130_fd_sc_hd__and3b_1 _1137_ (.A_N(net1889),
    .B(\mprj_logic1[133] ),
    .C(net86),
    .X(_0264_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1138_ (.A(net1456),
    .X(net545));
 sky130_fd_sc_hd__and3b_1 _1139_ (.A_N(net1886),
    .B(net2828),
    .C(net1639),
    .X(_0265_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1140_ (.A(net1453),
    .X(net547));
 sky130_fd_sc_hd__and3b_1 _1141_ (.A_N(net1885),
    .B(\mprj_logic1[135] ),
    .C(net1638),
    .X(_0266_));
 sky130_fd_sc_hd__clkbuf_2 _1142_ (.A(net1451),
    .X(net548));
 sky130_fd_sc_hd__and3b_1 _1143_ (.A_N(net1884),
    .B(\mprj_logic1[136] ),
    .C(net1637),
    .X(_0267_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1144_ (.A(net1449),
    .X(net549));
 sky130_fd_sc_hd__and3b_1 _1145_ (.A_N(net1882),
    .B(\mprj_logic1[137] ),
    .C(net1636),
    .X(_0268_));
 sky130_fd_sc_hd__clkbuf_2 _1146_ (.A(net1447),
    .X(net550));
 sky130_fd_sc_hd__and3b_1 _1147_ (.A_N(net348),
    .B(\mprj_logic1[138] ),
    .C(net92),
    .X(_0269_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1148_ (.A(net1446),
    .X(net551));
 sky130_fd_sc_hd__and3b_1 _1149_ (.A_N(net349),
    .B(\mprj_logic1[139] ),
    .C(net93),
    .X(_0270_));
 sky130_fd_sc_hd__clkbuf_2 _1150_ (.A(net1445),
    .X(net552));
 sky130_fd_sc_hd__and3b_1 _1151_ (.A_N(net1878),
    .B(\mprj_logic1[140] ),
    .C(net94),
    .X(_0271_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1152_ (.A(net1444),
    .X(net553));
 sky130_fd_sc_hd__and3b_1 _1153_ (.A_N(net1876),
    .B(net2827),
    .C(net1635),
    .X(_0272_));
 sky130_fd_sc_hd__clkbuf_2 _1154_ (.A(_0272_),
    .X(net554));
 sky130_fd_sc_hd__and3b_1 _1155_ (.A_N(net1875),
    .B(net2825),
    .C(net1634),
    .X(_0273_));
 sky130_fd_sc_hd__clkbuf_2 _1156_ (.A(_0273_),
    .X(net555));
 sky130_fd_sc_hd__and3b_1 _1157_ (.A_N(net1874),
    .B(net2824),
    .C(net97),
    .X(_0274_));
 sky130_fd_sc_hd__buf_2 _1158_ (.A(_0274_),
    .X(net556));
 sky130_fd_sc_hd__and3b_1 _1159_ (.A_N(net1873),
    .B(net2822),
    .C(net1633),
    .X(_0275_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1160_ (.A(_0275_),
    .X(net558));
 sky130_fd_sc_hd__and3b_1 _1161_ (.A_N(net1872),
    .B(net2820),
    .C(net2064),
    .X(_0276_));
 sky130_fd_sc_hd__clkbuf_2 _1162_ (.A(_0276_),
    .X(net559));
 sky130_fd_sc_hd__and3b_1 _1163_ (.A_N(net1871),
    .B(net2818),
    .C(net2063),
    .X(_0277_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1164_ (.A(_0277_),
    .X(net560));
 sky130_fd_sc_hd__and3b_1 _1165_ (.A_N(net1870),
    .B(net2816),
    .C(net2062),
    .X(_0278_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1166_ (.A(_0278_),
    .X(net561));
 sky130_fd_sc_hd__and3b_1 _1167_ (.A_N(net1868),
    .B(net2813),
    .C(net2060),
    .X(_0279_));
 sky130_fd_sc_hd__clkbuf_2 _1168_ (.A(_0279_),
    .X(net562));
 sky130_fd_sc_hd__and3b_1 _1169_ (.A_N(net1867),
    .B(net2811),
    .C(net2059),
    .X(_0280_));
 sky130_fd_sc_hd__clkbuf_2 _1170_ (.A(_0280_),
    .X(net563));
 sky130_fd_sc_hd__and3b_1 _1171_ (.A_N(net1865),
    .B(net2807),
    .C(net2057),
    .X(_0281_));
 sky130_fd_sc_hd__buf_2 _1172_ (.A(_0281_),
    .X(net564));
 sky130_fd_sc_hd__and3b_1 _1173_ (.A_N(net1863),
    .B(net2804),
    .C(net2054),
    .X(_0282_));
 sky130_fd_sc_hd__clkbuf_2 _1174_ (.A(net1443),
    .X(net565));
 sky130_fd_sc_hd__and3b_1 _1175_ (.A_N(net1861),
    .B(net2801),
    .C(net2052),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_2 _1176_ (.A(_0283_),
    .X(net566));
 sky130_fd_sc_hd__and3b_2 _1177_ (.A_N(net1860),
    .B(net2799),
    .C(net2051),
    .X(_0284_));
 sky130_fd_sc_hd__clkbuf_2 _1178_ (.A(_0284_),
    .X(net567));
 sky130_fd_sc_hd__and3b_1 _1179_ (.A_N(net1857),
    .B(net2795),
    .C(net2048),
    .X(_0285_));
 sky130_fd_sc_hd__clkbuf_2 _1180_ (.A(_0285_),
    .X(net569));
 sky130_fd_sc_hd__and3b_1 _1181_ (.A_N(net1855),
    .B(net2791),
    .C(net2046),
    .X(_0286_));
 sky130_fd_sc_hd__clkbuf_1 _1182_ (.A(_0286_),
    .X(net570));
 sky130_fd_sc_hd__and3b_1 _1183_ (.A_N(net1853),
    .B(net2787),
    .C(net2043),
    .X(_0287_));
 sky130_fd_sc_hd__clkbuf_2 _1184_ (.A(_0287_),
    .X(net571));
 sky130_fd_sc_hd__and3b_1 _1185_ (.A_N(net1851),
    .B(net2783),
    .C(net2040),
    .X(_0288_));
 sky130_fd_sc_hd__clkbuf_1 _1186_ (.A(_0288_),
    .X(net572));
 sky130_fd_sc_hd__and3b_1 _1187_ (.A_N(net1849),
    .B(net2780),
    .C(net2038),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_1 _1188_ (.A(_0289_),
    .X(net573));
 sky130_fd_sc_hd__and3b_1 _1189_ (.A_N(net1847),
    .B(net2776),
    .C(net2036),
    .X(_0290_));
 sky130_fd_sc_hd__buf_2 _1190_ (.A(_0290_),
    .X(net574));
 sky130_fd_sc_hd__and3b_1 _1191_ (.A_N(net1845),
    .B(net2772),
    .C(net2033),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_1 _1192_ (.A(_0291_),
    .X(net575));
 sky130_fd_sc_hd__and3b_1 _1193_ (.A_N(net1843),
    .B(net2767),
    .C(net2030),
    .X(_0292_));
 sky130_fd_sc_hd__clkbuf_2 _1194_ (.A(_0292_),
    .X(net576));
 sky130_fd_sc_hd__and3b_1 _1195_ (.A_N(net1842),
    .B(net2764),
    .C(net2029),
    .X(_0293_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1196_ (.A(_0293_),
    .X(net577));
 sky130_fd_sc_hd__and3b_1 _1197_ (.A_N(net375),
    .B(net2763),
    .C(net119),
    .X(_0294_));
 sky130_fd_sc_hd__clkbuf_1 _1198_ (.A(_0294_),
    .X(net578));
 sky130_fd_sc_hd__and3b_1 _1199_ (.A_N(net377),
    .B(net2762),
    .C(net121),
    .X(_0295_));
 sky130_fd_sc_hd__buf_2 _1200_ (.A(net1442),
    .X(net580));
 sky130_fd_sc_hd__and3b_1 _1201_ (.A_N(net378),
    .B(net2761),
    .C(net122),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_1 _1202_ (.A(net1440),
    .X(net581));
 sky130_fd_sc_hd__and3b_1 _1203_ (.A_N(net379),
    .B(net2760),
    .C(net123),
    .X(_0297_));
 sky130_fd_sc_hd__clkbuf_1 _1204_ (.A(net1438),
    .X(net582));
 sky130_fd_sc_hd__and3b_1 _1205_ (.A_N(net380),
    .B(\mprj_logic1[167] ),
    .C(net124),
    .X(_0298_));
 sky130_fd_sc_hd__clkbuf_2 _1206_ (.A(net1435),
    .X(net583));
 sky130_fd_sc_hd__and3b_1 _1207_ (.A_N(net381),
    .B(net2759),
    .C(net125),
    .X(_0299_));
 sky130_fd_sc_hd__clkbuf_2 _1208_ (.A(net1432),
    .X(net584));
 sky130_fd_sc_hd__and3b_1 _1209_ (.A_N(net382),
    .B(net2757),
    .C(net126),
    .X(_0300_));
 sky130_fd_sc_hd__clkbuf_2 _1210_ (.A(net1430),
    .X(net585));
 sky130_fd_sc_hd__and3b_1 _1211_ (.A_N(net1837),
    .B(net2756),
    .C(net127),
    .X(_0301_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1212_ (.A(net1428),
    .X(net586));
 sky130_fd_sc_hd__and3b_1 _1213_ (.A_N(net384),
    .B(net2755),
    .C(net128),
    .X(_0302_));
 sky130_fd_sc_hd__buf_2 _1214_ (.A(net1426),
    .X(net587));
 sky130_fd_sc_hd__and3b_1 _1215_ (.A_N(net385),
    .B(net2754),
    .C(net129),
    .X(_0303_));
 sky130_fd_sc_hd__clkbuf_1 _1216_ (.A(_0303_),
    .X(net588));
 sky130_fd_sc_hd__and3b_1 _1217_ (.A_N(net1832),
    .B(net2753),
    .C(net130),
    .X(_0304_));
 sky130_fd_sc_hd__buf_4 _1218_ (.A(_0304_),
    .X(net589));
 sky130_fd_sc_hd__and3b_1 _1219_ (.A_N(net1973),
    .B(net2751),
    .C(net5),
    .X(_0305_));
 sky130_fd_sc_hd__buf_2 _1220_ (.A(net1424),
    .X(net464));
 sky130_fd_sc_hd__and3b_1 _1221_ (.A_N(net262),
    .B(net2750),
    .C(net6),
    .X(_0306_));
 sky130_fd_sc_hd__clkbuf_1 _1222_ (.A(net1422),
    .X(net465));
 sky130_fd_sc_hd__and3b_1 _1223_ (.A_N(net1970),
    .B(net2748),
    .C(net7),
    .X(_0307_));
 sky130_fd_sc_hd__clkbuf_2 _1224_ (.A(net1421),
    .X(net466));
 sky130_fd_sc_hd__and3b_1 _1225_ (.A_N(net264),
    .B(net2746),
    .C(net8),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_1 _1226_ (.A(net1419),
    .X(net467));
 sky130_fd_sc_hd__and3b_1 _1227_ (.A_N(net265),
    .B(net2745),
    .C(net9),
    .X(_0309_));
 sky130_fd_sc_hd__clkbuf_2 _1228_ (.A(_0309_),
    .X(net468));
 sky130_fd_sc_hd__and3b_2 _1229_ (.A_N(net266),
    .B(net2743),
    .C(net10),
    .X(_0310_));
 sky130_fd_sc_hd__clkbuf_1 _1230_ (.A(_0310_),
    .X(net469));
 sky130_fd_sc_hd__and3b_1 _1231_ (.A_N(net267),
    .B(net2741),
    .C(net11),
    .X(_0311_));
 sky130_fd_sc_hd__buf_2 _1232_ (.A(net1417),
    .X(net470));
 sky130_fd_sc_hd__and3b_1 _1233_ (.A_N(net268),
    .B(net2739),
    .C(net12),
    .X(_0312_));
 sky130_fd_sc_hd__clkbuf_1 _1234_ (.A(net1415),
    .X(net471));
 sky130_fd_sc_hd__and3b_1 _1235_ (.A_N(net1961),
    .B(net2736),
    .C(net13),
    .X(_0313_));
 sky130_fd_sc_hd__buf_2 _1236_ (.A(net1414),
    .X(net472));
 sky130_fd_sc_hd__and3b_2 _1237_ (.A_N(net270),
    .B(net2734),
    .C(net14),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_1 _1238_ (.A(net1413),
    .X(net473));
 sky130_fd_sc_hd__and3b_1 _1239_ (.A_N(net1958),
    .B(net2732),
    .C(net16),
    .X(_0315_));
 sky130_fd_sc_hd__buf_2 _1240_ (.A(net1412),
    .X(net475));
 sky130_fd_sc_hd__and3b_1 _1241_ (.A_N(net1957),
    .B(net2729),
    .C(net2007),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_2 _1242_ (.A(_0316_),
    .X(net476));
 sky130_fd_sc_hd__and3b_1 _1243_ (.A_N(net1956),
    .B(net2727),
    .C(net18),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_2 _1244_ (.A(net1411),
    .X(net477));
 sky130_fd_sc_hd__and3b_1 _1245_ (.A_N(net1955),
    .B(net2725),
    .C(net19),
    .X(_0318_));
 sky130_fd_sc_hd__clkbuf_2 _1246_ (.A(_0318_),
    .X(net478));
 sky130_fd_sc_hd__and3b_1 _1247_ (.A_N(net1954),
    .B(net2722),
    .C(net20),
    .X(_0319_));
 sky130_fd_sc_hd__clkbuf_2 _1248_ (.A(net1410),
    .X(net479));
 sky130_fd_sc_hd__and3b_1 _1249_ (.A_N(net1952),
    .B(net2719),
    .C(net21),
    .X(_0320_));
 sky130_fd_sc_hd__clkbuf_2 _1250_ (.A(net1409),
    .X(net480));
 sky130_fd_sc_hd__and3b_1 _1251_ (.A_N(net1951),
    .B(net2716),
    .C(net22),
    .X(_0321_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1252_ (.A(_0321_),
    .X(net481));
 sky130_fd_sc_hd__and3b_1 _1253_ (.A_N(net1950),
    .B(net2714),
    .C(net23),
    .X(_0322_));
 sky130_fd_sc_hd__clkbuf_2 _1254_ (.A(net1408),
    .X(net482));
 sky130_fd_sc_hd__and3b_1 _1255_ (.A_N(net1948),
    .B(net2711),
    .C(net24),
    .X(_0323_));
 sky130_fd_sc_hd__clkbuf_2 _1256_ (.A(net1407),
    .X(net483));
 sky130_fd_sc_hd__and3b_1 _1257_ (.A_N(net281),
    .B(net2708),
    .C(net25),
    .X(_0324_));
 sky130_fd_sc_hd__clkbuf_2 _1258_ (.A(net1406),
    .X(net484));
 sky130_fd_sc_hd__and3b_2 _1259_ (.A_N(net1946),
    .B(net2705),
    .C(net1960),
    .X(_0325_));
 sky130_fd_sc_hd__clkbuf_2 _1260_ (.A(_0325_),
    .X(net486));
 sky130_fd_sc_hd__and3b_1 _1261_ (.A_N(net1944),
    .B(net2701),
    .C(net1949),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_2 _1262_ (.A(_0326_),
    .X(net487));
 sky130_fd_sc_hd__and3b_1 _1263_ (.A_N(net285),
    .B(net2698),
    .C(net29),
    .X(_0327_));
 sky130_fd_sc_hd__clkbuf_2 _1264_ (.A(net1405),
    .X(net488));
 sky130_fd_sc_hd__and3b_2 _1265_ (.A_N(net286),
    .B(net2695),
    .C(net30),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_2 _1266_ (.A(_0328_),
    .X(net489));
 sky130_fd_sc_hd__and3b_1 _1267_ (.A_N(net1941),
    .B(net2691),
    .C(net1923),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_2 _1268_ (.A(_0329_),
    .X(net490));
 sky130_fd_sc_hd__and3b_1 _1269_ (.A_N(net1940),
    .B(net2687),
    .C(net1919),
    .X(_0330_));
 sky130_fd_sc_hd__clkbuf_2 _1270_ (.A(_0330_),
    .X(net491));
 sky130_fd_sc_hd__and3b_1 _1271_ (.A_N(net1939),
    .B(net2683),
    .C(net1907),
    .X(_0331_));
 sky130_fd_sc_hd__clkbuf_2 _1272_ (.A(_0331_),
    .X(net492));
 sky130_fd_sc_hd__and3b_1 _1273_ (.A_N(net1938),
    .B(net2680),
    .C(net1894),
    .X(_0332_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1274_ (.A(_0332_),
    .X(net493));
 sky130_fd_sc_hd__and2_1 _1275_ (.A(net260),
    .B(net2678),
    .X(_0333_));
 sky130_fd_sc_hd__clkbuf_1 _1276_ (.A(_0333_),
    .X(net719));
 sky130_fd_sc_hd__and2_2 _1277_ (.A(net299),
    .B(net2675),
    .X(_0334_));
 sky130_fd_sc_hd__buf_2 _1278_ (.A(_0334_),
    .X(net758));
 sky130_fd_sc_hd__and2_1 _1279_ (.A(net310),
    .B(net2672),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_2 _1280_ (.A(net1404),
    .X(net769));
 sky130_fd_sc_hd__and2_1 _1281_ (.A(net321),
    .B(net2669),
    .X(_0336_));
 sky130_fd_sc_hd__clkbuf_2 _1282_ (.A(net1403),
    .X(net780));
 sky130_fd_sc_hd__and2_1 _1283_ (.A(net332),
    .B(net2667),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _1284_ (.A(net1402),
    .X(net791));
 sky130_fd_sc_hd__and2_2 _1285_ (.A(net343),
    .B(net2664),
    .X(_0338_));
 sky130_fd_sc_hd__clkbuf_2 _1286_ (.A(net1401),
    .X(net802));
 sky130_fd_sc_hd__and2_1 _1287_ (.A(net354),
    .B(net2661),
    .X(_0339_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1288_ (.A(net1399),
    .X(net813));
 sky130_fd_sc_hd__and2_1 _1289_ (.A(net365),
    .B(net2659),
    .X(_0340_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1290_ (.A(net1397),
    .X(net824));
 sky130_fd_sc_hd__and2_1 _1291_ (.A(net376),
    .B(net2657),
    .X(_0341_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1292_ (.A(net1395),
    .X(net835));
 sky130_fd_sc_hd__and2_1 _1293_ (.A(net387),
    .B(net2654),
    .X(_0342_));
 sky130_fd_sc_hd__clkbuf_1 _1294_ (.A(net1393),
    .X(net846));
 sky130_fd_sc_hd__and2_2 _1295_ (.A(net271),
    .B(net2651),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _1296_ (.A(net1392),
    .X(net730));
 sky130_fd_sc_hd__and2_1 _1297_ (.A(net282),
    .B(net2649),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_2 _1298_ (.A(net1391),
    .X(net741));
 sky130_fd_sc_hd__and2_1 _1299_ (.A(net291),
    .B(net2648),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_1 _1300_ (.A(net1390),
    .X(net750));
 sky130_fd_sc_hd__and2_1 _1301_ (.A(net292),
    .B(net2645),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_1 _1302_ (.A(net1388),
    .X(net751));
 sky130_fd_sc_hd__and2_1 _1303_ (.A(net293),
    .B(net2642),
    .X(_0347_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1304_ (.A(net1387),
    .X(net752));
 sky130_fd_sc_hd__and2_2 _1305_ (.A(net294),
    .B(net2640),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _1306_ (.A(net1386),
    .X(net753));
 sky130_fd_sc_hd__and2_1 _1307_ (.A(net295),
    .B(net2638),
    .X(_0349_));
 sky130_fd_sc_hd__clkbuf_1 _1308_ (.A(net1385),
    .X(net754));
 sky130_fd_sc_hd__and2_1 _1309_ (.A(net296),
    .B(net2636),
    .X(_0350_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1310_ (.A(net1383),
    .X(net755));
 sky130_fd_sc_hd__and2_2 _1311_ (.A(net1937),
    .B(net2632),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_2 _1312_ (.A(net1382),
    .X(net756));
 sky130_fd_sc_hd__and2_1 _1313_ (.A(net298),
    .B(net2630),
    .X(_0352_));
 sky130_fd_sc_hd__clkbuf_2 _1314_ (.A(net1381),
    .X(net757));
 sky130_fd_sc_hd__and2_1 _1315_ (.A(net1929),
    .B(net2628),
    .X(_0353_));
 sky130_fd_sc_hd__clkbuf_2 _1316_ (.A(net1379),
    .X(net759));
 sky130_fd_sc_hd__and2_1 _1317_ (.A(net301),
    .B(net2627),
    .X(_0354_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1318_ (.A(net1378),
    .X(net760));
 sky130_fd_sc_hd__and2_1 _1319_ (.A(net302),
    .B(net2626),
    .X(_0355_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1320_ (.A(net1377),
    .X(net761));
 sky130_fd_sc_hd__and2_1 _1321_ (.A(net303),
    .B(net2623),
    .X(_0356_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1322_ (.A(net1375),
    .X(net762));
 sky130_fd_sc_hd__and2_1 _1323_ (.A(net304),
    .B(net2622),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_1 _1324_ (.A(net1374),
    .X(net763));
 sky130_fd_sc_hd__and2_1 _1325_ (.A(net305),
    .B(net2620),
    .X(_0358_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1326_ (.A(net1372),
    .X(net764));
 sky130_fd_sc_hd__and2_1 _1327_ (.A(net1927),
    .B(\mprj_logic1[228] ),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _1328_ (.A(_0359_),
    .X(net765));
 sky130_fd_sc_hd__and2_1 _1329_ (.A(net1926),
    .B(net2618),
    .X(_0360_));
 sky130_fd_sc_hd__clkbuf_1 _1330_ (.A(net1371),
    .X(net766));
 sky130_fd_sc_hd__and2_1 _1331_ (.A(net308),
    .B(net2617),
    .X(_0361_));
 sky130_fd_sc_hd__clkbuf_1 _1332_ (.A(net1369),
    .X(net767));
 sky130_fd_sc_hd__and2_1 _1333_ (.A(net1925),
    .B(net2616),
    .X(_0362_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1334_ (.A(_0362_),
    .X(net768));
 sky130_fd_sc_hd__and2_1 _1335_ (.A(net311),
    .B(net2615),
    .X(_0363_));
 sky130_fd_sc_hd__clkbuf_1 _1336_ (.A(net1368),
    .X(net770));
 sky130_fd_sc_hd__and2_1 _1337_ (.A(net312),
    .B(net2613),
    .X(_0364_));
 sky130_fd_sc_hd__clkbuf_1 _1338_ (.A(net1367),
    .X(net771));
 sky130_fd_sc_hd__and2_1 _1339_ (.A(net313),
    .B(net2612),
    .X(_0365_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1340_ (.A(net1366),
    .X(net772));
 sky130_fd_sc_hd__and2_1 _1341_ (.A(net314),
    .B(net2611),
    .X(_0366_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1342_ (.A(net1365),
    .X(net773));
 sky130_fd_sc_hd__and2_1 _1343_ (.A(net315),
    .B(net2610),
    .X(_0367_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1344_ (.A(net1364),
    .X(net774));
 sky130_fd_sc_hd__and2_1 _1345_ (.A(net1922),
    .B(\mprj_logic1[237] ),
    .X(_0368_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1346_ (.A(_0368_),
    .X(net775));
 sky130_fd_sc_hd__and2_1 _1347_ (.A(net317),
    .B(net2609),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_2 _1348_ (.A(net1363),
    .X(net776));
 sky130_fd_sc_hd__and2_1 _1349_ (.A(net1920),
    .B(\mprj_logic1[239] ),
    .X(_0370_));
 sky130_fd_sc_hd__clkbuf_1 _1350_ (.A(net1362),
    .X(net777));
 sky130_fd_sc_hd__and2_1 _1351_ (.A(net319),
    .B(\mprj_logic1[240] ),
    .X(_0371_));
 sky130_fd_sc_hd__clkbuf_1 _1352_ (.A(net1361),
    .X(net778));
 sky130_fd_sc_hd__and2_1 _1353_ (.A(net320),
    .B(\mprj_logic1[241] ),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _1354_ (.A(_0372_),
    .X(net779));
 sky130_fd_sc_hd__and2_1 _1355_ (.A(net1917),
    .B(\mprj_logic1[242] ),
    .X(_0373_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1356_ (.A(_0373_),
    .X(net781));
 sky130_fd_sc_hd__and2_1 _1357_ (.A(net1916),
    .B(net2608),
    .X(_0374_));
 sky130_fd_sc_hd__clkbuf_2 _1358_ (.A(net1359),
    .X(net782));
 sky130_fd_sc_hd__and2_1 _1359_ (.A(net324),
    .B(\mprj_logic1[244] ),
    .X(_0375_));
 sky130_fd_sc_hd__buf_2 _1360_ (.A(_0375_),
    .X(net783));
 sky130_fd_sc_hd__and2_1 _1361_ (.A(net1914),
    .B(\mprj_logic1[245] ),
    .X(_0376_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1362_ (.A(_0376_),
    .X(net784));
 sky130_fd_sc_hd__and2_1 _1363_ (.A(net326),
    .B(\mprj_logic1[246] ),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_2 _1364_ (.A(net1358),
    .X(net785));
 sky130_fd_sc_hd__and2_1 _1365_ (.A(net327),
    .B(\mprj_logic1[247] ),
    .X(_0378_));
 sky130_fd_sc_hd__clkbuf_1 _1366_ (.A(_0378_),
    .X(net786));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(net1911),
    .B(net2607),
    .X(_0379_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1368_ (.A(net1357),
    .X(net787));
 sky130_fd_sc_hd__and2_2 _1369_ (.A(net1908),
    .B(\mprj_logic1[249] ),
    .X(_0380_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1370_ (.A(_0380_),
    .X(net788));
 sky130_fd_sc_hd__and2_2 _1371_ (.A(net1904),
    .B(net2606),
    .X(_0381_));
 sky130_fd_sc_hd__clkbuf_2 _1372_ (.A(_0381_),
    .X(net789));
 sky130_fd_sc_hd__and2_1 _1373_ (.A(net331),
    .B(\mprj_logic1[251] ),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_2 _1374_ (.A(_0382_),
    .X(net790));
 sky130_fd_sc_hd__and2_1 _1375_ (.A(net1903),
    .B(net2605),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_2 _1376_ (.A(net1355),
    .X(net792));
 sky130_fd_sc_hd__and2_1 _1377_ (.A(net1901),
    .B(\mprj_logic1[253] ),
    .X(_0384_));
 sky130_fd_sc_hd__clkbuf_2 _1378_ (.A(_0384_),
    .X(net793));
 sky130_fd_sc_hd__and2_1 _1379_ (.A(net1900),
    .B(net2604),
    .X(_0385_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1380_ (.A(net1353),
    .X(net794));
 sky130_fd_sc_hd__and2_1 _1381_ (.A(net1899),
    .B(net2603),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_2 _1382_ (.A(net1351),
    .X(net795));
 sky130_fd_sc_hd__and2_1 _1383_ (.A(net1897),
    .B(\mprj_logic1[256] ),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_1 _1384_ (.A(_0387_),
    .X(net796));
 sky130_fd_sc_hd__and2_1 _1385_ (.A(net1895),
    .B(net2602),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_1 _1386_ (.A(net1349),
    .X(net797));
 sky130_fd_sc_hd__and2_1 _1387_ (.A(net339),
    .B(\mprj_logic1[258] ),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_2 _1388_ (.A(net1348),
    .X(net798));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(net1892),
    .B(net2601),
    .X(_0390_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1390_ (.A(_0390_),
    .X(net799));
 sky130_fd_sc_hd__and2_1 _1391_ (.A(net1890),
    .B(\mprj_logic1[260] ),
    .X(_0391_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1392_ (.A(net1346),
    .X(net800));
 sky130_fd_sc_hd__and2_1 _1393_ (.A(net1887),
    .B(net2600),
    .X(_0392_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1394_ (.A(_0392_),
    .X(net801));
 sky130_fd_sc_hd__and2_1 _1395_ (.A(net1886),
    .B(\mprj_logic1[262] ),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_2 _1396_ (.A(net1344),
    .X(net803));
 sky130_fd_sc_hd__and2_2 _1397_ (.A(net1885),
    .B(\mprj_logic1[263] ),
    .X(_0394_));
 sky130_fd_sc_hd__clkbuf_1 _1398_ (.A(net1342),
    .X(net804));
 sky130_fd_sc_hd__and2_1 _1399_ (.A(net1884),
    .B(\mprj_logic1[264] ),
    .X(_0395_));
 sky130_fd_sc_hd__clkbuf_1 _1400_ (.A(net1340),
    .X(net805));
 sky130_fd_sc_hd__and2_1 _1401_ (.A(net1883),
    .B(\mprj_logic1[265] ),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_2 _1402_ (.A(net1339),
    .X(net806));
 sky130_fd_sc_hd__and2_1 _1403_ (.A(net1880),
    .B(net2599),
    .X(_0397_));
 sky130_fd_sc_hd__clkbuf_2 _1404_ (.A(_0397_),
    .X(net807));
 sky130_fd_sc_hd__and2_2 _1405_ (.A(net1879),
    .B(\mprj_logic1[267] ),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_1 _1406_ (.A(net1337),
    .X(net808));
 sky130_fd_sc_hd__and2_1 _1407_ (.A(net1877),
    .B(net2598),
    .X(_0399_));
 sky130_fd_sc_hd__clkbuf_2 _1408_ (.A(net1336),
    .X(net809));
 sky130_fd_sc_hd__and2_1 _1409_ (.A(net1876),
    .B(\mprj_logic1[269] ),
    .X(_0400_));
 sky130_fd_sc_hd__buf_2 _1410_ (.A(_0400_),
    .X(net810));
 sky130_fd_sc_hd__and2_1 _1411_ (.A(net1875),
    .B(net2595),
    .X(_0401_));
 sky130_fd_sc_hd__clkbuf_1 _1412_ (.A(_0401_),
    .X(net811));
 sky130_fd_sc_hd__and2_1 _1413_ (.A(net1874),
    .B(net2594),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_1 _1414_ (.A(_0402_),
    .X(net812));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(net1873),
    .B(net2593),
    .X(_0403_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1416_ (.A(_0403_),
    .X(net814));
 sky130_fd_sc_hd__and2_1 _1417_ (.A(net1872),
    .B(net2591),
    .X(_0404_));
 sky130_fd_sc_hd__clkbuf_1 _1418_ (.A(_0404_),
    .X(net815));
 sky130_fd_sc_hd__and2_1 _1419_ (.A(net1871),
    .B(net2589),
    .X(_0405_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1420_ (.A(_0405_),
    .X(net816));
 sky130_fd_sc_hd__and2_1 _1421_ (.A(net1870),
    .B(net2588),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _1422_ (.A(net1335),
    .X(net817));
 sky130_fd_sc_hd__and2_1 _1423_ (.A(net1868),
    .B(net2586),
    .X(_0407_));
 sky130_fd_sc_hd__buf_2 _1424_ (.A(_0407_),
    .X(net818));
 sky130_fd_sc_hd__and2_1 _1425_ (.A(net1867),
    .B(net2584),
    .X(_0408_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1426_ (.A(_0408_),
    .X(net819));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(net1865),
    .B(net2581),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_2 _1428_ (.A(_0409_),
    .X(net820));
 sky130_fd_sc_hd__and2_2 _1429_ (.A(net1863),
    .B(net2578),
    .X(_0410_));
 sky130_fd_sc_hd__clkbuf_2 _1430_ (.A(_0410_),
    .X(net821));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(net1861),
    .B(net2575),
    .X(_0411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1432_ (.A(_0411_),
    .X(net822));
 sky130_fd_sc_hd__and2_1 _1433_ (.A(net1859),
    .B(net2573),
    .X(_0412_));
 sky130_fd_sc_hd__clkbuf_2 _1434_ (.A(_0412_),
    .X(net823));
 sky130_fd_sc_hd__and2_1 _1435_ (.A(net1857),
    .B(net2570),
    .X(_0413_));
 sky130_fd_sc_hd__buf_2 _1436_ (.A(_0413_),
    .X(net825));
 sky130_fd_sc_hd__and2_1 _1437_ (.A(net1855),
    .B(net2568),
    .X(_0414_));
 sky130_fd_sc_hd__clkbuf_1 _1438_ (.A(_0414_),
    .X(net826));
 sky130_fd_sc_hd__and2_1 _1439_ (.A(net1853),
    .B(net2564),
    .X(_0415_));
 sky130_fd_sc_hd__clkbuf_2 _1440_ (.A(net1334),
    .X(net827));
 sky130_fd_sc_hd__and2_1 _1441_ (.A(net1851),
    .B(net2561),
    .X(_0416_));
 sky130_fd_sc_hd__clkbuf_2 _1442_ (.A(_0416_),
    .X(net828));
 sky130_fd_sc_hd__and2_2 _1443_ (.A(net1849),
    .B(net2558),
    .X(_0417_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1444_ (.A(_0417_),
    .X(net829));
 sky130_fd_sc_hd__and2_1 _1445_ (.A(net1847),
    .B(net2555),
    .X(_0418_));
 sky130_fd_sc_hd__clkbuf_2 _1446_ (.A(_0418_),
    .X(net830));
 sky130_fd_sc_hd__and2_1 _1447_ (.A(net1845),
    .B(net2551),
    .X(_0419_));
 sky130_fd_sc_hd__clkbuf_2 _1448_ (.A(_0419_),
    .X(net831));
 sky130_fd_sc_hd__and2_1 _1449_ (.A(net1843),
    .B(net2548),
    .X(_0420_));
 sky130_fd_sc_hd__clkbuf_1 _1450_ (.A(_0420_),
    .X(net832));
 sky130_fd_sc_hd__and2_1 _1451_ (.A(net1841),
    .B(net2544),
    .X(_0421_));
 sky130_fd_sc_hd__clkbuf_1 _1452_ (.A(_0421_),
    .X(net833));
 sky130_fd_sc_hd__and2_1 _1453_ (.A(net375),
    .B(net2543),
    .X(_0422_));
 sky130_fd_sc_hd__clkbuf_1 _1454_ (.A(net1333),
    .X(net834));
 sky130_fd_sc_hd__and2_1 _1455_ (.A(net377),
    .B(net2542),
    .X(_0423_));
 sky130_fd_sc_hd__clkbuf_1 _1456_ (.A(net1331),
    .X(net836));
 sky130_fd_sc_hd__and2_1 _1457_ (.A(net378),
    .B(net2541),
    .X(_0424_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1458_ (.A(net1330),
    .X(net837));
 sky130_fd_sc_hd__and2_1 _1459_ (.A(net379),
    .B(\mprj_logic1[294] ),
    .X(_0425_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1460_ (.A(net1329),
    .X(net838));
 sky130_fd_sc_hd__and2_1 _1461_ (.A(net1840),
    .B(net2539),
    .X(_0426_));
 sky130_fd_sc_hd__clkbuf_2 _1462_ (.A(_0426_),
    .X(net839));
 sky130_fd_sc_hd__and2_1 _1463_ (.A(net1839),
    .B(net2537),
    .X(_0427_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1464_ (.A(_0427_),
    .X(net840));
 sky130_fd_sc_hd__and2_1 _1465_ (.A(net1838),
    .B(net2534),
    .X(_0428_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1466_ (.A(_0428_),
    .X(net841));
 sky130_fd_sc_hd__and2_1 _1467_ (.A(net1836),
    .B(net2531),
    .X(_0429_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1468_ (.A(_0429_),
    .X(net842));
 sky130_fd_sc_hd__and2_1 _1469_ (.A(net1835),
    .B(net2529),
    .X(_0430_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1470_ (.A(_0430_),
    .X(net843));
 sky130_fd_sc_hd__and2_1 _1471_ (.A(net1833),
    .B(net2521),
    .X(_0431_));
 sky130_fd_sc_hd__clkbuf_2 _1472_ (.A(_0431_),
    .X(net844));
 sky130_fd_sc_hd__and2_1 _1473_ (.A(net1831),
    .B(net2518),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _1474_ (.A(_0432_),
    .X(net845));
 sky130_fd_sc_hd__and2_1 _1475_ (.A(net1972),
    .B(net2515),
    .X(_0433_));
 sky130_fd_sc_hd__clkbuf_2 _1476_ (.A(_0433_),
    .X(net720));
 sky130_fd_sc_hd__and2_1 _1477_ (.A(net1971),
    .B(net2512),
    .X(_0434_));
 sky130_fd_sc_hd__clkbuf_2 _1478_ (.A(_0434_),
    .X(net721));
 sky130_fd_sc_hd__and2_1 _1479_ (.A(net1969),
    .B(net2509),
    .X(_0435_));
 sky130_fd_sc_hd__clkbuf_2 _1480_ (.A(_0435_),
    .X(net722));
 sky130_fd_sc_hd__and2_1 _1481_ (.A(net1968),
    .B(net2506),
    .X(_0436_));
 sky130_fd_sc_hd__clkbuf_2 _1482_ (.A(_0436_),
    .X(net723));
 sky130_fd_sc_hd__and2_1 _1483_ (.A(net1967),
    .B(net2504),
    .X(_0437_));
 sky130_fd_sc_hd__clkbuf_2 _1484_ (.A(_0437_),
    .X(net724));
 sky130_fd_sc_hd__and2_1 _1485_ (.A(net1965),
    .B(net2501),
    .X(_0438_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1486_ (.A(_0438_),
    .X(net725));
 sky130_fd_sc_hd__and2_1 _1487_ (.A(net1963),
    .B(net2498),
    .X(_0439_));
 sky130_fd_sc_hd__clkbuf_2 _1488_ (.A(_0439_),
    .X(net726));
 sky130_fd_sc_hd__and2_1 _1489_ (.A(net1962),
    .B(net2495),
    .X(_0440_));
 sky130_fd_sc_hd__clkbuf_2 _1490_ (.A(_0440_),
    .X(net727));
 sky130_fd_sc_hd__and2_1 _1491_ (.A(net1961),
    .B(net2492),
    .X(_0441_));
 sky130_fd_sc_hd__clkbuf_2 _1492_ (.A(_0441_),
    .X(net728));
 sky130_fd_sc_hd__and2_1 _1493_ (.A(net1959),
    .B(net2489),
    .X(_0442_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1494_ (.A(_0442_),
    .X(net729));
 sky130_fd_sc_hd__and2_1 _1495_ (.A(net1958),
    .B(net2485),
    .X(_0443_));
 sky130_fd_sc_hd__clkbuf_2 _1496_ (.A(_0443_),
    .X(net731));
 sky130_fd_sc_hd__and2_1 _1497_ (.A(net1957),
    .B(net2482),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_2 _1498_ (.A(_0444_),
    .X(net732));
 sky130_fd_sc_hd__and2_1 _1499_ (.A(net1956),
    .B(net2480),
    .X(_0445_));
 sky130_fd_sc_hd__clkbuf_2 _1500_ (.A(_0445_),
    .X(net733));
 sky130_fd_sc_hd__and2_1 _1501_ (.A(net1955),
    .B(net2477),
    .X(_0446_));
 sky130_fd_sc_hd__buf_2 _1502_ (.A(_0446_),
    .X(net734));
 sky130_fd_sc_hd__and2_1 _1503_ (.A(net1953),
    .B(net2473),
    .X(_0447_));
 sky130_fd_sc_hd__clkbuf_2 _1504_ (.A(_0447_),
    .X(net735));
 sky130_fd_sc_hd__and2_1 _1505_ (.A(net1952),
    .B(net2469),
    .X(_0448_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1506_ (.A(_0448_),
    .X(net736));
 sky130_fd_sc_hd__and2_1 _1507_ (.A(net1951),
    .B(net2466),
    .X(_0449_));
 sky130_fd_sc_hd__clkbuf_2 _1508_ (.A(_0449_),
    .X(net737));
 sky130_fd_sc_hd__and2_1 _1509_ (.A(net1950),
    .B(net2463),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_1 _1510_ (.A(_0450_),
    .X(net738));
 sky130_fd_sc_hd__and2_1 _1511_ (.A(net1948),
    .B(net2459),
    .X(_0451_));
 sky130_fd_sc_hd__clkbuf_2 _1512_ (.A(_0451_),
    .X(net739));
 sky130_fd_sc_hd__and2_1 _1513_ (.A(net1947),
    .B(net2455),
    .X(_0452_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1514_ (.A(_0452_),
    .X(net740));
 sky130_fd_sc_hd__and2_1 _1515_ (.A(net1945),
    .B(net2451),
    .X(_0453_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1516_ (.A(_0453_),
    .X(net742));
 sky130_fd_sc_hd__and2_1 _1517_ (.A(net1944),
    .B(net2447),
    .X(_0454_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1518_ (.A(_0454_),
    .X(net743));
 sky130_fd_sc_hd__and2_1 _1519_ (.A(net1943),
    .B(net2443),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_2 _1520_ (.A(_0455_),
    .X(net744));
 sky130_fd_sc_hd__and2_1 _1521_ (.A(net1942),
    .B(net2439),
    .X(_0456_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1522_ (.A(_0456_),
    .X(net745));
 sky130_fd_sc_hd__and2_1 _1523_ (.A(net1941),
    .B(net2435),
    .X(_0457_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1524_ (.A(_0457_),
    .X(net746));
 sky130_fd_sc_hd__and2_1 _1525_ (.A(net1940),
    .B(net2431),
    .X(_0458_));
 sky130_fd_sc_hd__clkbuf_1 _1526_ (.A(_0458_),
    .X(net747));
 sky130_fd_sc_hd__and2_2 _1527_ (.A(net1939),
    .B(net2427),
    .X(_0459_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1528_ (.A(_0459_),
    .X(net748));
 sky130_fd_sc_hd__and2_1 _1529_ (.A(net1938),
    .B(net2422),
    .X(_0460_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1530_ (.A(_0460_),
    .X(net749));
 sky130_fd_sc_hd__and2_1 _1531_ (.A(net2420),
    .B(net132),
    .X(_0461_));
 sky130_fd_sc_hd__clkbuf_1 _1532_ (.A(_0461_),
    .X(\la_data_in_enable[0] ));
 sky130_fd_sc_hd__inv_2 _1533_ (.A(\la_data_in_mprj_bar[0] ),
    .Y(net591));
 sky130_fd_sc_hd__inv_2 _1534_ (.A(\la_data_in_mprj_bar[1] ),
    .Y(net630));
 sky130_fd_sc_hd__inv_2 _1535_ (.A(\la_data_in_mprj_bar[2] ),
    .Y(net641));
 sky130_fd_sc_hd__inv_2 _1536_ (.A(\la_data_in_mprj_bar[3] ),
    .Y(net652));
 sky130_fd_sc_hd__inv_2 _1537_ (.A(\la_data_in_mprj_bar[4] ),
    .Y(net663));
 sky130_fd_sc_hd__inv_2 _1538_ (.A(\la_data_in_mprj_bar[5] ),
    .Y(net674));
 sky130_fd_sc_hd__inv_2 _1539_ (.A(\la_data_in_mprj_bar[6] ),
    .Y(net685));
 sky130_fd_sc_hd__clkinv_2 _1540_ (.A(\la_data_in_mprj_bar[7] ),
    .Y(net696));
 sky130_fd_sc_hd__clkinv_2 _1541_ (.A(\la_data_in_mprj_bar[8] ),
    .Y(net707));
 sky130_fd_sc_hd__clkinv_2 _1542_ (.A(\la_data_in_mprj_bar[9] ),
    .Y(net718));
 sky130_fd_sc_hd__inv_2 _1543_ (.A(\la_data_in_mprj_bar[10] ),
    .Y(net602));
 sky130_fd_sc_hd__inv_2 _1544_ (.A(\la_data_in_mprj_bar[11] ),
    .Y(net613));
 sky130_fd_sc_hd__inv_2 _1545_ (.A(\la_data_in_mprj_bar[12] ),
    .Y(net622));
 sky130_fd_sc_hd__clkinv_2 _1546_ (.A(\la_data_in_mprj_bar[13] ),
    .Y(net623));
 sky130_fd_sc_hd__clkinv_2 _1547_ (.A(\la_data_in_mprj_bar[14] ),
    .Y(net624));
 sky130_fd_sc_hd__inv_2 _1548_ (.A(\la_data_in_mprj_bar[15] ),
    .Y(net625));
 sky130_fd_sc_hd__clkinv_2 _1549_ (.A(\la_data_in_mprj_bar[16] ),
    .Y(net626));
 mprj2_logic_high mprj2_logic_high_inst (.HI(net953));
 mprj_logic_high mprj_logic_high_inst (.HI({\mprj_logic1[462] ,
    net951,
    \mprj_logic1[460] ,
    \mprj_logic1[459] ,
    \mprj_logic1[458] ,
    \mprj_logic1[457] ,
    \mprj_logic1[456] ,
    \mprj_logic1[455] ,
    \mprj_logic1[454] ,
    \mprj_logic1[453] ,
    \mprj_logic1[452] ,
    \mprj_logic1[451] ,
    \mprj_logic1[450] ,
    \mprj_logic1[449] ,
    \mprj_logic1[448] ,
    \mprj_logic1[447] ,
    \mprj_logic1[446] ,
    \mprj_logic1[445] ,
    \mprj_logic1[444] ,
    \mprj_logic1[443] ,
    \mprj_logic1[442] ,
    \mprj_logic1[441] ,
    \mprj_logic1[440] ,
    \mprj_logic1[439] ,
    \mprj_logic1[438] ,
    \mprj_logic1[437] ,
    \mprj_logic1[436] ,
    \mprj_logic1[435] ,
    \mprj_logic1[434] ,
    \mprj_logic1[433] ,
    \mprj_logic1[432] ,
    \mprj_logic1[431] ,
    \mprj_logic1[430] ,
    \mprj_logic1[429] ,
    \mprj_logic1[428] ,
    \mprj_logic1[427] ,
    \mprj_logic1[426] ,
    \mprj_logic1[425] ,
    \mprj_logic1[424] ,
    \mprj_logic1[423] ,
    \mprj_logic1[422] ,
    \mprj_logic1[421] ,
    \mprj_logic1[420] ,
    \mprj_logic1[419] ,
    \mprj_logic1[418] ,
    \mprj_logic1[417] ,
    \mprj_logic1[416] ,
    \mprj_logic1[415] ,
    \mprj_logic1[414] ,
    \mprj_logic1[413] ,
    \mprj_logic1[412] ,
    \mprj_logic1[411] ,
    \mprj_logic1[410] ,
    \mprj_logic1[409] ,
    \mprj_logic1[408] ,
    \mprj_logic1[407] ,
    \mprj_logic1[406] ,
    \mprj_logic1[405] ,
    \mprj_logic1[404] ,
    \mprj_logic1[403] ,
    \mprj_logic1[402] ,
    \mprj_logic1[401] ,
    \mprj_logic1[400] ,
    \mprj_logic1[399] ,
    \mprj_logic1[398] ,
    \mprj_logic1[397] ,
    \mprj_logic1[396] ,
    \mprj_logic1[395] ,
    \mprj_logic1[394] ,
    \mprj_logic1[393] ,
    \mprj_logic1[392] ,
    \mprj_logic1[391] ,
    \mprj_logic1[390] ,
    \mprj_logic1[389] ,
    \mprj_logic1[388] ,
    \mprj_logic1[387] ,
    \mprj_logic1[386] ,
    \mprj_logic1[385] ,
    \mprj_logic1[384] ,
    \mprj_logic1[383] ,
    \mprj_logic1[382] ,
    \mprj_logic1[381] ,
    \mprj_logic1[380] ,
    \mprj_logic1[379] ,
    \mprj_logic1[378] ,
    \mprj_logic1[377] ,
    \mprj_logic1[376] ,
    \mprj_logic1[375] ,
    \mprj_logic1[374] ,
    \mprj_logic1[373] ,
    \mprj_logic1[372] ,
    \mprj_logic1[371] ,
    \mprj_logic1[370] ,
    \mprj_logic1[369] ,
    \mprj_logic1[368] ,
    \mprj_logic1[367] ,
    \mprj_logic1[366] ,
    \mprj_logic1[365] ,
    \mprj_logic1[364] ,
    \mprj_logic1[363] ,
    \mprj_logic1[362] ,
    \mprj_logic1[361] ,
    \mprj_logic1[360] ,
    \mprj_logic1[359] ,
    \mprj_logic1[358] ,
    \mprj_logic1[357] ,
    \mprj_logic1[356] ,
    \mprj_logic1[355] ,
    \mprj_logic1[354] ,
    \mprj_logic1[353] ,
    \mprj_logic1[352] ,
    \mprj_logic1[351] ,
    \mprj_logic1[350] ,
    \mprj_logic1[349] ,
    \mprj_logic1[348] ,
    \mprj_logic1[347] ,
    \mprj_logic1[346] ,
    \mprj_logic1[345] ,
    \mprj_logic1[344] ,
    \mprj_logic1[343] ,
    \mprj_logic1[342] ,
    \mprj_logic1[341] ,
    \mprj_logic1[340] ,
    \mprj_logic1[339] ,
    \mprj_logic1[338] ,
    \mprj_logic1[337] ,
    \mprj_logic1[336] ,
    \mprj_logic1[335] ,
    \mprj_logic1[334] ,
    \mprj_logic1[333] ,
    \mprj_logic1[332] ,
    \mprj_logic1[331] ,
    \mprj_logic1[330] ,
    \mprj_logic1[329] ,
    \mprj_logic1[328] ,
    \mprj_logic1[327] ,
    \mprj_logic1[326] ,
    \mprj_logic1[325] ,
    \mprj_logic1[324] ,
    \mprj_logic1[323] ,
    \mprj_logic1[322] ,
    \mprj_logic1[321] ,
    \mprj_logic1[320] ,
    \mprj_logic1[319] ,
    \mprj_logic1[318] ,
    \mprj_logic1[317] ,
    \mprj_logic1[316] ,
    \mprj_logic1[315] ,
    \mprj_logic1[314] ,
    \mprj_logic1[313] ,
    \mprj_logic1[312] ,
    \mprj_logic1[311] ,
    \mprj_logic1[310] ,
    \mprj_logic1[309] ,
    \mprj_logic1[308] ,
    \mprj_logic1[307] ,
    \mprj_logic1[306] ,
    \mprj_logic1[305] ,
    \mprj_logic1[304] ,
    \mprj_logic1[303] ,
    \mprj_logic1[302] ,
    \mprj_logic1[301] ,
    \mprj_logic1[300] ,
    \mprj_logic1[299] ,
    \mprj_logic1[298] ,
    \mprj_logic1[297] ,
    \mprj_logic1[296] ,
    \mprj_logic1[295] ,
    \mprj_logic1[294] ,
    \mprj_logic1[293] ,
    \mprj_logic1[292] ,
    \mprj_logic1[291] ,
    \mprj_logic1[290] ,
    \mprj_logic1[289] ,
    \mprj_logic1[288] ,
    \mprj_logic1[287] ,
    \mprj_logic1[286] ,
    \mprj_logic1[285] ,
    \mprj_logic1[284] ,
    \mprj_logic1[283] ,
    \mprj_logic1[282] ,
    \mprj_logic1[281] ,
    \mprj_logic1[280] ,
    \mprj_logic1[279] ,
    \mprj_logic1[278] ,
    \mprj_logic1[277] ,
    \mprj_logic1[276] ,
    \mprj_logic1[275] ,
    \mprj_logic1[274] ,
    \mprj_logic1[273] ,
    \mprj_logic1[272] ,
    \mprj_logic1[271] ,
    \mprj_logic1[270] ,
    \mprj_logic1[269] ,
    \mprj_logic1[268] ,
    \mprj_logic1[267] ,
    \mprj_logic1[266] ,
    \mprj_logic1[265] ,
    \mprj_logic1[264] ,
    \mprj_logic1[263] ,
    \mprj_logic1[262] ,
    \mprj_logic1[261] ,
    \mprj_logic1[260] ,
    \mprj_logic1[259] ,
    \mprj_logic1[258] ,
    \mprj_logic1[257] ,
    \mprj_logic1[256] ,
    \mprj_logic1[255] ,
    \mprj_logic1[254] ,
    \mprj_logic1[253] ,
    \mprj_logic1[252] ,
    \mprj_logic1[251] ,
    \mprj_logic1[250] ,
    \mprj_logic1[249] ,
    \mprj_logic1[248] ,
    \mprj_logic1[247] ,
    \mprj_logic1[246] ,
    \mprj_logic1[245] ,
    \mprj_logic1[244] ,
    \mprj_logic1[243] ,
    \mprj_logic1[242] ,
    \mprj_logic1[241] ,
    \mprj_logic1[240] ,
    \mprj_logic1[239] ,
    \mprj_logic1[238] ,
    \mprj_logic1[237] ,
    \mprj_logic1[236] ,
    \mprj_logic1[235] ,
    \mprj_logic1[234] ,
    \mprj_logic1[233] ,
    \mprj_logic1[232] ,
    \mprj_logic1[231] ,
    \mprj_logic1[230] ,
    \mprj_logic1[229] ,
    \mprj_logic1[228] ,
    \mprj_logic1[227] ,
    \mprj_logic1[226] ,
    \mprj_logic1[225] ,
    \mprj_logic1[224] ,
    \mprj_logic1[223] ,
    \mprj_logic1[222] ,
    \mprj_logic1[221] ,
    \mprj_logic1[220] ,
    \mprj_logic1[219] ,
    \mprj_logic1[218] ,
    \mprj_logic1[217] ,
    \mprj_logic1[216] ,
    \mprj_logic1[215] ,
    \mprj_logic1[214] ,
    \mprj_logic1[213] ,
    \mprj_logic1[212] ,
    \mprj_logic1[211] ,
    \mprj_logic1[210] ,
    \mprj_logic1[209] ,
    \mprj_logic1[208] ,
    \mprj_logic1[207] ,
    \mprj_logic1[206] ,
    \mprj_logic1[205] ,
    \mprj_logic1[204] ,
    \mprj_logic1[203] ,
    \mprj_logic1[202] ,
    \mprj_logic1[201] ,
    \mprj_logic1[200] ,
    \mprj_logic1[199] ,
    \mprj_logic1[198] ,
    \mprj_logic1[197] ,
    \mprj_logic1[196] ,
    \mprj_logic1[195] ,
    \mprj_logic1[194] ,
    \mprj_logic1[193] ,
    \mprj_logic1[192] ,
    \mprj_logic1[191] ,
    \mprj_logic1[190] ,
    \mprj_logic1[189] ,
    \mprj_logic1[188] ,
    \mprj_logic1[187] ,
    \mprj_logic1[186] ,
    \mprj_logic1[185] ,
    \mprj_logic1[184] ,
    \mprj_logic1[183] ,
    \mprj_logic1[182] ,
    \mprj_logic1[181] ,
    \mprj_logic1[180] ,
    \mprj_logic1[179] ,
    \mprj_logic1[178] ,
    \mprj_logic1[177] ,
    \mprj_logic1[176] ,
    \mprj_logic1[175] ,
    \mprj_logic1[174] ,
    \mprj_logic1[173] ,
    \mprj_logic1[172] ,
    \mprj_logic1[171] ,
    \mprj_logic1[170] ,
    \mprj_logic1[169] ,
    \mprj_logic1[168] ,
    \mprj_logic1[167] ,
    \mprj_logic1[166] ,
    \mprj_logic1[165] ,
    \mprj_logic1[164] ,
    \mprj_logic1[163] ,
    \mprj_logic1[162] ,
    \mprj_logic1[161] ,
    \mprj_logic1[160] ,
    \mprj_logic1[159] ,
    \mprj_logic1[158] ,
    \mprj_logic1[157] ,
    \mprj_logic1[156] ,
    \mprj_logic1[155] ,
    \mprj_logic1[154] ,
    \mprj_logic1[153] ,
    \mprj_logic1[152] ,
    \mprj_logic1[151] ,
    \mprj_logic1[150] ,
    \mprj_logic1[149] ,
    \mprj_logic1[148] ,
    \mprj_logic1[147] ,
    \mprj_logic1[146] ,
    \mprj_logic1[145] ,
    \mprj_logic1[144] ,
    \mprj_logic1[143] ,
    \mprj_logic1[142] ,
    \mprj_logic1[141] ,
    \mprj_logic1[140] ,
    \mprj_logic1[139] ,
    \mprj_logic1[138] ,
    \mprj_logic1[137] ,
    \mprj_logic1[136] ,
    \mprj_logic1[135] ,
    \mprj_logic1[134] ,
    \mprj_logic1[133] ,
    \mprj_logic1[132] ,
    \mprj_logic1[131] ,
    \mprj_logic1[130] ,
    \mprj_logic1[129] ,
    \mprj_logic1[128] ,
    \mprj_logic1[127] ,
    \mprj_logic1[126] ,
    \mprj_logic1[125] ,
    \mprj_logic1[124] ,
    \mprj_logic1[123] ,
    \mprj_logic1[122] ,
    \mprj_logic1[121] ,
    \mprj_logic1[120] ,
    \mprj_logic1[119] ,
    \mprj_logic1[118] ,
    \mprj_logic1[117] ,
    \mprj_logic1[116] ,
    \mprj_logic1[115] ,
    \mprj_logic1[114] ,
    \mprj_logic1[113] ,
    \mprj_logic1[112] ,
    \mprj_logic1[111] ,
    \mprj_logic1[110] ,
    \mprj_logic1[109] ,
    \mprj_logic1[108] ,
    \mprj_logic1[107] ,
    \mprj_logic1[106] ,
    \mprj_logic1[105] ,
    \mprj_logic1[104] ,
    \mprj_logic1[103] ,
    \mprj_logic1[102] ,
    \mprj_logic1[101] ,
    \mprj_logic1[100] ,
    \mprj_logic1[99] ,
    \mprj_logic1[98] ,
    \mprj_logic1[97] ,
    \mprj_logic1[96] ,
    \mprj_logic1[95] ,
    \mprj_logic1[94] ,
    \mprj_logic1[93] ,
    \mprj_logic1[92] ,
    \mprj_logic1[91] ,
    \mprj_logic1[90] ,
    \mprj_logic1[89] ,
    \mprj_logic1[88] ,
    \mprj_logic1[87] ,
    \mprj_logic1[86] ,
    \mprj_logic1[85] ,
    \mprj_logic1[84] ,
    \mprj_logic1[83] ,
    \mprj_logic1[82] ,
    \mprj_logic1[81] ,
    \mprj_logic1[80] ,
    \mprj_logic1[79] ,
    \mprj_logic1[78] ,
    \mprj_logic1[77] ,
    \mprj_logic1[76] ,
    \mprj_logic1[75] ,
    \mprj_logic1[74] ,
    \mprj_logic1[73] ,
    \mprj_logic1[72] ,
    \mprj_logic1[71] ,
    \mprj_logic1[70] ,
    \mprj_logic1[69] ,
    \mprj_logic1[68] ,
    \mprj_logic1[67] ,
    \mprj_logic1[66] ,
    \mprj_logic1[65] ,
    \mprj_logic1[64] ,
    \mprj_logic1[63] ,
    \mprj_logic1[62] ,
    \mprj_logic1[61] ,
    \mprj_logic1[60] ,
    \mprj_logic1[59] ,
    \mprj_logic1[58] ,
    \mprj_logic1[57] ,
    \mprj_logic1[56] ,
    \mprj_logic1[55] ,
    \mprj_logic1[54] ,
    \mprj_logic1[53] ,
    \mprj_logic1[52] ,
    \mprj_logic1[51] ,
    \mprj_logic1[50] ,
    \mprj_logic1[49] ,
    \mprj_logic1[48] ,
    \mprj_logic1[47] ,
    \mprj_logic1[46] ,
    \mprj_logic1[45] ,
    \mprj_logic1[44] ,
    \mprj_logic1[43] ,
    \mprj_logic1[42] ,
    \mprj_logic1[41] ,
    \mprj_logic1[40] ,
    \mprj_logic1[39] ,
    \mprj_logic1[38] ,
    \mprj_logic1[37] ,
    \mprj_logic1[36] ,
    \mprj_logic1[35] ,
    \mprj_logic1[34] ,
    \mprj_logic1[33] ,
    \mprj_logic1[32] ,
    \mprj_logic1[31] ,
    \mprj_logic1[30] ,
    \mprj_logic1[29] ,
    \mprj_logic1[28] ,
    \mprj_logic1[27] ,
    \mprj_logic1[26] ,
    \mprj_logic1[25] ,
    \mprj_logic1[24] ,
    \mprj_logic1[23] ,
    \mprj_logic1[22] ,
    \mprj_logic1[21] ,
    \mprj_logic1[20] ,
    \mprj_logic1[19] ,
    \mprj_logic1[18] ,
    \mprj_logic1[17] ,
    \mprj_logic1[16] ,
    \mprj_logic1[15] ,
    \mprj_logic1[14] ,
    \mprj_logic1[13] ,
    \mprj_logic1[12] ,
    \mprj_logic1[11] ,
    \mprj_logic1[10] ,
    \mprj_logic1[9] ,
    \mprj_logic1[8] ,
    \mprj_logic1[7] ,
    \mprj_logic1[6] ,
    \mprj_logic1[5] ,
    \mprj_logic1[4] ,
    \mprj_logic1[3] ,
    \mprj_logic1[2] ,
    \mprj_logic1[1] ,
    \mprj_logic1[0] }));
 mgmt_protect_hv powergood_check (.mprj2_vdd_logic1(net954),
    .mprj_vdd_logic1(net952));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[0]  (.A(user_irq_core[0]),
    .B(\user_irq_enable[0] ),
    .Y(\user_irq_bar[0] ));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[1]  (.A(user_irq_core[1]),
    .B(\user_irq_enable[1] ),
    .Y(\user_irq_bar[1] ));
 sky130_fd_sc_hd__nand2_1 \user_irq_gates[2]  (.A(user_irq_core[2]),
    .B(\user_irq_enable[2] ),
    .Y(\user_irq_bar[2] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[0]  (.A(la_data_out_core[0]),
    .B(\la_data_in_enable[0] ),
    .Y(\la_data_in_mprj_bar[0] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[100]  (.A(la_data_out_core[100]),
    .B(\la_data_in_enable[100] ),
    .Y(\la_data_in_mprj_bar[100] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[101]  (.A(la_data_out_core[101]),
    .B(\la_data_in_enable[101] ),
    .Y(\la_data_in_mprj_bar[101] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[102]  (.A(la_data_out_core[102]),
    .B(\la_data_in_enable[102] ),
    .Y(\la_data_in_mprj_bar[102] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[103]  (.A(la_data_out_core[103]),
    .B(\la_data_in_enable[103] ),
    .Y(\la_data_in_mprj_bar[103] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[104]  (.A(la_data_out_core[104]),
    .B(\la_data_in_enable[104] ),
    .Y(\la_data_in_mprj_bar[104] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[105]  (.A(la_data_out_core[105]),
    .B(net1328),
    .Y(\la_data_in_mprj_bar[105] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[106]  (.A(la_data_out_core[106]),
    .B(\la_data_in_enable[106] ),
    .Y(\la_data_in_mprj_bar[106] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[107]  (.A(la_data_out_core[107]),
    .B(\la_data_in_enable[107] ),
    .Y(\la_data_in_mprj_bar[107] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[108]  (.A(la_data_out_core[108]),
    .B(\la_data_in_enable[108] ),
    .Y(\la_data_in_mprj_bar[108] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[109]  (.A(la_data_out_core[109]),
    .B(\la_data_in_enable[109] ),
    .Y(\la_data_in_mprj_bar[109] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[10]  (.A(la_data_out_core[10]),
    .B(\la_data_in_enable[10] ),
    .Y(\la_data_in_mprj_bar[10] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[110]  (.A(la_data_out_core[110]),
    .B(\la_data_in_enable[110] ),
    .Y(\la_data_in_mprj_bar[110] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[111]  (.A(la_data_out_core[111]),
    .B(\la_data_in_enable[111] ),
    .Y(\la_data_in_mprj_bar[111] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[112]  (.A(la_data_out_core[112]),
    .B(\la_data_in_enable[112] ),
    .Y(\la_data_in_mprj_bar[112] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[113]  (.A(la_data_out_core[113]),
    .B(\la_data_in_enable[113] ),
    .Y(\la_data_in_mprj_bar[113] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[114]  (.A(la_data_out_core[114]),
    .B(\la_data_in_enable[114] ),
    .Y(\la_data_in_mprj_bar[114] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[115]  (.A(la_data_out_core[115]),
    .B(\la_data_in_enable[115] ),
    .Y(\la_data_in_mprj_bar[115] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[116]  (.A(la_data_out_core[116]),
    .B(\la_data_in_enable[116] ),
    .Y(\la_data_in_mprj_bar[116] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[117]  (.A(la_data_out_core[117]),
    .B(\la_data_in_enable[117] ),
    .Y(\la_data_in_mprj_bar[117] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[118]  (.A(la_data_out_core[118]),
    .B(\la_data_in_enable[118] ),
    .Y(\la_data_in_mprj_bar[118] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[119]  (.A(la_data_out_core[119]),
    .B(\la_data_in_enable[119] ),
    .Y(\la_data_in_mprj_bar[119] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[11]  (.A(la_data_out_core[11]),
    .B(\la_data_in_enable[11] ),
    .Y(\la_data_in_mprj_bar[11] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[120]  (.A(la_data_out_core[120]),
    .B(\la_data_in_enable[120] ),
    .Y(\la_data_in_mprj_bar[120] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[121]  (.A(la_data_out_core[121]),
    .B(\la_data_in_enable[121] ),
    .Y(\la_data_in_mprj_bar[121] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[122]  (.A(la_data_out_core[122]),
    .B(\la_data_in_enable[122] ),
    .Y(\la_data_in_mprj_bar[122] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[123]  (.A(la_data_out_core[123]),
    .B(\la_data_in_enable[123] ),
    .Y(\la_data_in_mprj_bar[123] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[124]  (.A(la_data_out_core[124]),
    .B(\la_data_in_enable[124] ),
    .Y(\la_data_in_mprj_bar[124] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[125]  (.A(la_data_out_core[125]),
    .B(\la_data_in_enable[125] ),
    .Y(\la_data_in_mprj_bar[125] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[126]  (.A(la_data_out_core[126]),
    .B(\la_data_in_enable[126] ),
    .Y(\la_data_in_mprj_bar[126] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[127]  (.A(la_data_out_core[127]),
    .B(\la_data_in_enable[127] ),
    .Y(\la_data_in_mprj_bar[127] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[12]  (.A(la_data_out_core[12]),
    .B(\la_data_in_enable[12] ),
    .Y(\la_data_in_mprj_bar[12] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[13]  (.A(la_data_out_core[13]),
    .B(\la_data_in_enable[13] ),
    .Y(\la_data_in_mprj_bar[13] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[14]  (.A(la_data_out_core[14]),
    .B(\la_data_in_enable[14] ),
    .Y(\la_data_in_mprj_bar[14] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[15]  (.A(la_data_out_core[15]),
    .B(\la_data_in_enable[15] ),
    .Y(\la_data_in_mprj_bar[15] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[16]  (.A(la_data_out_core[16]),
    .B(\la_data_in_enable[16] ),
    .Y(\la_data_in_mprj_bar[16] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[17]  (.A(la_data_out_core[17]),
    .B(\la_data_in_enable[17] ),
    .Y(\la_data_in_mprj_bar[17] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[18]  (.A(la_data_out_core[18]),
    .B(\la_data_in_enable[18] ),
    .Y(\la_data_in_mprj_bar[18] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[19]  (.A(la_data_out_core[19]),
    .B(\la_data_in_enable[19] ),
    .Y(\la_data_in_mprj_bar[19] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[1]  (.A(la_data_out_core[1]),
    .B(\la_data_in_enable[1] ),
    .Y(\la_data_in_mprj_bar[1] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[20]  (.A(la_data_out_core[20]),
    .B(\la_data_in_enable[20] ),
    .Y(\la_data_in_mprj_bar[20] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[21]  (.A(la_data_out_core[21]),
    .B(\la_data_in_enable[21] ),
    .Y(\la_data_in_mprj_bar[21] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[22]  (.A(la_data_out_core[22]),
    .B(\la_data_in_enable[22] ),
    .Y(\la_data_in_mprj_bar[22] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[23]  (.A(la_data_out_core[23]),
    .B(\la_data_in_enable[23] ),
    .Y(\la_data_in_mprj_bar[23] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[24]  (.A(la_data_out_core[24]),
    .B(\la_data_in_enable[24] ),
    .Y(\la_data_in_mprj_bar[24] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[25]  (.A(la_data_out_core[25]),
    .B(\la_data_in_enable[25] ),
    .Y(\la_data_in_mprj_bar[25] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[26]  (.A(la_data_out_core[26]),
    .B(\la_data_in_enable[26] ),
    .Y(\la_data_in_mprj_bar[26] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[27]  (.A(la_data_out_core[27]),
    .B(\la_data_in_enable[27] ),
    .Y(\la_data_in_mprj_bar[27] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[28]  (.A(la_data_out_core[28]),
    .B(\la_data_in_enable[28] ),
    .Y(\la_data_in_mprj_bar[28] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[29]  (.A(la_data_out_core[29]),
    .B(\la_data_in_enable[29] ),
    .Y(\la_data_in_mprj_bar[29] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[2]  (.A(la_data_out_core[2]),
    .B(\la_data_in_enable[2] ),
    .Y(\la_data_in_mprj_bar[2] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[30]  (.A(la_data_out_core[30]),
    .B(\la_data_in_enable[30] ),
    .Y(\la_data_in_mprj_bar[30] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[31]  (.A(la_data_out_core[31]),
    .B(\la_data_in_enable[31] ),
    .Y(\la_data_in_mprj_bar[31] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[32]  (.A(la_data_out_core[32]),
    .B(\la_data_in_enable[32] ),
    .Y(\la_data_in_mprj_bar[32] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[33]  (.A(la_data_out_core[33]),
    .B(\la_data_in_enable[33] ),
    .Y(\la_data_in_mprj_bar[33] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[34]  (.A(la_data_out_core[34]),
    .B(\la_data_in_enable[34] ),
    .Y(\la_data_in_mprj_bar[34] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[35]  (.A(la_data_out_core[35]),
    .B(\la_data_in_enable[35] ),
    .Y(\la_data_in_mprj_bar[35] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[36]  (.A(la_data_out_core[36]),
    .B(\la_data_in_enable[36] ),
    .Y(\la_data_in_mprj_bar[36] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[37]  (.A(la_data_out_core[37]),
    .B(\la_data_in_enable[37] ),
    .Y(\la_data_in_mprj_bar[37] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[38]  (.A(la_data_out_core[38]),
    .B(\la_data_in_enable[38] ),
    .Y(\la_data_in_mprj_bar[38] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[39]  (.A(la_data_out_core[39]),
    .B(\la_data_in_enable[39] ),
    .Y(\la_data_in_mprj_bar[39] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[3]  (.A(la_data_out_core[3]),
    .B(\la_data_in_enable[3] ),
    .Y(\la_data_in_mprj_bar[3] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[40]  (.A(la_data_out_core[40]),
    .B(\la_data_in_enable[40] ),
    .Y(\la_data_in_mprj_bar[40] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[41]  (.A(la_data_out_core[41]),
    .B(\la_data_in_enable[41] ),
    .Y(\la_data_in_mprj_bar[41] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[42]  (.A(la_data_out_core[42]),
    .B(\la_data_in_enable[42] ),
    .Y(\la_data_in_mprj_bar[42] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[43]  (.A(la_data_out_core[43]),
    .B(\la_data_in_enable[43] ),
    .Y(\la_data_in_mprj_bar[43] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[44]  (.A(la_data_out_core[44]),
    .B(\la_data_in_enable[44] ),
    .Y(\la_data_in_mprj_bar[44] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[45]  (.A(la_data_out_core[45]),
    .B(\la_data_in_enable[45] ),
    .Y(\la_data_in_mprj_bar[45] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[46]  (.A(la_data_out_core[46]),
    .B(\la_data_in_enable[46] ),
    .Y(\la_data_in_mprj_bar[46] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[47]  (.A(la_data_out_core[47]),
    .B(\la_data_in_enable[47] ),
    .Y(\la_data_in_mprj_bar[47] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[48]  (.A(la_data_out_core[48]),
    .B(\la_data_in_enable[48] ),
    .Y(\la_data_in_mprj_bar[48] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[49]  (.A(la_data_out_core[49]),
    .B(\la_data_in_enable[49] ),
    .Y(\la_data_in_mprj_bar[49] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[4]  (.A(la_data_out_core[4]),
    .B(\la_data_in_enable[4] ),
    .Y(\la_data_in_mprj_bar[4] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[50]  (.A(la_data_out_core[50]),
    .B(\la_data_in_enable[50] ),
    .Y(\la_data_in_mprj_bar[50] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[51]  (.A(la_data_out_core[51]),
    .B(\la_data_in_enable[51] ),
    .Y(\la_data_in_mprj_bar[51] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[52]  (.A(la_data_out_core[52]),
    .B(\la_data_in_enable[52] ),
    .Y(\la_data_in_mprj_bar[52] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[53]  (.A(la_data_out_core[53]),
    .B(\la_data_in_enable[53] ),
    .Y(\la_data_in_mprj_bar[53] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[54]  (.A(la_data_out_core[54]),
    .B(\la_data_in_enable[54] ),
    .Y(\la_data_in_mprj_bar[54] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[55]  (.A(la_data_out_core[55]),
    .B(\la_data_in_enable[55] ),
    .Y(\la_data_in_mprj_bar[55] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[56]  (.A(la_data_out_core[56]),
    .B(\la_data_in_enable[56] ),
    .Y(\la_data_in_mprj_bar[56] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[57]  (.A(la_data_out_core[57]),
    .B(\la_data_in_enable[57] ),
    .Y(\la_data_in_mprj_bar[57] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[58]  (.A(la_data_out_core[58]),
    .B(\la_data_in_enable[58] ),
    .Y(\la_data_in_mprj_bar[58] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[59]  (.A(la_data_out_core[59]),
    .B(\la_data_in_enable[59] ),
    .Y(\la_data_in_mprj_bar[59] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[5]  (.A(la_data_out_core[5]),
    .B(\la_data_in_enable[5] ),
    .Y(\la_data_in_mprj_bar[5] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[60]  (.A(la_data_out_core[60]),
    .B(\la_data_in_enable[60] ),
    .Y(\la_data_in_mprj_bar[60] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[61]  (.A(la_data_out_core[61]),
    .B(\la_data_in_enable[61] ),
    .Y(\la_data_in_mprj_bar[61] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[62]  (.A(la_data_out_core[62]),
    .B(\la_data_in_enable[62] ),
    .Y(\la_data_in_mprj_bar[62] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[63]  (.A(la_data_out_core[63]),
    .B(\la_data_in_enable[63] ),
    .Y(\la_data_in_mprj_bar[63] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[64]  (.A(la_data_out_core[64]),
    .B(\la_data_in_enable[64] ),
    .Y(\la_data_in_mprj_bar[64] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[65]  (.A(la_data_out_core[65]),
    .B(\la_data_in_enable[65] ),
    .Y(\la_data_in_mprj_bar[65] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[66]  (.A(la_data_out_core[66]),
    .B(\la_data_in_enable[66] ),
    .Y(\la_data_in_mprj_bar[66] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[67]  (.A(la_data_out_core[67]),
    .B(\la_data_in_enable[67] ),
    .Y(\la_data_in_mprj_bar[67] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[68]  (.A(la_data_out_core[68]),
    .B(\la_data_in_enable[68] ),
    .Y(\la_data_in_mprj_bar[68] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[69]  (.A(la_data_out_core[69]),
    .B(\la_data_in_enable[69] ),
    .Y(\la_data_in_mprj_bar[69] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[6]  (.A(la_data_out_core[6]),
    .B(\la_data_in_enable[6] ),
    .Y(\la_data_in_mprj_bar[6] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[70]  (.A(la_data_out_core[70]),
    .B(\la_data_in_enable[70] ),
    .Y(\la_data_in_mprj_bar[70] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[71]  (.A(la_data_out_core[71]),
    .B(\la_data_in_enable[71] ),
    .Y(\la_data_in_mprj_bar[71] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[72]  (.A(la_data_out_core[72]),
    .B(\la_data_in_enable[72] ),
    .Y(\la_data_in_mprj_bar[72] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[73]  (.A(la_data_out_core[73]),
    .B(\la_data_in_enable[73] ),
    .Y(\la_data_in_mprj_bar[73] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[74]  (.A(la_data_out_core[74]),
    .B(\la_data_in_enable[74] ),
    .Y(\la_data_in_mprj_bar[74] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[75]  (.A(la_data_out_core[75]),
    .B(\la_data_in_enable[75] ),
    .Y(\la_data_in_mprj_bar[75] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[76]  (.A(la_data_out_core[76]),
    .B(\la_data_in_enable[76] ),
    .Y(\la_data_in_mprj_bar[76] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[77]  (.A(la_data_out_core[77]),
    .B(\la_data_in_enable[77] ),
    .Y(\la_data_in_mprj_bar[77] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[78]  (.A(la_data_out_core[78]),
    .B(\la_data_in_enable[78] ),
    .Y(\la_data_in_mprj_bar[78] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[79]  (.A(la_data_out_core[79]),
    .B(\la_data_in_enable[79] ),
    .Y(\la_data_in_mprj_bar[79] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[7]  (.A(la_data_out_core[7]),
    .B(\la_data_in_enable[7] ),
    .Y(\la_data_in_mprj_bar[7] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[80]  (.A(la_data_out_core[80]),
    .B(\la_data_in_enable[80] ),
    .Y(\la_data_in_mprj_bar[80] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[81]  (.A(la_data_out_core[81]),
    .B(\la_data_in_enable[81] ),
    .Y(\la_data_in_mprj_bar[81] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[82]  (.A(la_data_out_core[82]),
    .B(\la_data_in_enable[82] ),
    .Y(\la_data_in_mprj_bar[82] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[83]  (.A(la_data_out_core[83]),
    .B(\la_data_in_enable[83] ),
    .Y(\la_data_in_mprj_bar[83] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[84]  (.A(la_data_out_core[84]),
    .B(\la_data_in_enable[84] ),
    .Y(\la_data_in_mprj_bar[84] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[85]  (.A(la_data_out_core[85]),
    .B(\la_data_in_enable[85] ),
    .Y(\la_data_in_mprj_bar[85] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[86]  (.A(la_data_out_core[86]),
    .B(\la_data_in_enable[86] ),
    .Y(\la_data_in_mprj_bar[86] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[87]  (.A(la_data_out_core[87]),
    .B(\la_data_in_enable[87] ),
    .Y(\la_data_in_mprj_bar[87] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[88]  (.A(la_data_out_core[88]),
    .B(\la_data_in_enable[88] ),
    .Y(\la_data_in_mprj_bar[88] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[89]  (.A(la_data_out_core[89]),
    .B(\la_data_in_enable[89] ),
    .Y(\la_data_in_mprj_bar[89] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[8]  (.A(la_data_out_core[8]),
    .B(\la_data_in_enable[8] ),
    .Y(\la_data_in_mprj_bar[8] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[90]  (.A(la_data_out_core[90]),
    .B(\la_data_in_enable[90] ),
    .Y(\la_data_in_mprj_bar[90] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[91]  (.A(la_data_out_core[91]),
    .B(\la_data_in_enable[91] ),
    .Y(\la_data_in_mprj_bar[91] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[92]  (.A(la_data_out_core[92]),
    .B(\la_data_in_enable[92] ),
    .Y(\la_data_in_mprj_bar[92] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[93]  (.A(la_data_out_core[93]),
    .B(\la_data_in_enable[93] ),
    .Y(\la_data_in_mprj_bar[93] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[94]  (.A(la_data_out_core[94]),
    .B(\la_data_in_enable[94] ),
    .Y(\la_data_in_mprj_bar[94] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[95]  (.A(la_data_out_core[95]),
    .B(\la_data_in_enable[95] ),
    .Y(\la_data_in_mprj_bar[95] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[96]  (.A(la_data_out_core[96]),
    .B(\la_data_in_enable[96] ),
    .Y(\la_data_in_mprj_bar[96] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[97]  (.A(la_data_out_core[97]),
    .B(\la_data_in_enable[97] ),
    .Y(\la_data_in_mprj_bar[97] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[98]  (.A(la_data_out_core[98]),
    .B(\la_data_in_enable[98] ),
    .Y(\la_data_in_mprj_bar[98] ));
 sky130_fd_sc_hd__nand2_2 \user_to_mprj_in_gates[99]  (.A(la_data_out_core[99]),
    .B(\la_data_in_enable[99] ),
    .Y(\la_data_in_mprj_bar[99] ));
 sky130_fd_sc_hd__nand2_1 \user_to_mprj_in_gates[9]  (.A(la_data_out_core[9]),
    .B(\la_data_in_enable[9] ),
    .Y(\la_data_in_mprj_bar[9] ));
 sky130_fd_sc_hd__nand2_1 user_wb_ack_gate (.A(mprj_ack_i_user),
    .B(net1326),
    .Y(mprj_ack_i_core_bar));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[0]  (.A(mprj_dat_i_user[0]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[0] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[10]  (.A(mprj_dat_i_user[10]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[10] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[11]  (.A(mprj_dat_i_user[11]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[11] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[12]  (.A(mprj_dat_i_user[12]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[12] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[13]  (.A(mprj_dat_i_user[13]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[13] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[14]  (.A(mprj_dat_i_user[14]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[14] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[15]  (.A(mprj_dat_i_user[15]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[15] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[16]  (.A(mprj_dat_i_user[16]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[16] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[17]  (.A(mprj_dat_i_user[17]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[17] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[18]  (.A(mprj_dat_i_user[18]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[18] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[19]  (.A(mprj_dat_i_user[19]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[19] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[1]  (.A(mprj_dat_i_user[1]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[1] ));
 sky130_fd_sc_hd__nand2_2 \user_wb_dat_gates[20]  (.A(mprj_dat_i_user[20]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[20] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[21]  (.A(mprj_dat_i_user[21]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[21] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[22]  (.A(mprj_dat_i_user[22]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[22] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[23]  (.A(mprj_dat_i_user[23]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[23] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[24]  (.A(mprj_dat_i_user[24]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[24] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[25]  (.A(mprj_dat_i_user[25]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[25] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[26]  (.A(mprj_dat_i_user[26]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[26] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[27]  (.A(mprj_dat_i_user[27]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[27] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[28]  (.A(mprj_dat_i_user[28]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[28] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[29]  (.A(mprj_dat_i_user[29]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[29] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[2]  (.A(mprj_dat_i_user[2]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[2] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[30]  (.A(mprj_dat_i_user[30]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[30] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[31]  (.A(mprj_dat_i_user[31]),
    .B(wb_in_enable),
    .Y(\mprj_dat_i_core_bar[31] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[3]  (.A(mprj_dat_i_user[3]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[3] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[4]  (.A(mprj_dat_i_user[4]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[4] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[5]  (.A(mprj_dat_i_user[5]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[5] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[6]  (.A(mprj_dat_i_user[6]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[6] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[7]  (.A(mprj_dat_i_user[7]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[7] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[8]  (.A(mprj_dat_i_user[8]),
    .B(net1326),
    .Y(\mprj_dat_i_core_bar[8] ));
 sky130_fd_sc_hd__nand2_1 \user_wb_dat_gates[9]  (.A(mprj_dat_i_user[9]),
    .B(net1327),
    .Y(\mprj_dat_i_core_bar[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(caravel_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(caravel_clk2),
    .X(net2));
 sky130_fd_sc_hd__buf_6 input3 (.A(caravel_rstn),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(la_data_out_mprj[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(la_data_out_mprj[100]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(la_data_out_mprj[101]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(la_data_out_mprj[102]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(la_data_out_mprj[103]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(la_data_out_mprj[104]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(la_data_out_mprj[105]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(la_data_out_mprj[106]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(la_data_out_mprj[107]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(la_data_out_mprj[108]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(la_data_out_mprj[109]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(la_data_out_mprj[10]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(la_data_out_mprj[110]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(la_data_out_mprj[111]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(la_data_out_mprj[112]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(la_data_out_mprj[113]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(la_data_out_mprj[114]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(la_data_out_mprj[115]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(la_data_out_mprj[116]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(la_data_out_mprj[117]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(la_data_out_mprj[118]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(la_data_out_mprj[119]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(la_data_out_mprj[11]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(la_data_out_mprj[120]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(la_data_out_mprj[121]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(la_data_out_mprj[122]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(la_data_out_mprj[123]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(la_data_out_mprj[124]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(la_data_out_mprj[125]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(la_data_out_mprj[126]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(la_data_out_mprj[127]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(la_data_out_mprj[12]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(la_data_out_mprj[13]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(la_data_out_mprj[14]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(la_data_out_mprj[15]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(la_data_out_mprj[16]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(la_data_out_mprj[17]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(la_data_out_mprj[18]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(la_data_out_mprj[19]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(la_data_out_mprj[1]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(la_data_out_mprj[20]),
    .X(net44));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(la_data_out_mprj[21]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(la_data_out_mprj[22]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(la_data_out_mprj[23]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(la_data_out_mprj[24]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(la_data_out_mprj[25]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input50 (.A(la_data_out_mprj[26]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(la_data_out_mprj[27]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(la_data_out_mprj[28]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(la_data_out_mprj[29]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(la_data_out_mprj[2]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(la_data_out_mprj[30]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(la_data_out_mprj[31]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(la_data_out_mprj[32]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(la_data_out_mprj[33]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(la_data_out_mprj[34]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(la_data_out_mprj[35]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(la_data_out_mprj[36]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(la_data_out_mprj[37]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(la_data_out_mprj[38]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(la_data_out_mprj[39]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(la_data_out_mprj[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(la_data_out_mprj[40]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(la_data_out_mprj[41]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(la_data_out_mprj[42]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(la_data_out_mprj[43]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(la_data_out_mprj[44]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(la_data_out_mprj[45]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(la_data_out_mprj[46]),
    .X(net72));
 sky130_fd_sc_hd__dlymetal6s2s_1 input73 (.A(la_data_out_mprj[47]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(la_data_out_mprj[48]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(la_data_out_mprj[49]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(la_data_out_mprj[4]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(la_data_out_mprj[50]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(la_data_out_mprj[51]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(la_data_out_mprj[52]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(la_data_out_mprj[53]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(la_data_out_mprj[54]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(la_data_out_mprj[55]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(la_data_out_mprj[56]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(la_data_out_mprj[57]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(la_data_out_mprj[58]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(la_data_out_mprj[59]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(la_data_out_mprj[5]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(la_data_out_mprj[60]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(la_data_out_mprj[61]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(la_data_out_mprj[62]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(la_data_out_mprj[63]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(la_data_out_mprj[64]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(la_data_out_mprj[65]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(la_data_out_mprj[66]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 input95 (.A(la_data_out_mprj[67]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 input96 (.A(la_data_out_mprj[68]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(la_data_out_mprj[69]),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 input98 (.A(la_data_out_mprj[6]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 input99 (.A(la_data_out_mprj[70]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(la_data_out_mprj[71]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(la_data_out_mprj[72]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(la_data_out_mprj[73]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_2 input103 (.A(la_data_out_mprj[74]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 input104 (.A(la_data_out_mprj[75]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input105 (.A(la_data_out_mprj[76]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(la_data_out_mprj[77]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(la_data_out_mprj[78]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(la_data_out_mprj[79]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 input109 (.A(la_data_out_mprj[7]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(la_data_out_mprj[80]),
    .X(net110));
 sky130_fd_sc_hd__buf_4 input111 (.A(la_data_out_mprj[81]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(la_data_out_mprj[82]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(la_data_out_mprj[83]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_2 input114 (.A(la_data_out_mprj[84]),
    .X(net114));
 sky130_fd_sc_hd__buf_4 input115 (.A(la_data_out_mprj[85]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(la_data_out_mprj[86]),
    .X(net116));
 sky130_fd_sc_hd__buf_6 input117 (.A(la_data_out_mprj[87]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(la_data_out_mprj[88]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(la_data_out_mprj[89]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(la_data_out_mprj[8]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(la_data_out_mprj[90]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(la_data_out_mprj[91]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(la_data_out_mprj[92]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(la_data_out_mprj[93]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(la_data_out_mprj[94]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(la_data_out_mprj[95]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(la_data_out_mprj[96]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(la_data_out_mprj[97]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(la_data_out_mprj[98]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(la_data_out_mprj[99]),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 input131 (.A(la_data_out_mprj[9]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(la_iena_mprj[0]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(la_iena_mprj[100]),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(la_iena_mprj[101]),
    .X(net134));
 sky130_fd_sc_hd__dlymetal6s2s_1 input135 (.A(la_iena_mprj[102]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(la_iena_mprj[103]),
    .X(net136));
 sky130_fd_sc_hd__dlymetal6s2s_1 input137 (.A(la_iena_mprj[104]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(la_iena_mprj[105]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_2 input139 (.A(la_iena_mprj[106]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(la_iena_mprj[107]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(la_iena_mprj[108]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 input142 (.A(la_iena_mprj[109]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 input143 (.A(la_iena_mprj[10]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(la_iena_mprj[110]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(la_iena_mprj[111]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(la_iena_mprj[112]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(la_iena_mprj[113]),
    .X(net147));
 sky130_fd_sc_hd__dlymetal6s2s_1 input148 (.A(la_iena_mprj[114]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(la_iena_mprj[115]),
    .X(net149));
 sky130_fd_sc_hd__dlymetal6s2s_1 input150 (.A(la_iena_mprj[116]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(la_iena_mprj[117]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(la_iena_mprj[118]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(la_iena_mprj[119]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 input154 (.A(la_iena_mprj[11]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 input155 (.A(la_iena_mprj[120]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 input156 (.A(la_iena_mprj[121]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 input157 (.A(la_iena_mprj[122]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 input158 (.A(la_iena_mprj[123]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 input159 (.A(la_iena_mprj[124]),
    .X(net159));
 sky130_fd_sc_hd__dlymetal6s2s_1 input160 (.A(la_iena_mprj[125]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 input161 (.A(la_iena_mprj[126]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(la_iena_mprj[127]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 input163 (.A(la_iena_mprj[12]),
    .X(net163));
 sky130_fd_sc_hd__dlymetal6s2s_1 input164 (.A(la_iena_mprj[13]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(la_iena_mprj[14]),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 input166 (.A(la_iena_mprj[15]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(la_iena_mprj[16]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 input168 (.A(la_iena_mprj[17]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(la_iena_mprj[18]),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 input170 (.A(la_iena_mprj[19]),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 input171 (.A(la_iena_mprj[1]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(la_iena_mprj[20]),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 input173 (.A(la_iena_mprj[21]),
    .X(net173));
 sky130_fd_sc_hd__dlymetal6s2s_1 input174 (.A(la_iena_mprj[22]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(la_iena_mprj[23]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(la_iena_mprj[24]),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 input177 (.A(la_iena_mprj[25]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(la_iena_mprj[26]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(la_iena_mprj[27]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(la_iena_mprj[28]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(la_iena_mprj[29]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(la_iena_mprj[2]),
    .X(net182));
 sky130_fd_sc_hd__dlymetal6s2s_1 input183 (.A(la_iena_mprj[30]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(la_iena_mprj[31]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(la_iena_mprj[32]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(la_iena_mprj[33]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(la_iena_mprj[34]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(la_iena_mprj[35]),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 input189 (.A(la_iena_mprj[36]),
    .X(net189));
 sky130_fd_sc_hd__dlymetal6s2s_1 input190 (.A(la_iena_mprj[37]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(la_iena_mprj[38]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(la_iena_mprj[39]),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 input193 (.A(la_iena_mprj[3]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(la_iena_mprj[40]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(la_iena_mprj[41]),
    .X(net195));
 sky130_fd_sc_hd__dlymetal6s2s_1 input196 (.A(la_iena_mprj[42]),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(la_iena_mprj[43]),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(la_iena_mprj[44]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(la_iena_mprj[45]),
    .X(net199));
 sky130_fd_sc_hd__dlymetal6s2s_1 input200 (.A(la_iena_mprj[46]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(la_iena_mprj[47]),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(la_iena_mprj[48]),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(la_iena_mprj[49]),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(la_iena_mprj[4]),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(la_iena_mprj[50]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(la_iena_mprj[51]),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 input207 (.A(la_iena_mprj[52]),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(la_iena_mprj[53]),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(la_iena_mprj[54]),
    .X(net209));
 sky130_fd_sc_hd__dlymetal6s2s_1 input210 (.A(la_iena_mprj[55]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 input211 (.A(la_iena_mprj[56]),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 input212 (.A(la_iena_mprj[57]),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_2 input213 (.A(la_iena_mprj[58]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 input214 (.A(la_iena_mprj[59]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(la_iena_mprj[5]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_1 input216 (.A(la_iena_mprj[60]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_1 input217 (.A(la_iena_mprj[61]),
    .X(net217));
 sky130_fd_sc_hd__dlymetal6s2s_1 input218 (.A(la_iena_mprj[62]),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 input219 (.A(la_iena_mprj[63]),
    .X(net219));
 sky130_fd_sc_hd__dlymetal6s2s_1 input220 (.A(la_iena_mprj[64]),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(la_iena_mprj[65]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(la_iena_mprj[66]),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 input223 (.A(la_iena_mprj[67]),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(la_iena_mprj[68]),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(la_iena_mprj[69]),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 input226 (.A(la_iena_mprj[6]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(la_iena_mprj[70]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 input228 (.A(la_iena_mprj[71]),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 input229 (.A(la_iena_mprj[72]),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(la_iena_mprj[73]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(la_iena_mprj[74]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_2 input232 (.A(la_iena_mprj[75]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(la_iena_mprj[76]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 input234 (.A(la_iena_mprj[77]),
    .X(net234));
 sky130_fd_sc_hd__dlymetal6s2s_1 input235 (.A(la_iena_mprj[78]),
    .X(net235));
 sky130_fd_sc_hd__dlymetal6s2s_1 input236 (.A(la_iena_mprj[79]),
    .X(net236));
 sky130_fd_sc_hd__dlymetal6s2s_1 input237 (.A(la_iena_mprj[7]),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input238 (.A(la_iena_mprj[80]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(la_iena_mprj[81]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(la_iena_mprj[82]),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(la_iena_mprj[83]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(la_iena_mprj[84]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(la_iena_mprj[85]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(la_iena_mprj[86]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 input245 (.A(la_iena_mprj[87]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 input246 (.A(la_iena_mprj[88]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 input247 (.A(la_iena_mprj[89]),
    .X(net247));
 sky130_fd_sc_hd__dlymetal6s2s_1 input248 (.A(la_iena_mprj[8]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(la_iena_mprj[90]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(la_iena_mprj[91]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(la_iena_mprj[92]),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(la_iena_mprj[93]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(la_iena_mprj[94]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(la_iena_mprj[95]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 input255 (.A(la_iena_mprj[96]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(la_iena_mprj[97]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 input257 (.A(la_iena_mprj[98]),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(la_iena_mprj[99]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(la_iena_mprj[9]),
    .X(net259));
 sky130_fd_sc_hd__dlymetal6s2s_1 input260 (.A(la_oenb_mprj[0]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 input261 (.A(la_oenb_mprj[100]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 input262 (.A(la_oenb_mprj[101]),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 input263 (.A(la_oenb_mprj[102]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 input264 (.A(la_oenb_mprj[103]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 input265 (.A(la_oenb_mprj[104]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 input266 (.A(la_oenb_mprj[105]),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 input267 (.A(la_oenb_mprj[106]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(la_oenb_mprj[107]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 input269 (.A(la_oenb_mprj[108]),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 input270 (.A(la_oenb_mprj[109]),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 input271 (.A(la_oenb_mprj[10]),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 input272 (.A(la_oenb_mprj[110]),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 input273 (.A(la_oenb_mprj[111]),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 input274 (.A(la_oenb_mprj[112]),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 input275 (.A(la_oenb_mprj[113]),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 input276 (.A(la_oenb_mprj[114]),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 input277 (.A(la_oenb_mprj[115]),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 input278 (.A(la_oenb_mprj[116]),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 input279 (.A(la_oenb_mprj[117]),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 input280 (.A(la_oenb_mprj[118]),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 input281 (.A(la_oenb_mprj[119]),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 input282 (.A(la_oenb_mprj[11]),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 input283 (.A(la_oenb_mprj[120]),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 input284 (.A(la_oenb_mprj[121]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 input285 (.A(la_oenb_mprj[122]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 input286 (.A(la_oenb_mprj[123]),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 input287 (.A(la_oenb_mprj[124]),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_2 input288 (.A(la_oenb_mprj[125]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 input289 (.A(la_oenb_mprj[126]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 input290 (.A(la_oenb_mprj[127]),
    .X(net290));
 sky130_fd_sc_hd__dlymetal6s2s_1 input291 (.A(la_oenb_mprj[12]),
    .X(net291));
 sky130_fd_sc_hd__dlymetal6s2s_1 input292 (.A(la_oenb_mprj[13]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 input293 (.A(la_oenb_mprj[14]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 input294 (.A(la_oenb_mprj[15]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 input295 (.A(la_oenb_mprj[16]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 input296 (.A(la_oenb_mprj[17]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 input297 (.A(la_oenb_mprj[18]),
    .X(net297));
 sky130_fd_sc_hd__dlymetal6s2s_1 input298 (.A(la_oenb_mprj[19]),
    .X(net298));
 sky130_fd_sc_hd__dlymetal6s2s_1 input299 (.A(la_oenb_mprj[1]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 input300 (.A(la_oenb_mprj[20]),
    .X(net300));
 sky130_fd_sc_hd__buf_2 input301 (.A(la_oenb_mprj[21]),
    .X(net301));
 sky130_fd_sc_hd__buf_2 input302 (.A(la_oenb_mprj[22]),
    .X(net302));
 sky130_fd_sc_hd__dlymetal6s2s_1 input303 (.A(la_oenb_mprj[23]),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 input304 (.A(la_oenb_mprj[24]),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 input305 (.A(la_oenb_mprj[25]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(la_oenb_mprj[26]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(la_oenb_mprj[27]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_2 input308 (.A(la_oenb_mprj[28]),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 input309 (.A(la_oenb_mprj[29]),
    .X(net309));
 sky130_fd_sc_hd__buf_2 input310 (.A(la_oenb_mprj[2]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(la_oenb_mprj[30]),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 input312 (.A(la_oenb_mprj[31]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 input313 (.A(la_oenb_mprj[32]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 input314 (.A(la_oenb_mprj[33]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(la_oenb_mprj[34]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(la_oenb_mprj[35]),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 input317 (.A(la_oenb_mprj[36]),
    .X(net317));
 sky130_fd_sc_hd__buf_4 input318 (.A(la_oenb_mprj[37]),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 input319 (.A(la_oenb_mprj[38]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(la_oenb_mprj[39]),
    .X(net320));
 sky130_fd_sc_hd__buf_2 input321 (.A(la_oenb_mprj[3]),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 input322 (.A(la_oenb_mprj[40]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 input323 (.A(la_oenb_mprj[41]),
    .X(net323));
 sky130_fd_sc_hd__buf_2 input324 (.A(la_oenb_mprj[42]),
    .X(net324));
 sky130_fd_sc_hd__buf_6 input325 (.A(la_oenb_mprj[43]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 input326 (.A(la_oenb_mprj[44]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 input327 (.A(la_oenb_mprj[45]),
    .X(net327));
 sky130_fd_sc_hd__buf_2 input328 (.A(la_oenb_mprj[46]),
    .X(net328));
 sky130_fd_sc_hd__buf_6 input329 (.A(la_oenb_mprj[47]),
    .X(net329));
 sky130_fd_sc_hd__buf_6 input330 (.A(la_oenb_mprj[48]),
    .X(net330));
 sky130_fd_sc_hd__buf_2 input331 (.A(la_oenb_mprj[49]),
    .X(net331));
 sky130_fd_sc_hd__dlymetal6s2s_1 input332 (.A(la_oenb_mprj[4]),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 input333 (.A(la_oenb_mprj[50]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 input334 (.A(la_oenb_mprj[51]),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 input335 (.A(la_oenb_mprj[52]),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 input336 (.A(la_oenb_mprj[53]),
    .X(net336));
 sky130_fd_sc_hd__buf_6 input337 (.A(la_oenb_mprj[54]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 input338 (.A(la_oenb_mprj[55]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 input339 (.A(la_oenb_mprj[56]),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 input340 (.A(la_oenb_mprj[57]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 input341 (.A(la_oenb_mprj[58]),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 input342 (.A(la_oenb_mprj[59]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 input343 (.A(la_oenb_mprj[5]),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 input344 (.A(la_oenb_mprj[60]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 input345 (.A(la_oenb_mprj[61]),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 input346 (.A(la_oenb_mprj[62]),
    .X(net346));
 sky130_fd_sc_hd__buf_2 input347 (.A(la_oenb_mprj[63]),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 input348 (.A(la_oenb_mprj[64]),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 input349 (.A(la_oenb_mprj[65]),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 input350 (.A(la_oenb_mprj[66]),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 input351 (.A(la_oenb_mprj[67]),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 input352 (.A(la_oenb_mprj[68]),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 input353 (.A(la_oenb_mprj[69]),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 input354 (.A(la_oenb_mprj[6]),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 input355 (.A(la_oenb_mprj[70]),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 input356 (.A(la_oenb_mprj[71]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_2 input357 (.A(la_oenb_mprj[72]),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 input358 (.A(la_oenb_mprj[73]),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 input359 (.A(la_oenb_mprj[74]),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 input360 (.A(la_oenb_mprj[75]),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 input361 (.A(la_oenb_mprj[76]),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_2 input362 (.A(la_oenb_mprj[77]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 input363 (.A(la_oenb_mprj[78]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 input364 (.A(la_oenb_mprj[79]),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 input365 (.A(la_oenb_mprj[7]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 input366 (.A(la_oenb_mprj[80]),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 input367 (.A(la_oenb_mprj[81]),
    .X(net367));
 sky130_fd_sc_hd__buf_4 input368 (.A(la_oenb_mprj[82]),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_2 input369 (.A(la_oenb_mprj[83]),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 input370 (.A(la_oenb_mprj[84]),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_2 input371 (.A(la_oenb_mprj[85]),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_2 input372 (.A(la_oenb_mprj[86]),
    .X(net372));
 sky130_fd_sc_hd__buf_6 input373 (.A(la_oenb_mprj[87]),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 input374 (.A(la_oenb_mprj[88]),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 input375 (.A(la_oenb_mprj[89]),
    .X(net375));
 sky130_fd_sc_hd__dlymetal6s2s_1 input376 (.A(la_oenb_mprj[8]),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 input377 (.A(la_oenb_mprj[90]),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 input378 (.A(la_oenb_mprj[91]),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 input379 (.A(la_oenb_mprj[92]),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_2 input380 (.A(la_oenb_mprj[93]),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 input381 (.A(la_oenb_mprj[94]),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_2 input382 (.A(la_oenb_mprj[95]),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 input383 (.A(la_oenb_mprj[96]),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 input384 (.A(la_oenb_mprj[97]),
    .X(net384));
 sky130_fd_sc_hd__dlymetal6s2s_1 input385 (.A(la_oenb_mprj[98]),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 input386 (.A(la_oenb_mprj[99]),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 input387 (.A(la_oenb_mprj[9]),
    .X(net387));
 sky130_fd_sc_hd__buf_2 input388 (.A(mprj_adr_o_core[0]),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 input389 (.A(mprj_adr_o_core[10]),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 input390 (.A(mprj_adr_o_core[11]),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 input391 (.A(mprj_adr_o_core[12]),
    .X(net391));
 sky130_fd_sc_hd__buf_6 input392 (.A(mprj_adr_o_core[13]),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 input393 (.A(mprj_adr_o_core[14]),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 input394 (.A(mprj_adr_o_core[15]),
    .X(net394));
 sky130_fd_sc_hd__buf_4 input395 (.A(mprj_adr_o_core[16]),
    .X(net395));
 sky130_fd_sc_hd__buf_6 input396 (.A(mprj_adr_o_core[17]),
    .X(net396));
 sky130_fd_sc_hd__buf_2 input397 (.A(mprj_adr_o_core[18]),
    .X(net397));
 sky130_fd_sc_hd__buf_6 input398 (.A(mprj_adr_o_core[19]),
    .X(net398));
 sky130_fd_sc_hd__buf_6 input399 (.A(mprj_adr_o_core[1]),
    .X(net399));
 sky130_fd_sc_hd__buf_6 input400 (.A(mprj_adr_o_core[20]),
    .X(net400));
 sky130_fd_sc_hd__buf_4 input401 (.A(mprj_adr_o_core[21]),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 input402 (.A(mprj_adr_o_core[22]),
    .X(net402));
 sky130_fd_sc_hd__buf_6 input403 (.A(mprj_adr_o_core[23]),
    .X(net403));
 sky130_fd_sc_hd__buf_6 input404 (.A(mprj_adr_o_core[24]),
    .X(net404));
 sky130_fd_sc_hd__buf_6 input405 (.A(mprj_adr_o_core[25]),
    .X(net405));
 sky130_fd_sc_hd__buf_6 input406 (.A(mprj_adr_o_core[26]),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 input407 (.A(mprj_adr_o_core[27]),
    .X(net407));
 sky130_fd_sc_hd__buf_6 input408 (.A(mprj_adr_o_core[28]),
    .X(net408));
 sky130_fd_sc_hd__buf_6 input409 (.A(mprj_adr_o_core[29]),
    .X(net409));
 sky130_fd_sc_hd__buf_2 input410 (.A(mprj_adr_o_core[2]),
    .X(net410));
 sky130_fd_sc_hd__buf_6 input411 (.A(mprj_adr_o_core[30]),
    .X(net411));
 sky130_fd_sc_hd__buf_6 input412 (.A(mprj_adr_o_core[31]),
    .X(net412));
 sky130_fd_sc_hd__buf_6 input413 (.A(mprj_adr_o_core[3]),
    .X(net413));
 sky130_fd_sc_hd__buf_6 input414 (.A(mprj_adr_o_core[4]),
    .X(net414));
 sky130_fd_sc_hd__buf_6 input415 (.A(mprj_adr_o_core[5]),
    .X(net415));
 sky130_fd_sc_hd__buf_6 input416 (.A(mprj_adr_o_core[6]),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 input417 (.A(mprj_adr_o_core[7]),
    .X(net417));
 sky130_fd_sc_hd__buf_6 input418 (.A(mprj_adr_o_core[8]),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 input419 (.A(mprj_adr_o_core[9]),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 input420 (.A(mprj_cyc_o_core),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_1 input421 (.A(mprj_dat_o_core[0]),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_2 input422 (.A(mprj_dat_o_core[10]),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 input423 (.A(mprj_dat_o_core[11]),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 input424 (.A(mprj_dat_o_core[12]),
    .X(net424));
 sky130_fd_sc_hd__dlymetal6s2s_1 input425 (.A(mprj_dat_o_core[13]),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 input426 (.A(mprj_dat_o_core[14]),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 input427 (.A(mprj_dat_o_core[15]),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 input428 (.A(mprj_dat_o_core[16]),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 input429 (.A(mprj_dat_o_core[17]),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 input430 (.A(mprj_dat_o_core[18]),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 input431 (.A(mprj_dat_o_core[19]),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 input432 (.A(mprj_dat_o_core[1]),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 input433 (.A(mprj_dat_o_core[20]),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 input434 (.A(mprj_dat_o_core[21]),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 input435 (.A(mprj_dat_o_core[22]),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 input436 (.A(mprj_dat_o_core[23]),
    .X(net436));
 sky130_fd_sc_hd__dlymetal6s2s_1 input437 (.A(mprj_dat_o_core[24]),
    .X(net437));
 sky130_fd_sc_hd__dlymetal6s2s_1 input438 (.A(mprj_dat_o_core[25]),
    .X(net438));
 sky130_fd_sc_hd__dlymetal6s2s_1 input439 (.A(mprj_dat_o_core[26]),
    .X(net439));
 sky130_fd_sc_hd__dlymetal6s2s_1 input440 (.A(mprj_dat_o_core[27]),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 input441 (.A(mprj_dat_o_core[28]),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 input442 (.A(mprj_dat_o_core[29]),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 input443 (.A(mprj_dat_o_core[2]),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 input444 (.A(mprj_dat_o_core[30]),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 input445 (.A(mprj_dat_o_core[31]),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 input446 (.A(mprj_dat_o_core[3]),
    .X(net446));
 sky130_fd_sc_hd__buf_4 input447 (.A(mprj_dat_o_core[4]),
    .X(net447));
 sky130_fd_sc_hd__buf_2 input448 (.A(mprj_dat_o_core[5]),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 input449 (.A(mprj_dat_o_core[6]),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 input450 (.A(mprj_dat_o_core[7]),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 input451 (.A(mprj_dat_o_core[8]),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_2 input452 (.A(mprj_dat_o_core[9]),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 input453 (.A(mprj_iena_wb),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 input454 (.A(mprj_sel_o_core[0]),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 input455 (.A(mprj_sel_o_core[1]),
    .X(net455));
 sky130_fd_sc_hd__dlymetal6s2s_1 input456 (.A(mprj_sel_o_core[2]),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_2 input457 (.A(mprj_sel_o_core[3]),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 input458 (.A(mprj_stb_o_core),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 input459 (.A(mprj_we_o_core),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_1 input460 (.A(user_irq_ena[0]),
    .X(net460));
 sky130_fd_sc_hd__dlymetal6s2s_1 input461 (.A(user_irq_ena[1]),
    .X(net461));
 sky130_fd_sc_hd__dlymetal6s2s_1 input462 (.A(user_irq_ena[2]),
    .X(net462));
 sky130_fd_sc_hd__buf_12 output463 (.A(net1148),
    .X(la_data_in_core[0]));
 sky130_fd_sc_hd__buf_12 output464 (.A(net464),
    .X(la_data_in_core[100]));
 sky130_fd_sc_hd__buf_12 output465 (.A(net1101),
    .X(la_data_in_core[101]));
 sky130_fd_sc_hd__buf_12 output466 (.A(net466),
    .X(la_data_in_core[102]));
 sky130_fd_sc_hd__buf_12 output467 (.A(net1100),
    .X(la_data_in_core[103]));
 sky130_fd_sc_hd__buf_12 output468 (.A(net1099),
    .X(la_data_in_core[104]));
 sky130_fd_sc_hd__buf_12 output469 (.A(net1098),
    .X(la_data_in_core[105]));
 sky130_fd_sc_hd__buf_12 output470 (.A(net470),
    .X(la_data_in_core[106]));
 sky130_fd_sc_hd__buf_12 output471 (.A(net1097),
    .X(la_data_in_core[107]));
 sky130_fd_sc_hd__buf_12 output472 (.A(net472),
    .X(la_data_in_core[108]));
 sky130_fd_sc_hd__buf_12 output473 (.A(net1096),
    .X(la_data_in_core[109]));
 sky130_fd_sc_hd__buf_12 output474 (.A(net474),
    .X(la_data_in_core[10]));
 sky130_fd_sc_hd__buf_12 output475 (.A(net475),
    .X(la_data_in_core[110]));
 sky130_fd_sc_hd__buf_12 output476 (.A(net476),
    .X(la_data_in_core[111]));
 sky130_fd_sc_hd__buf_12 output477 (.A(net477),
    .X(la_data_in_core[112]));
 sky130_fd_sc_hd__buf_12 output478 (.A(net478),
    .X(la_data_in_core[113]));
 sky130_fd_sc_hd__buf_12 output479 (.A(net479),
    .X(la_data_in_core[114]));
 sky130_fd_sc_hd__buf_12 output480 (.A(net480),
    .X(la_data_in_core[115]));
 sky130_fd_sc_hd__buf_12 output481 (.A(net481),
    .X(la_data_in_core[116]));
 sky130_fd_sc_hd__buf_12 output482 (.A(net482),
    .X(la_data_in_core[117]));
 sky130_fd_sc_hd__buf_12 output483 (.A(net483),
    .X(la_data_in_core[118]));
 sky130_fd_sc_hd__buf_12 output484 (.A(net484),
    .X(la_data_in_core[119]));
 sky130_fd_sc_hd__buf_12 output485 (.A(net485),
    .X(la_data_in_core[11]));
 sky130_fd_sc_hd__buf_12 output486 (.A(net486),
    .X(la_data_in_core[120]));
 sky130_fd_sc_hd__buf_12 output487 (.A(net487),
    .X(la_data_in_core[121]));
 sky130_fd_sc_hd__buf_12 output488 (.A(net488),
    .X(la_data_in_core[122]));
 sky130_fd_sc_hd__buf_12 output489 (.A(net489),
    .X(la_data_in_core[123]));
 sky130_fd_sc_hd__buf_12 output490 (.A(net490),
    .X(la_data_in_core[124]));
 sky130_fd_sc_hd__buf_12 output491 (.A(net491),
    .X(la_data_in_core[125]));
 sky130_fd_sc_hd__buf_12 output492 (.A(net492),
    .X(la_data_in_core[126]));
 sky130_fd_sc_hd__buf_12 output493 (.A(net493),
    .X(la_data_in_core[127]));
 sky130_fd_sc_hd__buf_12 output494 (.A(net1138),
    .X(la_data_in_core[12]));
 sky130_fd_sc_hd__buf_12 output495 (.A(net1137),
    .X(la_data_in_core[13]));
 sky130_fd_sc_hd__buf_12 output496 (.A(net496),
    .X(la_data_in_core[14]));
 sky130_fd_sc_hd__buf_12 output497 (.A(net497),
    .X(la_data_in_core[15]));
 sky130_fd_sc_hd__buf_12 output498 (.A(net1135),
    .X(la_data_in_core[16]));
 sky130_fd_sc_hd__buf_12 output499 (.A(net499),
    .X(la_data_in_core[17]));
 sky130_fd_sc_hd__buf_12 output500 (.A(net500),
    .X(la_data_in_core[18]));
 sky130_fd_sc_hd__buf_12 output501 (.A(net1133),
    .X(la_data_in_core[19]));
 sky130_fd_sc_hd__buf_12 output502 (.A(net1146),
    .X(la_data_in_core[1]));
 sky130_fd_sc_hd__buf_12 output503 (.A(net1132),
    .X(la_data_in_core[20]));
 sky130_fd_sc_hd__buf_12 output504 (.A(net504),
    .X(la_data_in_core[21]));
 sky130_fd_sc_hd__buf_12 output505 (.A(net505),
    .X(la_data_in_core[22]));
 sky130_fd_sc_hd__buf_12 output506 (.A(net506),
    .X(la_data_in_core[23]));
 sky130_fd_sc_hd__buf_12 output507 (.A(net507),
    .X(la_data_in_core[24]));
 sky130_fd_sc_hd__buf_12 output508 (.A(net508),
    .X(la_data_in_core[25]));
 sky130_fd_sc_hd__buf_12 output509 (.A(net1131),
    .X(la_data_in_core[26]));
 sky130_fd_sc_hd__buf_12 output510 (.A(net1129),
    .X(la_data_in_core[27]));
 sky130_fd_sc_hd__buf_12 output511 (.A(net1128),
    .X(la_data_in_core[28]));
 sky130_fd_sc_hd__buf_12 output512 (.A(net1127),
    .X(la_data_in_core[29]));
 sky130_fd_sc_hd__buf_12 output513 (.A(net1145),
    .X(la_data_in_core[2]));
 sky130_fd_sc_hd__buf_12 output514 (.A(net514),
    .X(la_data_in_core[30]));
 sky130_fd_sc_hd__buf_12 output515 (.A(net1126),
    .X(la_data_in_core[31]));
 sky130_fd_sc_hd__buf_12 output516 (.A(net1124),
    .X(la_data_in_core[32]));
 sky130_fd_sc_hd__buf_12 output517 (.A(net1122),
    .X(la_data_in_core[33]));
 sky130_fd_sc_hd__buf_12 output518 (.A(net1121),
    .X(la_data_in_core[34]));
 sky130_fd_sc_hd__buf_12 output519 (.A(net519),
    .X(la_data_in_core[35]));
 sky130_fd_sc_hd__buf_12 output520 (.A(net520),
    .X(la_data_in_core[36]));
 sky130_fd_sc_hd__buf_12 output521 (.A(net521),
    .X(la_data_in_core[37]));
 sky130_fd_sc_hd__buf_12 output522 (.A(net522),
    .X(la_data_in_core[38]));
 sky130_fd_sc_hd__buf_12 output523 (.A(net523),
    .X(la_data_in_core[39]));
 sky130_fd_sc_hd__buf_12 output524 (.A(net1144),
    .X(la_data_in_core[3]));
 sky130_fd_sc_hd__buf_12 output525 (.A(net1120),
    .X(la_data_in_core[40]));
 sky130_fd_sc_hd__buf_12 output526 (.A(net526),
    .X(la_data_in_core[41]));
 sky130_fd_sc_hd__buf_12 output527 (.A(net527),
    .X(la_data_in_core[42]));
 sky130_fd_sc_hd__buf_12 output528 (.A(net528),
    .X(la_data_in_core[43]));
 sky130_fd_sc_hd__buf_12 output529 (.A(net529),
    .X(la_data_in_core[44]));
 sky130_fd_sc_hd__buf_12 output530 (.A(net530),
    .X(la_data_in_core[45]));
 sky130_fd_sc_hd__buf_12 output531 (.A(net531),
    .X(la_data_in_core[46]));
 sky130_fd_sc_hd__buf_12 output532 (.A(net532),
    .X(la_data_in_core[47]));
 sky130_fd_sc_hd__buf_12 output533 (.A(net1119),
    .X(la_data_in_core[48]));
 sky130_fd_sc_hd__buf_12 output534 (.A(net534),
    .X(la_data_in_core[49]));
 sky130_fd_sc_hd__buf_12 output535 (.A(net1143),
    .X(la_data_in_core[4]));
 sky130_fd_sc_hd__buf_12 output536 (.A(net536),
    .X(la_data_in_core[50]));
 sky130_fd_sc_hd__buf_12 output537 (.A(net537),
    .X(la_data_in_core[51]));
 sky130_fd_sc_hd__buf_12 output538 (.A(net538),
    .X(la_data_in_core[52]));
 sky130_fd_sc_hd__buf_12 output539 (.A(net539),
    .X(la_data_in_core[53]));
 sky130_fd_sc_hd__buf_12 output540 (.A(net540),
    .X(la_data_in_core[54]));
 sky130_fd_sc_hd__buf_12 output541 (.A(net541),
    .X(la_data_in_core[55]));
 sky130_fd_sc_hd__buf_12 output542 (.A(net542),
    .X(la_data_in_core[56]));
 sky130_fd_sc_hd__buf_12 output543 (.A(net543),
    .X(la_data_in_core[57]));
 sky130_fd_sc_hd__buf_12 output544 (.A(net544),
    .X(la_data_in_core[58]));
 sky130_fd_sc_hd__buf_12 output545 (.A(net545),
    .X(la_data_in_core[59]));
 sky130_fd_sc_hd__buf_12 output546 (.A(net1142),
    .X(la_data_in_core[5]));
 sky130_fd_sc_hd__buf_12 output547 (.A(net547),
    .X(la_data_in_core[60]));
 sky130_fd_sc_hd__buf_12 output548 (.A(net548),
    .X(la_data_in_core[61]));
 sky130_fd_sc_hd__buf_12 output549 (.A(net549),
    .X(la_data_in_core[62]));
 sky130_fd_sc_hd__buf_12 output550 (.A(net550),
    .X(la_data_in_core[63]));
 sky130_fd_sc_hd__buf_12 output551 (.A(net551),
    .X(la_data_in_core[64]));
 sky130_fd_sc_hd__buf_12 output552 (.A(net552),
    .X(la_data_in_core[65]));
 sky130_fd_sc_hd__buf_12 output553 (.A(net553),
    .X(la_data_in_core[66]));
 sky130_fd_sc_hd__buf_12 output554 (.A(net554),
    .X(la_data_in_core[67]));
 sky130_fd_sc_hd__buf_12 output555 (.A(net555),
    .X(la_data_in_core[68]));
 sky130_fd_sc_hd__buf_12 output556 (.A(net556),
    .X(la_data_in_core[69]));
 sky130_fd_sc_hd__buf_12 output557 (.A(net1141),
    .X(la_data_in_core[6]));
 sky130_fd_sc_hd__buf_12 output558 (.A(net558),
    .X(la_data_in_core[70]));
 sky130_fd_sc_hd__buf_12 output559 (.A(net559),
    .X(la_data_in_core[71]));
 sky130_fd_sc_hd__buf_12 output560 (.A(net560),
    .X(la_data_in_core[72]));
 sky130_fd_sc_hd__buf_12 output561 (.A(net561),
    .X(la_data_in_core[73]));
 sky130_fd_sc_hd__buf_12 output562 (.A(net562),
    .X(la_data_in_core[74]));
 sky130_fd_sc_hd__buf_12 output563 (.A(net563),
    .X(la_data_in_core[75]));
 sky130_fd_sc_hd__buf_12 output564 (.A(net564),
    .X(la_data_in_core[76]));
 sky130_fd_sc_hd__buf_12 output565 (.A(net565),
    .X(la_data_in_core[77]));
 sky130_fd_sc_hd__buf_12 output566 (.A(net566),
    .X(la_data_in_core[78]));
 sky130_fd_sc_hd__buf_12 output567 (.A(net567),
    .X(la_data_in_core[79]));
 sky130_fd_sc_hd__buf_12 output568 (.A(net1140),
    .X(la_data_in_core[7]));
 sky130_fd_sc_hd__buf_12 output569 (.A(net1118),
    .X(la_data_in_core[80]));
 sky130_fd_sc_hd__buf_12 output570 (.A(net1117),
    .X(la_data_in_core[81]));
 sky130_fd_sc_hd__buf_12 output571 (.A(net1116),
    .X(la_data_in_core[82]));
 sky130_fd_sc_hd__buf_12 output572 (.A(net1115),
    .X(la_data_in_core[83]));
 sky130_fd_sc_hd__buf_12 output573 (.A(net1114),
    .X(la_data_in_core[84]));
 sky130_fd_sc_hd__buf_12 output574 (.A(net574),
    .X(la_data_in_core[85]));
 sky130_fd_sc_hd__buf_12 output575 (.A(net1113),
    .X(la_data_in_core[86]));
 sky130_fd_sc_hd__buf_12 output576 (.A(net1112),
    .X(la_data_in_core[87]));
 sky130_fd_sc_hd__buf_12 output577 (.A(net577),
    .X(la_data_in_core[88]));
 sky130_fd_sc_hd__buf_12 output578 (.A(net1111),
    .X(la_data_in_core[89]));
 sky130_fd_sc_hd__buf_12 output579 (.A(net579),
    .X(la_data_in_core[8]));
 sky130_fd_sc_hd__buf_12 output580 (.A(net580),
    .X(la_data_in_core[90]));
 sky130_fd_sc_hd__buf_12 output581 (.A(net1110),
    .X(la_data_in_core[91]));
 sky130_fd_sc_hd__buf_12 output582 (.A(net1109),
    .X(la_data_in_core[92]));
 sky130_fd_sc_hd__buf_12 output583 (.A(net1108),
    .X(la_data_in_core[93]));
 sky130_fd_sc_hd__buf_12 output584 (.A(net1107),
    .X(la_data_in_core[94]));
 sky130_fd_sc_hd__buf_12 output585 (.A(net1106),
    .X(la_data_in_core[95]));
 sky130_fd_sc_hd__buf_12 output586 (.A(net1105),
    .X(la_data_in_core[96]));
 sky130_fd_sc_hd__buf_12 output587 (.A(net587),
    .X(la_data_in_core[97]));
 sky130_fd_sc_hd__buf_12 output588 (.A(net1103),
    .X(la_data_in_core[98]));
 sky130_fd_sc_hd__buf_12 output589 (.A(net1102),
    .X(la_data_in_core[99]));
 sky130_fd_sc_hd__buf_12 output590 (.A(net1139),
    .X(la_data_in_core[9]));
 sky130_fd_sc_hd__buf_12 output591 (.A(net591),
    .X(la_data_in_mprj[0]));
 sky130_fd_sc_hd__buf_12 output592 (.A(net592),
    .X(la_data_in_mprj[100]));
 sky130_fd_sc_hd__buf_12 output593 (.A(net593),
    .X(la_data_in_mprj[101]));
 sky130_fd_sc_hd__buf_12 output594 (.A(net594),
    .X(la_data_in_mprj[102]));
 sky130_fd_sc_hd__buf_12 output595 (.A(net595),
    .X(la_data_in_mprj[103]));
 sky130_fd_sc_hd__buf_12 output596 (.A(net993),
    .X(la_data_in_mprj[104]));
 sky130_fd_sc_hd__buf_12 output597 (.A(net597),
    .X(la_data_in_mprj[105]));
 sky130_fd_sc_hd__buf_12 output598 (.A(net991),
    .X(la_data_in_mprj[106]));
 sky130_fd_sc_hd__buf_12 output599 (.A(net990),
    .X(la_data_in_mprj[107]));
 sky130_fd_sc_hd__buf_12 output600 (.A(net989),
    .X(la_data_in_mprj[108]));
 sky130_fd_sc_hd__buf_12 output601 (.A(net987),
    .X(la_data_in_mprj[109]));
 sky130_fd_sc_hd__buf_12 output602 (.A(net962),
    .X(la_data_in_mprj[10]));
 sky130_fd_sc_hd__buf_12 output603 (.A(net986),
    .X(la_data_in_mprj[110]));
 sky130_fd_sc_hd__buf_12 output604 (.A(net984),
    .X(la_data_in_mprj[111]));
 sky130_fd_sc_hd__buf_12 output605 (.A(net982),
    .X(la_data_in_mprj[112]));
 sky130_fd_sc_hd__buf_12 output606 (.A(net980),
    .X(la_data_in_mprj[113]));
 sky130_fd_sc_hd__buf_12 output607 (.A(net978),
    .X(la_data_in_mprj[114]));
 sky130_fd_sc_hd__buf_12 output608 (.A(net976),
    .X(la_data_in_mprj[115]));
 sky130_fd_sc_hd__buf_12 output609 (.A(net974),
    .X(la_data_in_mprj[116]));
 sky130_fd_sc_hd__buf_12 output610 (.A(net972),
    .X(la_data_in_mprj[117]));
 sky130_fd_sc_hd__buf_12 output611 (.A(net971),
    .X(la_data_in_mprj[118]));
 sky130_fd_sc_hd__buf_12 output612 (.A(net612),
    .X(la_data_in_mprj[119]));
 sky130_fd_sc_hd__buf_12 output613 (.A(net613),
    .X(la_data_in_mprj[11]));
 sky130_fd_sc_hd__buf_12 output614 (.A(net970),
    .X(la_data_in_mprj[120]));
 sky130_fd_sc_hd__buf_12 output615 (.A(net969),
    .X(la_data_in_mprj[121]));
 sky130_fd_sc_hd__buf_12 output616 (.A(net968),
    .X(la_data_in_mprj[122]));
 sky130_fd_sc_hd__buf_12 output617 (.A(net967),
    .X(la_data_in_mprj[123]));
 sky130_fd_sc_hd__buf_12 output618 (.A(net618),
    .X(la_data_in_mprj[124]));
 sky130_fd_sc_hd__buf_12 output619 (.A(net966),
    .X(la_data_in_mprj[125]));
 sky130_fd_sc_hd__buf_12 output620 (.A(net620),
    .X(la_data_in_mprj[126]));
 sky130_fd_sc_hd__buf_12 output621 (.A(net621),
    .X(la_data_in_mprj[127]));
 sky130_fd_sc_hd__buf_12 output622 (.A(net622),
    .X(la_data_in_mprj[12]));
 sky130_fd_sc_hd__buf_12 output623 (.A(net623),
    .X(la_data_in_mprj[13]));
 sky130_fd_sc_hd__buf_12 output624 (.A(net624),
    .X(la_data_in_mprj[14]));
 sky130_fd_sc_hd__buf_12 output625 (.A(net961),
    .X(la_data_in_mprj[15]));
 sky130_fd_sc_hd__buf_12 output626 (.A(net626),
    .X(la_data_in_mprj[16]));
 sky130_fd_sc_hd__buf_12 output627 (.A(net627),
    .X(la_data_in_mprj[17]));
 sky130_fd_sc_hd__buf_12 output628 (.A(net628),
    .X(la_data_in_mprj[18]));
 sky130_fd_sc_hd__buf_12 output629 (.A(net1012),
    .X(la_data_in_mprj[19]));
 sky130_fd_sc_hd__buf_12 output630 (.A(net630),
    .X(la_data_in_mprj[1]));
 sky130_fd_sc_hd__buf_12 output631 (.A(net1011),
    .X(la_data_in_mprj[20]));
 sky130_fd_sc_hd__buf_12 output632 (.A(net632),
    .X(la_data_in_mprj[21]));
 sky130_fd_sc_hd__buf_12 output633 (.A(net633),
    .X(la_data_in_mprj[22]));
 sky130_fd_sc_hd__buf_12 output634 (.A(net1010),
    .X(la_data_in_mprj[23]));
 sky130_fd_sc_hd__buf_12 output635 (.A(net635),
    .X(la_data_in_mprj[24]));
 sky130_fd_sc_hd__buf_12 output636 (.A(net1009),
    .X(la_data_in_mprj[25]));
 sky130_fd_sc_hd__buf_12 output637 (.A(net1008),
    .X(la_data_in_mprj[26]));
 sky130_fd_sc_hd__buf_12 output638 (.A(net638),
    .X(la_data_in_mprj[27]));
 sky130_fd_sc_hd__buf_12 output639 (.A(net1007),
    .X(la_data_in_mprj[28]));
 sky130_fd_sc_hd__buf_12 output640 (.A(net1006),
    .X(la_data_in_mprj[29]));
 sky130_fd_sc_hd__buf_12 output641 (.A(net641),
    .X(la_data_in_mprj[2]));
 sky130_fd_sc_hd__buf_12 output642 (.A(net1005),
    .X(la_data_in_mprj[30]));
 sky130_fd_sc_hd__buf_12 output643 (.A(net1004),
    .X(la_data_in_mprj[31]));
 sky130_fd_sc_hd__buf_12 output644 (.A(net644),
    .X(la_data_in_mprj[32]));
 sky130_fd_sc_hd__buf_12 output645 (.A(net1003),
    .X(la_data_in_mprj[33]));
 sky130_fd_sc_hd__buf_12 output646 (.A(net1002),
    .X(la_data_in_mprj[34]));
 sky130_fd_sc_hd__buf_12 output647 (.A(net1001),
    .X(la_data_in_mprj[35]));
 sky130_fd_sc_hd__buf_12 output648 (.A(net648),
    .X(la_data_in_mprj[36]));
 sky130_fd_sc_hd__buf_12 output649 (.A(net1000),
    .X(la_data_in_mprj[37]));
 sky130_fd_sc_hd__buf_12 output650 (.A(net999),
    .X(la_data_in_mprj[38]));
 sky130_fd_sc_hd__buf_12 output651 (.A(net651),
    .X(la_data_in_mprj[39]));
 sky130_fd_sc_hd__buf_12 output652 (.A(net652),
    .X(la_data_in_mprj[3]));
 sky130_fd_sc_hd__buf_12 output653 (.A(net653),
    .X(la_data_in_mprj[40]));
 sky130_fd_sc_hd__buf_12 output654 (.A(net654),
    .X(la_data_in_mprj[41]));
 sky130_fd_sc_hd__buf_12 output655 (.A(net998),
    .X(la_data_in_mprj[42]));
 sky130_fd_sc_hd__buf_12 output656 (.A(net656),
    .X(la_data_in_mprj[43]));
 sky130_fd_sc_hd__buf_12 output657 (.A(net657),
    .X(la_data_in_mprj[44]));
 sky130_fd_sc_hd__buf_12 output658 (.A(net997),
    .X(la_data_in_mprj[45]));
 sky130_fd_sc_hd__buf_12 output659 (.A(net659),
    .X(la_data_in_mprj[46]));
 sky130_fd_sc_hd__buf_12 output660 (.A(net996),
    .X(la_data_in_mprj[47]));
 sky130_fd_sc_hd__buf_12 output661 (.A(net661),
    .X(la_data_in_mprj[48]));
 sky130_fd_sc_hd__buf_12 output662 (.A(net662),
    .X(la_data_in_mprj[49]));
 sky130_fd_sc_hd__buf_12 output663 (.A(net663),
    .X(la_data_in_mprj[4]));
 sky130_fd_sc_hd__buf_12 output664 (.A(net664),
    .X(la_data_in_mprj[50]));
 sky130_fd_sc_hd__buf_12 output665 (.A(net995),
    .X(la_data_in_mprj[51]));
 sky130_fd_sc_hd__buf_12 output666 (.A(net994),
    .X(la_data_in_mprj[52]));
 sky130_fd_sc_hd__buf_12 output667 (.A(net667),
    .X(la_data_in_mprj[53]));
 sky130_fd_sc_hd__buf_12 output668 (.A(net668),
    .X(la_data_in_mprj[54]));
 sky130_fd_sc_hd__buf_12 output669 (.A(net669),
    .X(la_data_in_mprj[55]));
 sky130_fd_sc_hd__buf_12 output670 (.A(net670),
    .X(la_data_in_mprj[56]));
 sky130_fd_sc_hd__buf_12 output671 (.A(net671),
    .X(la_data_in_mprj[57]));
 sky130_fd_sc_hd__buf_12 output672 (.A(net672),
    .X(la_data_in_mprj[58]));
 sky130_fd_sc_hd__buf_12 output673 (.A(net673),
    .X(la_data_in_mprj[59]));
 sky130_fd_sc_hd__buf_12 output674 (.A(net674),
    .X(la_data_in_mprj[5]));
 sky130_fd_sc_hd__buf_12 output675 (.A(net675),
    .X(la_data_in_mprj[60]));
 sky130_fd_sc_hd__buf_12 output676 (.A(net676),
    .X(la_data_in_mprj[61]));
 sky130_fd_sc_hd__buf_12 output677 (.A(net677),
    .X(la_data_in_mprj[62]));
 sky130_fd_sc_hd__buf_12 output678 (.A(net678),
    .X(la_data_in_mprj[63]));
 sky130_fd_sc_hd__buf_12 output679 (.A(net679),
    .X(la_data_in_mprj[64]));
 sky130_fd_sc_hd__buf_12 output680 (.A(net680),
    .X(la_data_in_mprj[65]));
 sky130_fd_sc_hd__buf_12 output681 (.A(net681),
    .X(la_data_in_mprj[66]));
 sky130_fd_sc_hd__buf_12 output682 (.A(net682),
    .X(la_data_in_mprj[67]));
 sky130_fd_sc_hd__buf_12 output683 (.A(net683),
    .X(la_data_in_mprj[68]));
 sky130_fd_sc_hd__buf_12 output684 (.A(net684),
    .X(la_data_in_mprj[69]));
 sky130_fd_sc_hd__buf_12 output685 (.A(net685),
    .X(la_data_in_mprj[6]));
 sky130_fd_sc_hd__buf_12 output686 (.A(net686),
    .X(la_data_in_mprj[70]));
 sky130_fd_sc_hd__buf_12 output687 (.A(net687),
    .X(la_data_in_mprj[71]));
 sky130_fd_sc_hd__buf_12 output688 (.A(net688),
    .X(la_data_in_mprj[72]));
 sky130_fd_sc_hd__buf_12 output689 (.A(net689),
    .X(la_data_in_mprj[73]));
 sky130_fd_sc_hd__buf_12 output690 (.A(net690),
    .X(la_data_in_mprj[74]));
 sky130_fd_sc_hd__buf_12 output691 (.A(net691),
    .X(la_data_in_mprj[75]));
 sky130_fd_sc_hd__buf_12 output692 (.A(net692),
    .X(la_data_in_mprj[76]));
 sky130_fd_sc_hd__buf_12 output693 (.A(net693),
    .X(la_data_in_mprj[77]));
 sky130_fd_sc_hd__buf_12 output694 (.A(net694),
    .X(la_data_in_mprj[78]));
 sky130_fd_sc_hd__buf_12 output695 (.A(net695),
    .X(la_data_in_mprj[79]));
 sky130_fd_sc_hd__buf_12 output696 (.A(net696),
    .X(la_data_in_mprj[7]));
 sky130_fd_sc_hd__buf_12 output697 (.A(net697),
    .X(la_data_in_mprj[80]));
 sky130_fd_sc_hd__buf_12 output698 (.A(net698),
    .X(la_data_in_mprj[81]));
 sky130_fd_sc_hd__buf_12 output699 (.A(net699),
    .X(la_data_in_mprj[82]));
 sky130_fd_sc_hd__buf_12 output700 (.A(net700),
    .X(la_data_in_mprj[83]));
 sky130_fd_sc_hd__buf_12 output701 (.A(net701),
    .X(la_data_in_mprj[84]));
 sky130_fd_sc_hd__buf_12 output702 (.A(net702),
    .X(la_data_in_mprj[85]));
 sky130_fd_sc_hd__buf_12 output703 (.A(net703),
    .X(la_data_in_mprj[86]));
 sky130_fd_sc_hd__buf_12 output704 (.A(net704),
    .X(la_data_in_mprj[87]));
 sky130_fd_sc_hd__buf_12 output705 (.A(net705),
    .X(la_data_in_mprj[88]));
 sky130_fd_sc_hd__buf_12 output706 (.A(net706),
    .X(la_data_in_mprj[89]));
 sky130_fd_sc_hd__buf_12 output707 (.A(net707),
    .X(la_data_in_mprj[8]));
 sky130_fd_sc_hd__buf_12 output708 (.A(net708),
    .X(la_data_in_mprj[90]));
 sky130_fd_sc_hd__buf_12 output709 (.A(net709),
    .X(la_data_in_mprj[91]));
 sky130_fd_sc_hd__buf_12 output710 (.A(net710),
    .X(la_data_in_mprj[92]));
 sky130_fd_sc_hd__buf_12 output711 (.A(net711),
    .X(la_data_in_mprj[93]));
 sky130_fd_sc_hd__buf_12 output712 (.A(net712),
    .X(la_data_in_mprj[94]));
 sky130_fd_sc_hd__buf_12 output713 (.A(net713),
    .X(la_data_in_mprj[95]));
 sky130_fd_sc_hd__buf_12 output714 (.A(net714),
    .X(la_data_in_mprj[96]));
 sky130_fd_sc_hd__buf_12 output715 (.A(net715),
    .X(la_data_in_mprj[97]));
 sky130_fd_sc_hd__buf_12 output716 (.A(net716),
    .X(la_data_in_mprj[98]));
 sky130_fd_sc_hd__buf_12 output717 (.A(net717),
    .X(la_data_in_mprj[99]));
 sky130_fd_sc_hd__buf_12 output718 (.A(net718),
    .X(la_data_in_mprj[9]));
 sky130_fd_sc_hd__buf_12 output719 (.A(net1095),
    .X(la_oenb_core[0]));
 sky130_fd_sc_hd__buf_12 output720 (.A(net720),
    .X(la_oenb_core[100]));
 sky130_fd_sc_hd__buf_12 output721 (.A(net721),
    .X(la_oenb_core[101]));
 sky130_fd_sc_hd__buf_12 output722 (.A(net722),
    .X(la_oenb_core[102]));
 sky130_fd_sc_hd__buf_12 output723 (.A(net723),
    .X(la_oenb_core[103]));
 sky130_fd_sc_hd__buf_12 output724 (.A(net724),
    .X(la_oenb_core[104]));
 sky130_fd_sc_hd__buf_12 output725 (.A(net725),
    .X(la_oenb_core[105]));
 sky130_fd_sc_hd__buf_12 output726 (.A(net726),
    .X(la_oenb_core[106]));
 sky130_fd_sc_hd__buf_12 output727 (.A(net727),
    .X(la_oenb_core[107]));
 sky130_fd_sc_hd__buf_12 output728 (.A(net728),
    .X(la_oenb_core[108]));
 sky130_fd_sc_hd__buf_12 output729 (.A(net729),
    .X(la_oenb_core[109]));
 sky130_fd_sc_hd__buf_12 output730 (.A(net730),
    .X(la_oenb_core[10]));
 sky130_fd_sc_hd__buf_12 output731 (.A(net731),
    .X(la_oenb_core[110]));
 sky130_fd_sc_hd__buf_12 output732 (.A(net732),
    .X(la_oenb_core[111]));
 sky130_fd_sc_hd__buf_12 output733 (.A(net733),
    .X(la_oenb_core[112]));
 sky130_fd_sc_hd__buf_12 output734 (.A(net734),
    .X(la_oenb_core[113]));
 sky130_fd_sc_hd__buf_12 output735 (.A(net735),
    .X(la_oenb_core[114]));
 sky130_fd_sc_hd__buf_12 output736 (.A(net736),
    .X(la_oenb_core[115]));
 sky130_fd_sc_hd__buf_12 output737 (.A(net737),
    .X(la_oenb_core[116]));
 sky130_fd_sc_hd__buf_12 output738 (.A(net738),
    .X(la_oenb_core[117]));
 sky130_fd_sc_hd__buf_12 output739 (.A(net739),
    .X(la_oenb_core[118]));
 sky130_fd_sc_hd__buf_12 output740 (.A(net740),
    .X(la_oenb_core[119]));
 sky130_fd_sc_hd__buf_12 output741 (.A(net741),
    .X(la_oenb_core[11]));
 sky130_fd_sc_hd__buf_12 output742 (.A(net742),
    .X(la_oenb_core[120]));
 sky130_fd_sc_hd__buf_12 output743 (.A(net743),
    .X(la_oenb_core[121]));
 sky130_fd_sc_hd__buf_12 output744 (.A(net744),
    .X(la_oenb_core[122]));
 sky130_fd_sc_hd__buf_12 output745 (.A(net745),
    .X(la_oenb_core[123]));
 sky130_fd_sc_hd__buf_12 output746 (.A(net746),
    .X(la_oenb_core[124]));
 sky130_fd_sc_hd__buf_12 output747 (.A(net747),
    .X(la_oenb_core[125]));
 sky130_fd_sc_hd__buf_12 output748 (.A(net748),
    .X(la_oenb_core[126]));
 sky130_fd_sc_hd__buf_12 output749 (.A(net749),
    .X(la_oenb_core[127]));
 sky130_fd_sc_hd__buf_12 output750 (.A(net750),
    .X(la_oenb_core[12]));
 sky130_fd_sc_hd__buf_12 output751 (.A(net751),
    .X(la_oenb_core[13]));
 sky130_fd_sc_hd__buf_12 output752 (.A(net752),
    .X(la_oenb_core[14]));
 sky130_fd_sc_hd__buf_12 output753 (.A(net753),
    .X(la_oenb_core[15]));
 sky130_fd_sc_hd__buf_12 output754 (.A(net754),
    .X(la_oenb_core[16]));
 sky130_fd_sc_hd__buf_12 output755 (.A(net755),
    .X(la_oenb_core[17]));
 sky130_fd_sc_hd__buf_12 output756 (.A(net756),
    .X(la_oenb_core[18]));
 sky130_fd_sc_hd__buf_12 output757 (.A(net757),
    .X(la_oenb_core[19]));
 sky130_fd_sc_hd__buf_12 output758 (.A(net758),
    .X(la_oenb_core[1]));
 sky130_fd_sc_hd__buf_12 output759 (.A(net759),
    .X(la_oenb_core[20]));
 sky130_fd_sc_hd__buf_12 output760 (.A(net760),
    .X(la_oenb_core[21]));
 sky130_fd_sc_hd__buf_12 output761 (.A(net761),
    .X(la_oenb_core[22]));
 sky130_fd_sc_hd__buf_12 output762 (.A(net762),
    .X(la_oenb_core[23]));
 sky130_fd_sc_hd__buf_12 output763 (.A(net763),
    .X(la_oenb_core[24]));
 sky130_fd_sc_hd__buf_12 output764 (.A(net764),
    .X(la_oenb_core[25]));
 sky130_fd_sc_hd__buf_12 output765 (.A(net765),
    .X(la_oenb_core[26]));
 sky130_fd_sc_hd__buf_12 output766 (.A(net1093),
    .X(la_oenb_core[27]));
 sky130_fd_sc_hd__buf_12 output767 (.A(net767),
    .X(la_oenb_core[28]));
 sky130_fd_sc_hd__buf_12 output768 (.A(net768),
    .X(la_oenb_core[29]));
 sky130_fd_sc_hd__buf_12 output769 (.A(net769),
    .X(la_oenb_core[2]));
 sky130_fd_sc_hd__buf_12 output770 (.A(net770),
    .X(la_oenb_core[30]));
 sky130_fd_sc_hd__buf_12 output771 (.A(net771),
    .X(la_oenb_core[31]));
 sky130_fd_sc_hd__buf_12 output772 (.A(net772),
    .X(la_oenb_core[32]));
 sky130_fd_sc_hd__buf_12 output773 (.A(net773),
    .X(la_oenb_core[33]));
 sky130_fd_sc_hd__buf_12 output774 (.A(net774),
    .X(la_oenb_core[34]));
 sky130_fd_sc_hd__buf_12 output775 (.A(net775),
    .X(la_oenb_core[35]));
 sky130_fd_sc_hd__buf_12 output776 (.A(net776),
    .X(la_oenb_core[36]));
 sky130_fd_sc_hd__buf_12 output777 (.A(net777),
    .X(la_oenb_core[37]));
 sky130_fd_sc_hd__buf_12 output778 (.A(net778),
    .X(la_oenb_core[38]));
 sky130_fd_sc_hd__buf_12 output779 (.A(net1092),
    .X(la_oenb_core[39]));
 sky130_fd_sc_hd__buf_12 output780 (.A(net780),
    .X(la_oenb_core[3]));
 sky130_fd_sc_hd__buf_12 output781 (.A(net781),
    .X(la_oenb_core[40]));
 sky130_fd_sc_hd__buf_12 output782 (.A(net782),
    .X(la_oenb_core[41]));
 sky130_fd_sc_hd__buf_12 output783 (.A(net783),
    .X(la_oenb_core[42]));
 sky130_fd_sc_hd__buf_12 output784 (.A(net784),
    .X(la_oenb_core[43]));
 sky130_fd_sc_hd__buf_12 output785 (.A(net785),
    .X(la_oenb_core[44]));
 sky130_fd_sc_hd__buf_12 output786 (.A(net1091),
    .X(la_oenb_core[45]));
 sky130_fd_sc_hd__buf_12 output787 (.A(net787),
    .X(la_oenb_core[46]));
 sky130_fd_sc_hd__buf_12 output788 (.A(net788),
    .X(la_oenb_core[47]));
 sky130_fd_sc_hd__buf_12 output789 (.A(net789),
    .X(la_oenb_core[48]));
 sky130_fd_sc_hd__buf_12 output790 (.A(net790),
    .X(la_oenb_core[49]));
 sky130_fd_sc_hd__buf_12 output791 (.A(net1094),
    .X(la_oenb_core[4]));
 sky130_fd_sc_hd__buf_12 output792 (.A(net792),
    .X(la_oenb_core[50]));
 sky130_fd_sc_hd__buf_12 output793 (.A(net793),
    .X(la_oenb_core[51]));
 sky130_fd_sc_hd__buf_12 output794 (.A(net794),
    .X(la_oenb_core[52]));
 sky130_fd_sc_hd__buf_12 output795 (.A(net795),
    .X(la_oenb_core[53]));
 sky130_fd_sc_hd__buf_12 output796 (.A(net796),
    .X(la_oenb_core[54]));
 sky130_fd_sc_hd__buf_12 output797 (.A(net797),
    .X(la_oenb_core[55]));
 sky130_fd_sc_hd__buf_12 output798 (.A(net798),
    .X(la_oenb_core[56]));
 sky130_fd_sc_hd__buf_12 output799 (.A(net799),
    .X(la_oenb_core[57]));
 sky130_fd_sc_hd__buf_12 output800 (.A(net800),
    .X(la_oenb_core[58]));
 sky130_fd_sc_hd__buf_12 output801 (.A(net801),
    .X(la_oenb_core[59]));
 sky130_fd_sc_hd__buf_12 output802 (.A(net802),
    .X(la_oenb_core[5]));
 sky130_fd_sc_hd__buf_12 output803 (.A(net803),
    .X(la_oenb_core[60]));
 sky130_fd_sc_hd__buf_12 output804 (.A(net804),
    .X(la_oenb_core[61]));
 sky130_fd_sc_hd__buf_12 output805 (.A(net805),
    .X(la_oenb_core[62]));
 sky130_fd_sc_hd__buf_12 output806 (.A(net806),
    .X(la_oenb_core[63]));
 sky130_fd_sc_hd__buf_12 output807 (.A(net807),
    .X(la_oenb_core[64]));
 sky130_fd_sc_hd__buf_12 output808 (.A(net808),
    .X(la_oenb_core[65]));
 sky130_fd_sc_hd__buf_12 output809 (.A(net809),
    .X(la_oenb_core[66]));
 sky130_fd_sc_hd__buf_12 output810 (.A(net810),
    .X(la_oenb_core[67]));
 sky130_fd_sc_hd__buf_12 output811 (.A(net811),
    .X(la_oenb_core[68]));
 sky130_fd_sc_hd__buf_12 output812 (.A(net812),
    .X(la_oenb_core[69]));
 sky130_fd_sc_hd__buf_12 output813 (.A(net813),
    .X(la_oenb_core[6]));
 sky130_fd_sc_hd__buf_12 output814 (.A(net814),
    .X(la_oenb_core[70]));
 sky130_fd_sc_hd__buf_12 output815 (.A(net815),
    .X(la_oenb_core[71]));
 sky130_fd_sc_hd__buf_12 output816 (.A(net816),
    .X(la_oenb_core[72]));
 sky130_fd_sc_hd__buf_12 output817 (.A(net1090),
    .X(la_oenb_core[73]));
 sky130_fd_sc_hd__buf_12 output818 (.A(net818),
    .X(la_oenb_core[74]));
 sky130_fd_sc_hd__buf_12 output819 (.A(net819),
    .X(la_oenb_core[75]));
 sky130_fd_sc_hd__buf_12 output820 (.A(net820),
    .X(la_oenb_core[76]));
 sky130_fd_sc_hd__buf_12 output821 (.A(net821),
    .X(la_oenb_core[77]));
 sky130_fd_sc_hd__buf_12 output822 (.A(net822),
    .X(la_oenb_core[78]));
 sky130_fd_sc_hd__buf_12 output823 (.A(net823),
    .X(la_oenb_core[79]));
 sky130_fd_sc_hd__buf_12 output824 (.A(net824),
    .X(la_oenb_core[7]));
 sky130_fd_sc_hd__buf_12 output825 (.A(net825),
    .X(la_oenb_core[80]));
 sky130_fd_sc_hd__buf_12 output826 (.A(net1089),
    .X(la_oenb_core[81]));
 sky130_fd_sc_hd__buf_12 output827 (.A(net827),
    .X(la_oenb_core[82]));
 sky130_fd_sc_hd__buf_12 output828 (.A(net828),
    .X(la_oenb_core[83]));
 sky130_fd_sc_hd__buf_12 output829 (.A(net829),
    .X(la_oenb_core[84]));
 sky130_fd_sc_hd__buf_12 output830 (.A(net830),
    .X(la_oenb_core[85]));
 sky130_fd_sc_hd__buf_12 output831 (.A(net831),
    .X(la_oenb_core[86]));
 sky130_fd_sc_hd__buf_12 output832 (.A(net1088),
    .X(la_oenb_core[87]));
 sky130_fd_sc_hd__buf_12 output833 (.A(net1087),
    .X(la_oenb_core[88]));
 sky130_fd_sc_hd__buf_12 output834 (.A(net834),
    .X(la_oenb_core[89]));
 sky130_fd_sc_hd__buf_12 output835 (.A(net835),
    .X(la_oenb_core[8]));
 sky130_fd_sc_hd__buf_12 output836 (.A(net836),
    .X(la_oenb_core[90]));
 sky130_fd_sc_hd__buf_12 output837 (.A(net837),
    .X(la_oenb_core[91]));
 sky130_fd_sc_hd__buf_12 output838 (.A(net838),
    .X(la_oenb_core[92]));
 sky130_fd_sc_hd__buf_12 output839 (.A(net839),
    .X(la_oenb_core[93]));
 sky130_fd_sc_hd__buf_12 output840 (.A(net840),
    .X(la_oenb_core[94]));
 sky130_fd_sc_hd__buf_12 output841 (.A(net841),
    .X(la_oenb_core[95]));
 sky130_fd_sc_hd__buf_12 output842 (.A(net842),
    .X(la_oenb_core[96]));
 sky130_fd_sc_hd__buf_12 output843 (.A(net843),
    .X(la_oenb_core[97]));
 sky130_fd_sc_hd__buf_12 output844 (.A(net844),
    .X(la_oenb_core[98]));
 sky130_fd_sc_hd__buf_12 output845 (.A(net845),
    .X(la_oenb_core[99]));
 sky130_fd_sc_hd__buf_12 output846 (.A(net846),
    .X(la_oenb_core[9]));
 sky130_fd_sc_hd__buf_12 output847 (.A(net847),
    .X(mprj_ack_i_core));
 sky130_fd_sc_hd__buf_12 output848 (.A(net1291),
    .X(mprj_adr_o_user[0]));
 sky130_fd_sc_hd__buf_12 output849 (.A(net1277),
    .X(mprj_adr_o_user[10]));
 sky130_fd_sc_hd__buf_12 output850 (.A(net1274),
    .X(mprj_adr_o_user[11]));
 sky130_fd_sc_hd__buf_12 output851 (.A(net1272),
    .X(mprj_adr_o_user[12]));
 sky130_fd_sc_hd__buf_12 output852 (.A(net1270),
    .X(mprj_adr_o_user[13]));
 sky130_fd_sc_hd__buf_12 output853 (.A(net1267),
    .X(mprj_adr_o_user[14]));
 sky130_fd_sc_hd__buf_12 output854 (.A(net1266),
    .X(mprj_adr_o_user[15]));
 sky130_fd_sc_hd__buf_12 output855 (.A(net855),
    .X(mprj_adr_o_user[16]));
 sky130_fd_sc_hd__buf_12 output856 (.A(net1263),
    .X(mprj_adr_o_user[17]));
 sky130_fd_sc_hd__buf_12 output857 (.A(net857),
    .X(mprj_adr_o_user[18]));
 sky130_fd_sc_hd__buf_12 output858 (.A(net1262),
    .X(mprj_adr_o_user[19]));
 sky130_fd_sc_hd__buf_12 output859 (.A(net1290),
    .X(mprj_adr_o_user[1]));
 sky130_fd_sc_hd__buf_12 output860 (.A(net1260),
    .X(mprj_adr_o_user[20]));
 sky130_fd_sc_hd__buf_12 output861 (.A(net861),
    .X(mprj_adr_o_user[21]));
 sky130_fd_sc_hd__buf_12 output862 (.A(net1257),
    .X(mprj_adr_o_user[22]));
 sky130_fd_sc_hd__buf_12 output863 (.A(net1255),
    .X(mprj_adr_o_user[23]));
 sky130_fd_sc_hd__buf_12 output864 (.A(net864),
    .X(mprj_adr_o_user[24]));
 sky130_fd_sc_hd__buf_12 output865 (.A(net865),
    .X(mprj_adr_o_user[25]));
 sky130_fd_sc_hd__buf_12 output866 (.A(net1254),
    .X(mprj_adr_o_user[26]));
 sky130_fd_sc_hd__buf_12 output867 (.A(net1253),
    .X(mprj_adr_o_user[27]));
 sky130_fd_sc_hd__buf_12 output868 (.A(net1252),
    .X(mprj_adr_o_user[28]));
 sky130_fd_sc_hd__buf_12 output869 (.A(net1251),
    .X(mprj_adr_o_user[29]));
 sky130_fd_sc_hd__buf_12 output870 (.A(net870),
    .X(mprj_adr_o_user[2]));
 sky130_fd_sc_hd__buf_12 output871 (.A(net1249),
    .X(mprj_adr_o_user[30]));
 sky130_fd_sc_hd__buf_12 output872 (.A(net1247),
    .X(mprj_adr_o_user[31]));
 sky130_fd_sc_hd__buf_12 output873 (.A(net1289),
    .X(mprj_adr_o_user[3]));
 sky130_fd_sc_hd__buf_12 output874 (.A(net874),
    .X(mprj_adr_o_user[4]));
 sky130_fd_sc_hd__buf_12 output875 (.A(net1287),
    .X(mprj_adr_o_user[5]));
 sky130_fd_sc_hd__buf_12 output876 (.A(net1284),
    .X(mprj_adr_o_user[6]));
 sky130_fd_sc_hd__buf_12 output877 (.A(net877),
    .X(mprj_adr_o_user[7]));
 sky130_fd_sc_hd__buf_12 output878 (.A(net878),
    .X(mprj_adr_o_user[8]));
 sky130_fd_sc_hd__buf_12 output879 (.A(net1281),
    .X(mprj_adr_o_user[9]));
 sky130_fd_sc_hd__buf_12 output880 (.A(net1319),
    .X(mprj_cyc_o_user));
 sky130_fd_sc_hd__buf_12 output881 (.A(net881),
    .X(mprj_dat_i_core[0]));
 sky130_fd_sc_hd__buf_12 output882 (.A(net882),
    .X(mprj_dat_i_core[10]));
 sky130_fd_sc_hd__buf_12 output883 (.A(net883),
    .X(mprj_dat_i_core[11]));
 sky130_fd_sc_hd__buf_12 output884 (.A(net884),
    .X(mprj_dat_i_core[12]));
 sky130_fd_sc_hd__buf_12 output885 (.A(net885),
    .X(mprj_dat_i_core[13]));
 sky130_fd_sc_hd__buf_12 output886 (.A(net886),
    .X(mprj_dat_i_core[14]));
 sky130_fd_sc_hd__buf_12 output887 (.A(net887),
    .X(mprj_dat_i_core[15]));
 sky130_fd_sc_hd__buf_12 output888 (.A(net888),
    .X(mprj_dat_i_core[16]));
 sky130_fd_sc_hd__buf_12 output889 (.A(net889),
    .X(mprj_dat_i_core[17]));
 sky130_fd_sc_hd__buf_12 output890 (.A(net890),
    .X(mprj_dat_i_core[18]));
 sky130_fd_sc_hd__buf_12 output891 (.A(net891),
    .X(mprj_dat_i_core[19]));
 sky130_fd_sc_hd__buf_12 output892 (.A(net892),
    .X(mprj_dat_i_core[1]));
 sky130_fd_sc_hd__buf_12 output893 (.A(net893),
    .X(mprj_dat_i_core[20]));
 sky130_fd_sc_hd__buf_12 output894 (.A(net894),
    .X(mprj_dat_i_core[21]));
 sky130_fd_sc_hd__buf_12 output895 (.A(net895),
    .X(mprj_dat_i_core[22]));
 sky130_fd_sc_hd__buf_12 output896 (.A(net896),
    .X(mprj_dat_i_core[23]));
 sky130_fd_sc_hd__buf_12 output897 (.A(net897),
    .X(mprj_dat_i_core[24]));
 sky130_fd_sc_hd__buf_12 output898 (.A(net898),
    .X(mprj_dat_i_core[25]));
 sky130_fd_sc_hd__buf_12 output899 (.A(net899),
    .X(mprj_dat_i_core[26]));
 sky130_fd_sc_hd__buf_12 output900 (.A(net900),
    .X(mprj_dat_i_core[27]));
 sky130_fd_sc_hd__buf_12 output901 (.A(net901),
    .X(mprj_dat_i_core[28]));
 sky130_fd_sc_hd__buf_12 output902 (.A(net902),
    .X(mprj_dat_i_core[29]));
 sky130_fd_sc_hd__buf_12 output903 (.A(net965),
    .X(mprj_dat_i_core[2]));
 sky130_fd_sc_hd__buf_12 output904 (.A(net904),
    .X(mprj_dat_i_core[30]));
 sky130_fd_sc_hd__buf_12 output905 (.A(net905),
    .X(mprj_dat_i_core[31]));
 sky130_fd_sc_hd__buf_12 output906 (.A(net906),
    .X(mprj_dat_i_core[3]));
 sky130_fd_sc_hd__buf_12 output907 (.A(net964),
    .X(mprj_dat_i_core[4]));
 sky130_fd_sc_hd__buf_12 output908 (.A(net908),
    .X(mprj_dat_i_core[5]));
 sky130_fd_sc_hd__buf_12 output909 (.A(net909),
    .X(mprj_dat_i_core[6]));
 sky130_fd_sc_hd__buf_12 output910 (.A(net963),
    .X(mprj_dat_i_core[7]));
 sky130_fd_sc_hd__buf_12 output911 (.A(net911),
    .X(mprj_dat_i_core[8]));
 sky130_fd_sc_hd__buf_12 output912 (.A(net912),
    .X(mprj_dat_i_core[9]));
 sky130_fd_sc_hd__buf_12 output913 (.A(net1244),
    .X(mprj_dat_o_user[0]));
 sky130_fd_sc_hd__buf_12 output914 (.A(net1211),
    .X(mprj_dat_o_user[10]));
 sky130_fd_sc_hd__buf_12 output915 (.A(net1208),
    .X(mprj_dat_o_user[11]));
 sky130_fd_sc_hd__buf_12 output916 (.A(net1204),
    .X(mprj_dat_o_user[12]));
 sky130_fd_sc_hd__buf_12 output917 (.A(net1200),
    .X(mprj_dat_o_user[13]));
 sky130_fd_sc_hd__buf_12 output918 (.A(net1197),
    .X(mprj_dat_o_user[14]));
 sky130_fd_sc_hd__buf_12 output919 (.A(net1194),
    .X(mprj_dat_o_user[15]));
 sky130_fd_sc_hd__buf_12 output920 (.A(net1191),
    .X(mprj_dat_o_user[16]));
 sky130_fd_sc_hd__buf_12 output921 (.A(net1188),
    .X(mprj_dat_o_user[17]));
 sky130_fd_sc_hd__buf_12 output922 (.A(net1186),
    .X(mprj_dat_o_user[18]));
 sky130_fd_sc_hd__buf_12 output923 (.A(net1183),
    .X(mprj_dat_o_user[19]));
 sky130_fd_sc_hd__buf_12 output924 (.A(net1241),
    .X(mprj_dat_o_user[1]));
 sky130_fd_sc_hd__buf_12 output925 (.A(net1180),
    .X(mprj_dat_o_user[20]));
 sky130_fd_sc_hd__buf_12 output926 (.A(net1177),
    .X(mprj_dat_o_user[21]));
 sky130_fd_sc_hd__buf_12 output927 (.A(net1174),
    .X(mprj_dat_o_user[22]));
 sky130_fd_sc_hd__buf_12 output928 (.A(net1171),
    .X(mprj_dat_o_user[23]));
 sky130_fd_sc_hd__buf_12 output929 (.A(net1168),
    .X(mprj_dat_o_user[24]));
 sky130_fd_sc_hd__buf_12 output930 (.A(net1165),
    .X(mprj_dat_o_user[25]));
 sky130_fd_sc_hd__buf_12 output931 (.A(net1162),
    .X(mprj_dat_o_user[26]));
 sky130_fd_sc_hd__buf_12 output932 (.A(net1159),
    .X(mprj_dat_o_user[27]));
 sky130_fd_sc_hd__buf_12 output933 (.A(net1156),
    .X(mprj_dat_o_user[28]));
 sky130_fd_sc_hd__buf_12 output934 (.A(net1153),
    .X(mprj_dat_o_user[29]));
 sky130_fd_sc_hd__buf_12 output935 (.A(net1238),
    .X(mprj_dat_o_user[2]));
 sky130_fd_sc_hd__buf_12 output936 (.A(net1151),
    .X(mprj_dat_o_user[30]));
 sky130_fd_sc_hd__buf_12 output937 (.A(net1149),
    .X(mprj_dat_o_user[31]));
 sky130_fd_sc_hd__buf_12 output938 (.A(net1235),
    .X(mprj_dat_o_user[3]));
 sky130_fd_sc_hd__buf_12 output939 (.A(net1232),
    .X(mprj_dat_o_user[4]));
 sky130_fd_sc_hd__buf_12 output940 (.A(net1228),
    .X(mprj_dat_o_user[5]));
 sky130_fd_sc_hd__buf_12 output941 (.A(net1224),
    .X(mprj_dat_o_user[6]));
 sky130_fd_sc_hd__buf_12 output942 (.A(net1221),
    .X(mprj_dat_o_user[7]));
 sky130_fd_sc_hd__buf_12 output943 (.A(net1217),
    .X(mprj_dat_o_user[8]));
 sky130_fd_sc_hd__buf_12 output944 (.A(net1214),
    .X(mprj_dat_o_user[9]));
 sky130_fd_sc_hd__buf_12 output945 (.A(net1306),
    .X(mprj_sel_o_user[0]));
 sky130_fd_sc_hd__buf_12 output946 (.A(net1301),
    .X(mprj_sel_o_user[1]));
 sky130_fd_sc_hd__buf_12 output947 (.A(net1296),
    .X(mprj_sel_o_user[2]));
 sky130_fd_sc_hd__buf_12 output948 (.A(net1292),
    .X(mprj_sel_o_user[3]));
 sky130_fd_sc_hd__buf_12 output949 (.A(net1315),
    .X(mprj_stb_o_user));
 sky130_fd_sc_hd__buf_12 output950 (.A(net1311),
    .X(mprj_we_o_user));
 sky130_fd_sc_hd__buf_12 output951 (.A(net2214),
    .X(user1_vcc_powergood));
 sky130_fd_sc_hd__buf_12 output952 (.A(net2070),
    .X(user1_vdd_powergood));
 sky130_fd_sc_hd__buf_12 output953 (.A(net2850),
    .X(user2_vcc_powergood));
 sky130_fd_sc_hd__buf_12 output954 (.A(net2072),
    .X(user2_vdd_powergood));
 sky130_fd_sc_hd__buf_12 output955 (.A(net1322),
    .X(user_clock));
 sky130_fd_sc_hd__buf_12 output956 (.A(net956),
    .X(user_clock2));
 sky130_fd_sc_hd__buf_12 output957 (.A(net957),
    .X(user_irq[0]));
 sky130_fd_sc_hd__buf_12 output958 (.A(net958),
    .X(user_irq[1]));
 sky130_fd_sc_hd__buf_12 output959 (.A(net959),
    .X(user_irq[2]));
 sky130_fd_sc_hd__buf_12 output960 (.A(net960),
    .X(user_reset));
 sky130_fd_sc_hd__buf_2 wire961 (.A(net625),
    .X(net961));
 sky130_fd_sc_hd__buf_2 wire962 (.A(net602),
    .X(net962));
 sky130_fd_sc_hd__buf_2 wire963 (.A(net910),
    .X(net963));
 sky130_fd_sc_hd__buf_2 wire964 (.A(net907),
    .X(net964));
 sky130_fd_sc_hd__buf_2 wire965 (.A(net903),
    .X(net965));
 sky130_fd_sc_hd__buf_2 wire966 (.A(net619),
    .X(net966));
 sky130_fd_sc_hd__buf_2 wire967 (.A(net617),
    .X(net967));
 sky130_fd_sc_hd__buf_2 wire968 (.A(net616),
    .X(net968));
 sky130_fd_sc_hd__buf_2 wire969 (.A(net615),
    .X(net969));
 sky130_fd_sc_hd__buf_2 wire970 (.A(net614),
    .X(net970));
 sky130_fd_sc_hd__buf_2 wire971 (.A(net611),
    .X(net971));
 sky130_fd_sc_hd__buf_4 wire972 (.A(net973),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 wire973 (.A(net610),
    .X(net973));
 sky130_fd_sc_hd__buf_4 wire974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_2 wire975 (.A(net609),
    .X(net975));
 sky130_fd_sc_hd__buf_4 wire976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_2 wire977 (.A(net608),
    .X(net977));
 sky130_fd_sc_hd__buf_4 wire978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_2 wire979 (.A(net607),
    .X(net979));
 sky130_fd_sc_hd__buf_4 wire980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_2 wire981 (.A(net606),
    .X(net981));
 sky130_fd_sc_hd__buf_4 wire982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_2 wire983 (.A(net605),
    .X(net983));
 sky130_fd_sc_hd__buf_4 wire984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_2 wire985 (.A(net604),
    .X(net985));
 sky130_fd_sc_hd__buf_4 wire986 (.A(net603),
    .X(net986));
 sky130_fd_sc_hd__buf_4 wire987 (.A(net988),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_2 wire988 (.A(net601),
    .X(net988));
 sky130_fd_sc_hd__buf_2 wire989 (.A(net600),
    .X(net989));
 sky130_fd_sc_hd__buf_2 wire990 (.A(net599),
    .X(net990));
 sky130_fd_sc_hd__buf_4 wire991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_2 wire992 (.A(net598),
    .X(net992));
 sky130_fd_sc_hd__buf_2 wire993 (.A(net596),
    .X(net993));
 sky130_fd_sc_hd__buf_2 wire994 (.A(net666),
    .X(net994));
 sky130_fd_sc_hd__buf_2 wire995 (.A(net665),
    .X(net995));
 sky130_fd_sc_hd__buf_2 wire996 (.A(net660),
    .X(net996));
 sky130_fd_sc_hd__buf_2 wire997 (.A(net658),
    .X(net997));
 sky130_fd_sc_hd__buf_2 wire998 (.A(net655),
    .X(net998));
 sky130_fd_sc_hd__buf_2 wire999 (.A(net650),
    .X(net999));
 sky130_fd_sc_hd__buf_2 wire1000 (.A(net649),
    .X(net1000));
 sky130_fd_sc_hd__buf_2 wire1001 (.A(net647),
    .X(net1001));
 sky130_fd_sc_hd__buf_2 wire1002 (.A(net646),
    .X(net1002));
 sky130_fd_sc_hd__buf_2 wire1003 (.A(net645),
    .X(net1003));
 sky130_fd_sc_hd__buf_2 wire1004 (.A(net643),
    .X(net1004));
 sky130_fd_sc_hd__buf_2 wire1005 (.A(net642),
    .X(net1005));
 sky130_fd_sc_hd__buf_2 wire1006 (.A(net640),
    .X(net1006));
 sky130_fd_sc_hd__buf_2 wire1007 (.A(net639),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 wire1008 (.A(net637),
    .X(net1008));
 sky130_fd_sc_hd__buf_2 wire1009 (.A(net636),
    .X(net1009));
 sky130_fd_sc_hd__buf_2 wire1010 (.A(net634),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 wire1011 (.A(net631),
    .X(net1011));
 sky130_fd_sc_hd__buf_2 wire1012 (.A(net629),
    .X(net1012));
 sky130_fd_sc_hd__buf_4 wire1013 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_2 wire1014 (.A(\la_data_in_mprj_bar[99] ),
    .X(net1014));
 sky130_fd_sc_hd__buf_4 wire1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_2 wire1016 (.A(\la_data_in_mprj_bar[98] ),
    .X(net1016));
 sky130_fd_sc_hd__buf_4 wire1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_2 wire1018 (.A(\la_data_in_mprj_bar[97] ),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 wire1019 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_2 wire1020 (.A(\la_data_in_mprj_bar[96] ),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 wire1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_2 wire1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_2 wire1023 (.A(\la_data_in_mprj_bar[95] ),
    .X(net1023));
 sky130_fd_sc_hd__buf_4 wire1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_2 wire1025 (.A(\la_data_in_mprj_bar[94] ),
    .X(net1025));
 sky130_fd_sc_hd__buf_4 wire1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_2 wire1027 (.A(\la_data_in_mprj_bar[93] ),
    .X(net1027));
 sky130_fd_sc_hd__buf_4 wire1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_2 wire1029 (.A(\la_data_in_mprj_bar[92] ),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 wire1030 (.A(net1031),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_2 wire1031 (.A(\la_data_in_mprj_bar[91] ),
    .X(net1031));
 sky130_fd_sc_hd__buf_6 wire1032 (.A(net1033),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 wire1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_2 wire1034 (.A(\la_data_in_mprj_bar[90] ),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_2 wire1035 (.A(\la_data_in_mprj_bar[89] ),
    .X(net1035));
 sky130_fd_sc_hd__buf_6 wire1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 wire1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_2 wire1038 (.A(\la_data_in_mprj_bar[88] ),
    .X(net1038));
 sky130_fd_sc_hd__buf_4 wire1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_2 wire1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_2 wire1041 (.A(\la_data_in_mprj_bar[87] ),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_2 wire1042 (.A(net1043),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_2 wire1043 (.A(\la_data_in_mprj_bar[86] ),
    .X(net1043));
 sky130_fd_sc_hd__buf_4 wire1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_2 wire1045 (.A(\la_data_in_mprj_bar[85] ),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 wire1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_2 wire1047 (.A(net1048),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_2 wire1048 (.A(\la_data_in_mprj_bar[84] ),
    .X(net1048));
 sky130_fd_sc_hd__buf_4 wire1049 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_2 wire1050 (.A(\la_data_in_mprj_bar[83] ),
    .X(net1050));
 sky130_fd_sc_hd__buf_4 wire1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_2 wire1052 (.A(\la_data_in_mprj_bar[82] ),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 wire1053 (.A(net1054),
    .X(net1053));
 sky130_fd_sc_hd__buf_4 wire1054 (.A(net1055),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_2 wire1055 (.A(\la_data_in_mprj_bar[81] ),
    .X(net1055));
 sky130_fd_sc_hd__buf_6 wire1056 (.A(net1057),
    .X(net1056));
 sky130_fd_sc_hd__buf_4 wire1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_2 wire1058 (.A(\la_data_in_mprj_bar[80] ),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 wire1059 (.A(net1060),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_2 wire1060 (.A(\la_data_in_mprj_bar[79] ),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 wire1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__clkbuf_2 wire1062 (.A(\la_data_in_mprj_bar[78] ),
    .X(net1062));
 sky130_fd_sc_hd__buf_6 wire1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_4 wire1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__buf_2 wire1065 (.A(net1066),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_2 wire1066 (.A(\la_data_in_mprj_bar[77] ),
    .X(net1066));
 sky130_fd_sc_hd__buf_6 wire1067 (.A(net1068),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 wire1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__clkbuf_2 wire1069 (.A(\la_data_in_mprj_bar[76] ),
    .X(net1069));
 sky130_fd_sc_hd__buf_4 wire1070 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 wire1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_2 wire1072 (.A(\la_data_in_mprj_bar[75] ),
    .X(net1072));
 sky130_fd_sc_hd__buf_4 wire1073 (.A(net1074),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_2 wire1074 (.A(\la_data_in_mprj_bar[74] ),
    .X(net1074));
 sky130_fd_sc_hd__buf_4 wire1075 (.A(net1076),
    .X(net1075));
 sky130_fd_sc_hd__clkbuf_2 wire1076 (.A(\la_data_in_mprj_bar[73] ),
    .X(net1076));
 sky130_fd_sc_hd__buf_4 wire1077 (.A(net1078),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_2 wire1078 (.A(\la_data_in_mprj_bar[72] ),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 wire1079 (.A(\la_data_in_mprj_bar[71] ),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_2 wire1080 (.A(\la_data_in_mprj_bar[70] ),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 wire1081 (.A(net1082),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_2 wire1082 (.A(\la_data_in_mprj_bar[103] ),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_2 wire1083 (.A(\la_data_in_mprj_bar[102] ),
    .X(net1083));
 sky130_fd_sc_hd__buf_4 wire1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_2 wire1085 (.A(\la_data_in_mprj_bar[101] ),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_2 wire1086 (.A(\la_data_in_mprj_bar[100] ),
    .X(net1086));
 sky130_fd_sc_hd__buf_2 wire1087 (.A(net833),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 wire1088 (.A(net832),
    .X(net1088));
 sky130_fd_sc_hd__buf_2 wire1089 (.A(net826),
    .X(net1089));
 sky130_fd_sc_hd__buf_2 wire1090 (.A(net817),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 wire1091 (.A(net786),
    .X(net1091));
 sky130_fd_sc_hd__buf_2 wire1092 (.A(net779),
    .X(net1092));
 sky130_fd_sc_hd__buf_2 wire1093 (.A(net766),
    .X(net1093));
 sky130_fd_sc_hd__buf_2 wire1094 (.A(net791),
    .X(net1094));
 sky130_fd_sc_hd__buf_2 wire1095 (.A(net719),
    .X(net1095));
 sky130_fd_sc_hd__buf_2 wire1096 (.A(net473),
    .X(net1096));
 sky130_fd_sc_hd__buf_2 wire1097 (.A(net471),
    .X(net1097));
 sky130_fd_sc_hd__buf_2 wire1098 (.A(net469),
    .X(net1098));
 sky130_fd_sc_hd__buf_2 wire1099 (.A(net468),
    .X(net1099));
 sky130_fd_sc_hd__buf_2 wire1100 (.A(net467),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 wire1101 (.A(net465),
    .X(net1101));
 sky130_fd_sc_hd__buf_4 wire1102 (.A(net589),
    .X(net1102));
 sky130_fd_sc_hd__buf_4 wire1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_2 wire1104 (.A(net588),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 wire1105 (.A(net586),
    .X(net1105));
 sky130_fd_sc_hd__buf_2 wire1106 (.A(net585),
    .X(net1106));
 sky130_fd_sc_hd__buf_2 wire1107 (.A(net584),
    .X(net1107));
 sky130_fd_sc_hd__buf_2 wire1108 (.A(net583),
    .X(net1108));
 sky130_fd_sc_hd__buf_2 wire1109 (.A(net582),
    .X(net1109));
 sky130_fd_sc_hd__buf_2 wire1110 (.A(net581),
    .X(net1110));
 sky130_fd_sc_hd__buf_2 wire1111 (.A(net578),
    .X(net1111));
 sky130_fd_sc_hd__buf_2 wire1112 (.A(net576),
    .X(net1112));
 sky130_fd_sc_hd__buf_2 wire1113 (.A(net575),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 wire1114 (.A(net573),
    .X(net1114));
 sky130_fd_sc_hd__buf_2 wire1115 (.A(net572),
    .X(net1115));
 sky130_fd_sc_hd__buf_2 wire1116 (.A(net571),
    .X(net1116));
 sky130_fd_sc_hd__buf_2 wire1117 (.A(net570),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 wire1118 (.A(net569),
    .X(net1118));
 sky130_fd_sc_hd__buf_2 wire1119 (.A(net533),
    .X(net1119));
 sky130_fd_sc_hd__buf_4 wire1120 (.A(net525),
    .X(net1120));
 sky130_fd_sc_hd__buf_2 wire1121 (.A(net518),
    .X(net1121));
 sky130_fd_sc_hd__buf_4 wire1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_2 wire1123 (.A(net517),
    .X(net1123));
 sky130_fd_sc_hd__buf_4 wire1124 (.A(net1125),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_2 wire1125 (.A(net516),
    .X(net1125));
 sky130_fd_sc_hd__buf_2 wire1126 (.A(net515),
    .X(net1126));
 sky130_fd_sc_hd__buf_2 wire1127 (.A(net512),
    .X(net1127));
 sky130_fd_sc_hd__buf_2 wire1128 (.A(net511),
    .X(net1128));
 sky130_fd_sc_hd__buf_4 wire1129 (.A(net1130),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_2 wire1130 (.A(net510),
    .X(net1130));
 sky130_fd_sc_hd__buf_2 wire1131 (.A(net509),
    .X(net1131));
 sky130_fd_sc_hd__buf_2 wire1132 (.A(net503),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 wire1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_2 wire1134 (.A(net501),
    .X(net1134));
 sky130_fd_sc_hd__buf_4 wire1135 (.A(net1136),
    .X(net1135));
 sky130_fd_sc_hd__clkbuf_2 wire1136 (.A(net498),
    .X(net1136));
 sky130_fd_sc_hd__buf_2 wire1137 (.A(net495),
    .X(net1137));
 sky130_fd_sc_hd__buf_2 wire1138 (.A(net494),
    .X(net1138));
 sky130_fd_sc_hd__buf_2 wire1139 (.A(net590),
    .X(net1139));
 sky130_fd_sc_hd__buf_2 wire1140 (.A(net568),
    .X(net1140));
 sky130_fd_sc_hd__buf_2 wire1141 (.A(net557),
    .X(net1141));
 sky130_fd_sc_hd__buf_2 wire1142 (.A(net546),
    .X(net1142));
 sky130_fd_sc_hd__buf_2 wire1143 (.A(net535),
    .X(net1143));
 sky130_fd_sc_hd__buf_2 wire1144 (.A(net524),
    .X(net1144));
 sky130_fd_sc_hd__buf_2 wire1145 (.A(net513),
    .X(net1145));
 sky130_fd_sc_hd__buf_4 wire1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_2 wire1147 (.A(net502),
    .X(net1147));
 sky130_fd_sc_hd__buf_2 wire1148 (.A(net463),
    .X(net1148));
 sky130_fd_sc_hd__buf_4 wire1149 (.A(net1150),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_2 wire1150 (.A(net937),
    .X(net1150));
 sky130_fd_sc_hd__buf_4 wire1151 (.A(net1152),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_2 wire1152 (.A(net936),
    .X(net1152));
 sky130_fd_sc_hd__buf_6 wire1153 (.A(net1154),
    .X(net1153));
 sky130_fd_sc_hd__buf_4 wire1154 (.A(net1155),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_2 wire1155 (.A(net934),
    .X(net1155));
 sky130_fd_sc_hd__buf_6 wire1156 (.A(net1157),
    .X(net1156));
 sky130_fd_sc_hd__buf_4 wire1157 (.A(net1158),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_2 wire1158 (.A(net933),
    .X(net1158));
 sky130_fd_sc_hd__buf_6 wire1159 (.A(net1160),
    .X(net1159));
 sky130_fd_sc_hd__buf_4 wire1160 (.A(net1161),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_2 wire1161 (.A(net932),
    .X(net1161));
 sky130_fd_sc_hd__buf_6 wire1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__buf_4 wire1163 (.A(net1164),
    .X(net1163));
 sky130_fd_sc_hd__clkbuf_2 wire1164 (.A(net931),
    .X(net1164));
 sky130_fd_sc_hd__buf_6 wire1165 (.A(net1166),
    .X(net1165));
 sky130_fd_sc_hd__buf_4 wire1166 (.A(net1167),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_2 wire1167 (.A(net930),
    .X(net1167));
 sky130_fd_sc_hd__buf_6 wire1168 (.A(net1169),
    .X(net1168));
 sky130_fd_sc_hd__buf_4 wire1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_2 wire1170 (.A(net929),
    .X(net1170));
 sky130_fd_sc_hd__buf_6 wire1171 (.A(net1172),
    .X(net1171));
 sky130_fd_sc_hd__buf_4 wire1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__clkbuf_2 wire1173 (.A(net928),
    .X(net1173));
 sky130_fd_sc_hd__buf_6 wire1174 (.A(net1175),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_2 wire1175 (.A(net1176),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_2 wire1176 (.A(net927),
    .X(net1176));
 sky130_fd_sc_hd__buf_6 wire1177 (.A(net1178),
    .X(net1177));
 sky130_fd_sc_hd__clkbuf_2 wire1178 (.A(net1179),
    .X(net1178));
 sky130_fd_sc_hd__clkbuf_2 wire1179 (.A(net926),
    .X(net1179));
 sky130_fd_sc_hd__buf_6 wire1180 (.A(net1181),
    .X(net1180));
 sky130_fd_sc_hd__buf_4 wire1181 (.A(net1182),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_2 wire1182 (.A(net925),
    .X(net1182));
 sky130_fd_sc_hd__buf_6 wire1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_2 wire1184 (.A(net1185),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_2 wire1185 (.A(net923),
    .X(net1185));
 sky130_fd_sc_hd__buf_4 wire1186 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_2 wire1187 (.A(net922),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 wire1188 (.A(net1189),
    .X(net1188));
 sky130_fd_sc_hd__buf_4 wire1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__clkbuf_2 wire1190 (.A(net921),
    .X(net1190));
 sky130_fd_sc_hd__buf_6 wire1191 (.A(net1192),
    .X(net1191));
 sky130_fd_sc_hd__buf_4 wire1192 (.A(net1193),
    .X(net1192));
 sky130_fd_sc_hd__clkbuf_2 wire1193 (.A(net920),
    .X(net1193));
 sky130_fd_sc_hd__buf_6 wire1194 (.A(net1195),
    .X(net1194));
 sky130_fd_sc_hd__buf_4 wire1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_2 wire1196 (.A(net919),
    .X(net1196));
 sky130_fd_sc_hd__buf_6 wire1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__buf_4 wire1198 (.A(net1199),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_2 wire1199 (.A(net918),
    .X(net1199));
 sky130_fd_sc_hd__buf_6 wire1200 (.A(net1201),
    .X(net1200));
 sky130_fd_sc_hd__buf_4 wire1201 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_2 wire1202 (.A(net1203),
    .X(net1202));
 sky130_fd_sc_hd__clkbuf_2 wire1203 (.A(net917),
    .X(net1203));
 sky130_fd_sc_hd__buf_6 wire1204 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__buf_4 wire1205 (.A(net1206),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_2 wire1206 (.A(net1207),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_2 wire1207 (.A(net916),
    .X(net1207));
 sky130_fd_sc_hd__buf_6 wire1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_4 wire1209 (.A(net1210),
    .X(net1209));
 sky130_fd_sc_hd__clkbuf_2 wire1210 (.A(net915),
    .X(net1210));
 sky130_fd_sc_hd__buf_6 wire1211 (.A(net1212),
    .X(net1211));
 sky130_fd_sc_hd__buf_4 wire1212 (.A(net1213),
    .X(net1212));
 sky130_fd_sc_hd__clkbuf_2 wire1213 (.A(net914),
    .X(net1213));
 sky130_fd_sc_hd__buf_6 wire1214 (.A(net1215),
    .X(net1214));
 sky130_fd_sc_hd__buf_4 wire1215 (.A(net1216),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_2 wire1216 (.A(net944),
    .X(net1216));
 sky130_fd_sc_hd__buf_6 wire1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__buf_4 wire1218 (.A(net1219),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_2 wire1219 (.A(net1220),
    .X(net1219));
 sky130_fd_sc_hd__clkbuf_2 wire1220 (.A(net943),
    .X(net1220));
 sky130_fd_sc_hd__buf_6 wire1221 (.A(net1222),
    .X(net1221));
 sky130_fd_sc_hd__buf_4 wire1222 (.A(net1223),
    .X(net1222));
 sky130_fd_sc_hd__clkbuf_2 wire1223 (.A(net942),
    .X(net1223));
 sky130_fd_sc_hd__buf_6 wire1224 (.A(net1225),
    .X(net1224));
 sky130_fd_sc_hd__buf_4 wire1225 (.A(net1226),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_2 wire1226 (.A(net1227),
    .X(net1226));
 sky130_fd_sc_hd__clkbuf_2 wire1227 (.A(net941),
    .X(net1227));
 sky130_fd_sc_hd__buf_6 wire1228 (.A(net1229),
    .X(net1228));
 sky130_fd_sc_hd__buf_4 wire1229 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_2 wire1230 (.A(net1231),
    .X(net1230));
 sky130_fd_sc_hd__clkbuf_2 wire1231 (.A(net940),
    .X(net1231));
 sky130_fd_sc_hd__buf_6 wire1232 (.A(net1233),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 wire1233 (.A(net1234),
    .X(net1233));
 sky130_fd_sc_hd__clkbuf_2 wire1234 (.A(net939),
    .X(net1234));
 sky130_fd_sc_hd__buf_6 wire1235 (.A(net1236),
    .X(net1235));
 sky130_fd_sc_hd__buf_4 wire1236 (.A(net1237),
    .X(net1236));
 sky130_fd_sc_hd__clkbuf_2 wire1237 (.A(net938),
    .X(net1237));
 sky130_fd_sc_hd__buf_6 wire1238 (.A(net1239),
    .X(net1238));
 sky130_fd_sc_hd__buf_4 wire1239 (.A(net1240),
    .X(net1239));
 sky130_fd_sc_hd__clkbuf_2 wire1240 (.A(net935),
    .X(net1240));
 sky130_fd_sc_hd__buf_6 wire1241 (.A(net1242),
    .X(net1241));
 sky130_fd_sc_hd__buf_4 wire1242 (.A(net1243),
    .X(net1242));
 sky130_fd_sc_hd__clkbuf_2 wire1243 (.A(net924),
    .X(net1243));
 sky130_fd_sc_hd__buf_6 wire1244 (.A(net1245),
    .X(net1244));
 sky130_fd_sc_hd__buf_4 wire1245 (.A(net1246),
    .X(net1245));
 sky130_fd_sc_hd__clkbuf_2 wire1246 (.A(net913),
    .X(net1246));
 sky130_fd_sc_hd__buf_4 wire1247 (.A(net1248),
    .X(net1247));
 sky130_fd_sc_hd__clkbuf_2 wire1248 (.A(net872),
    .X(net1248));
 sky130_fd_sc_hd__buf_4 wire1249 (.A(net1250),
    .X(net1249));
 sky130_fd_sc_hd__clkbuf_2 wire1250 (.A(net871),
    .X(net1250));
 sky130_fd_sc_hd__buf_2 wire1251 (.A(net869),
    .X(net1251));
 sky130_fd_sc_hd__buf_4 wire1252 (.A(net868),
    .X(net1252));
 sky130_fd_sc_hd__buf_2 wire1253 (.A(net867),
    .X(net1253));
 sky130_fd_sc_hd__buf_2 wire1254 (.A(net866),
    .X(net1254));
 sky130_fd_sc_hd__buf_4 wire1255 (.A(net1256),
    .X(net1255));
 sky130_fd_sc_hd__clkbuf_2 wire1256 (.A(net863),
    .X(net1256));
 sky130_fd_sc_hd__buf_6 wire1257 (.A(net1258),
    .X(net1257));
 sky130_fd_sc_hd__buf_4 wire1258 (.A(net1259),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_2 wire1259 (.A(net862),
    .X(net1259));
 sky130_fd_sc_hd__buf_4 wire1260 (.A(net1261),
    .X(net1260));
 sky130_fd_sc_hd__clkbuf_2 wire1261 (.A(net860),
    .X(net1261));
 sky130_fd_sc_hd__buf_2 wire1262 (.A(net858),
    .X(net1262));
 sky130_fd_sc_hd__buf_6 wire1263 (.A(net1264),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_2 wire1264 (.A(net1265),
    .X(net1264));
 sky130_fd_sc_hd__clkbuf_2 wire1265 (.A(net856),
    .X(net1265));
 sky130_fd_sc_hd__buf_2 wire1266 (.A(net854),
    .X(net1266));
 sky130_fd_sc_hd__buf_6 wire1267 (.A(net1268),
    .X(net1267));
 sky130_fd_sc_hd__clkbuf_2 wire1268 (.A(net1269),
    .X(net1268));
 sky130_fd_sc_hd__clkbuf_2 wire1269 (.A(net853),
    .X(net1269));
 sky130_fd_sc_hd__buf_4 wire1270 (.A(net1271),
    .X(net1270));
 sky130_fd_sc_hd__clkbuf_2 wire1271 (.A(net852),
    .X(net1271));
 sky130_fd_sc_hd__buf_4 wire1272 (.A(net1273),
    .X(net1272));
 sky130_fd_sc_hd__clkbuf_2 wire1273 (.A(net851),
    .X(net1273));
 sky130_fd_sc_hd__buf_6 wire1274 (.A(net1275),
    .X(net1274));
 sky130_fd_sc_hd__buf_4 wire1275 (.A(net1276),
    .X(net1275));
 sky130_fd_sc_hd__clkbuf_2 wire1276 (.A(net850),
    .X(net1276));
 sky130_fd_sc_hd__buf_6 wire1277 (.A(net1278),
    .X(net1277));
 sky130_fd_sc_hd__buf_4 wire1278 (.A(net1279),
    .X(net1278));
 sky130_fd_sc_hd__clkbuf_2 wire1279 (.A(net1280),
    .X(net1279));
 sky130_fd_sc_hd__clkbuf_2 wire1280 (.A(net849),
    .X(net1280));
 sky130_fd_sc_hd__buf_6 wire1281 (.A(net1282),
    .X(net1281));
 sky130_fd_sc_hd__buf_4 wire1282 (.A(net1283),
    .X(net1282));
 sky130_fd_sc_hd__clkbuf_2 wire1283 (.A(net879),
    .X(net1283));
 sky130_fd_sc_hd__buf_6 wire1284 (.A(net1285),
    .X(net1284));
 sky130_fd_sc_hd__clkbuf_2 wire1285 (.A(net1286),
    .X(net1285));
 sky130_fd_sc_hd__clkbuf_2 wire1286 (.A(net876),
    .X(net1286));
 sky130_fd_sc_hd__buf_4 wire1287 (.A(net1288),
    .X(net1287));
 sky130_fd_sc_hd__clkbuf_2 wire1288 (.A(net875),
    .X(net1288));
 sky130_fd_sc_hd__buf_2 wire1289 (.A(net873),
    .X(net1289));
 sky130_fd_sc_hd__buf_2 wire1290 (.A(net859),
    .X(net1290));
 sky130_fd_sc_hd__buf_2 wire1291 (.A(net848),
    .X(net1291));
 sky130_fd_sc_hd__buf_6 wire1292 (.A(net1293),
    .X(net1292));
 sky130_fd_sc_hd__buf_6 wire1293 (.A(net1294),
    .X(net1293));
 sky130_fd_sc_hd__buf_4 wire1294 (.A(net1295),
    .X(net1294));
 sky130_fd_sc_hd__clkbuf_2 wire1295 (.A(net948),
    .X(net1295));
 sky130_fd_sc_hd__buf_6 wire1296 (.A(net1297),
    .X(net1296));
 sky130_fd_sc_hd__buf_6 wire1297 (.A(net1298),
    .X(net1297));
 sky130_fd_sc_hd__buf_4 wire1298 (.A(net1299),
    .X(net1298));
 sky130_fd_sc_hd__clkbuf_2 wire1299 (.A(net1300),
    .X(net1299));
 sky130_fd_sc_hd__clkbuf_2 wire1300 (.A(net947),
    .X(net1300));
 sky130_fd_sc_hd__buf_4 wire1301 (.A(net1302),
    .X(net1301));
 sky130_fd_sc_hd__buf_6 wire1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_6 wire1303 (.A(net1304),
    .X(net1303));
 sky130_fd_sc_hd__buf_4 wire1304 (.A(net1305),
    .X(net1304));
 sky130_fd_sc_hd__clkbuf_2 wire1305 (.A(net946),
    .X(net1305));
 sky130_fd_sc_hd__buf_6 wire1306 (.A(net1307),
    .X(net1306));
 sky130_fd_sc_hd__buf_6 wire1307 (.A(net1308),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 wire1308 (.A(net1309),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_2 wire1309 (.A(net1310),
    .X(net1309));
 sky130_fd_sc_hd__clkbuf_2 wire1310 (.A(net945),
    .X(net1310));
 sky130_fd_sc_hd__buf_6 wire1311 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_6 wire1312 (.A(net1313),
    .X(net1312));
 sky130_fd_sc_hd__buf_4 wire1313 (.A(net1314),
    .X(net1313));
 sky130_fd_sc_hd__clkbuf_2 wire1314 (.A(net950),
    .X(net1314));
 sky130_fd_sc_hd__buf_6 wire1315 (.A(net1316),
    .X(net1315));
 sky130_fd_sc_hd__buf_6 wire1316 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__buf_4 wire1317 (.A(net1318),
    .X(net1317));
 sky130_fd_sc_hd__clkbuf_2 wire1318 (.A(net949),
    .X(net1318));
 sky130_fd_sc_hd__buf_6 wire1319 (.A(net1320),
    .X(net1319));
 sky130_fd_sc_hd__buf_4 wire1320 (.A(net1321),
    .X(net1320));
 sky130_fd_sc_hd__clkbuf_2 wire1321 (.A(net880),
    .X(net1321));
 sky130_fd_sc_hd__buf_6 wire1322 (.A(net1323),
    .X(net1322));
 sky130_fd_sc_hd__buf_4 wire1323 (.A(net1324),
    .X(net1323));
 sky130_fd_sc_hd__clkbuf_2 wire1324 (.A(net1325),
    .X(net1324));
 sky130_fd_sc_hd__clkbuf_2 wire1325 (.A(net955),
    .X(net1325));
 sky130_fd_sc_hd__buf_4 wire1326 (.A(net1327),
    .X(net1326));
 sky130_fd_sc_hd__buf_4 max_length1327 (.A(wb_in_enable),
    .X(net1327));
 sky130_fd_sc_hd__clkbuf_2 wire1328 (.A(\la_data_in_enable[105] ),
    .X(net1328));
 sky130_fd_sc_hd__clkbuf_2 wire1329 (.A(_0425_),
    .X(net1329));
 sky130_fd_sc_hd__clkbuf_2 wire1330 (.A(_0424_),
    .X(net1330));
 sky130_fd_sc_hd__clkbuf_2 wire1331 (.A(net1332),
    .X(net1331));
 sky130_fd_sc_hd__clkbuf_2 wire1332 (.A(_0423_),
    .X(net1332));
 sky130_fd_sc_hd__clkbuf_2 wire1333 (.A(_0422_),
    .X(net1333));
 sky130_fd_sc_hd__clkbuf_2 wire1334 (.A(_0415_),
    .X(net1334));
 sky130_fd_sc_hd__clkbuf_2 wire1335 (.A(_0406_),
    .X(net1335));
 sky130_fd_sc_hd__clkbuf_2 wire1336 (.A(_0399_),
    .X(net1336));
 sky130_fd_sc_hd__buf_2 wire1337 (.A(net1338),
    .X(net1337));
 sky130_fd_sc_hd__clkbuf_2 wire1338 (.A(_0398_),
    .X(net1338));
 sky130_fd_sc_hd__clkbuf_2 wire1339 (.A(_0396_),
    .X(net1339));
 sky130_fd_sc_hd__buf_2 wire1340 (.A(net1341),
    .X(net1340));
 sky130_fd_sc_hd__clkbuf_2 wire1341 (.A(_0395_),
    .X(net1341));
 sky130_fd_sc_hd__buf_2 wire1342 (.A(net1343),
    .X(net1342));
 sky130_fd_sc_hd__clkbuf_2 wire1343 (.A(_0394_),
    .X(net1343));
 sky130_fd_sc_hd__clkbuf_2 wire1344 (.A(net1345),
    .X(net1344));
 sky130_fd_sc_hd__clkbuf_2 wire1345 (.A(_0393_),
    .X(net1345));
 sky130_fd_sc_hd__buf_2 wire1346 (.A(net1347),
    .X(net1346));
 sky130_fd_sc_hd__clkbuf_2 wire1347 (.A(_0391_),
    .X(net1347));
 sky130_fd_sc_hd__clkbuf_2 wire1348 (.A(_0389_),
    .X(net1348));
 sky130_fd_sc_hd__buf_2 wire1349 (.A(net1350),
    .X(net1349));
 sky130_fd_sc_hd__clkbuf_2 wire1350 (.A(_0388_),
    .X(net1350));
 sky130_fd_sc_hd__clkbuf_2 wire1351 (.A(net1352),
    .X(net1351));
 sky130_fd_sc_hd__clkbuf_2 wire1352 (.A(_0386_),
    .X(net1352));
 sky130_fd_sc_hd__buf_2 wire1353 (.A(net1354),
    .X(net1353));
 sky130_fd_sc_hd__clkbuf_2 wire1354 (.A(_0385_),
    .X(net1354));
 sky130_fd_sc_hd__clkbuf_2 wire1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__clkbuf_2 wire1356 (.A(_0383_),
    .X(net1356));
 sky130_fd_sc_hd__clkbuf_2 wire1357 (.A(_0379_),
    .X(net1357));
 sky130_fd_sc_hd__clkbuf_2 wire1358 (.A(_0377_),
    .X(net1358));
 sky130_fd_sc_hd__clkbuf_2 wire1359 (.A(net1360),
    .X(net1359));
 sky130_fd_sc_hd__clkbuf_2 wire1360 (.A(_0374_),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_2 wire1361 (.A(_0371_),
    .X(net1361));
 sky130_fd_sc_hd__clkbuf_2 wire1362 (.A(_0370_),
    .X(net1362));
 sky130_fd_sc_hd__clkbuf_2 wire1363 (.A(_0369_),
    .X(net1363));
 sky130_fd_sc_hd__clkbuf_2 wire1364 (.A(_0367_),
    .X(net1364));
 sky130_fd_sc_hd__clkbuf_2 wire1365 (.A(_0366_),
    .X(net1365));
 sky130_fd_sc_hd__clkbuf_2 wire1366 (.A(_0365_),
    .X(net1366));
 sky130_fd_sc_hd__clkbuf_2 wire1367 (.A(_0364_),
    .X(net1367));
 sky130_fd_sc_hd__clkbuf_2 wire1368 (.A(_0363_),
    .X(net1368));
 sky130_fd_sc_hd__clkbuf_2 wire1369 (.A(net1370),
    .X(net1369));
 sky130_fd_sc_hd__clkbuf_2 wire1370 (.A(_0361_),
    .X(net1370));
 sky130_fd_sc_hd__clkbuf_2 wire1371 (.A(_0360_),
    .X(net1371));
 sky130_fd_sc_hd__clkbuf_2 wire1372 (.A(net1373),
    .X(net1372));
 sky130_fd_sc_hd__clkbuf_2 wire1373 (.A(_0358_),
    .X(net1373));
 sky130_fd_sc_hd__clkbuf_2 wire1374 (.A(_0357_),
    .X(net1374));
 sky130_fd_sc_hd__clkbuf_2 wire1375 (.A(net1376),
    .X(net1375));
 sky130_fd_sc_hd__clkbuf_2 wire1376 (.A(_0356_),
    .X(net1376));
 sky130_fd_sc_hd__clkbuf_2 wire1377 (.A(_0355_),
    .X(net1377));
 sky130_fd_sc_hd__clkbuf_2 wire1378 (.A(_0354_),
    .X(net1378));
 sky130_fd_sc_hd__clkbuf_2 wire1379 (.A(net1380),
    .X(net1379));
 sky130_fd_sc_hd__clkbuf_2 wire1380 (.A(_0353_),
    .X(net1380));
 sky130_fd_sc_hd__clkbuf_2 wire1381 (.A(_0352_),
    .X(net1381));
 sky130_fd_sc_hd__clkbuf_2 wire1382 (.A(_0351_),
    .X(net1382));
 sky130_fd_sc_hd__clkbuf_2 wire1383 (.A(net1384),
    .X(net1383));
 sky130_fd_sc_hd__clkbuf_2 wire1384 (.A(_0350_),
    .X(net1384));
 sky130_fd_sc_hd__clkbuf_2 wire1385 (.A(_0349_),
    .X(net1385));
 sky130_fd_sc_hd__clkbuf_2 wire1386 (.A(_0348_),
    .X(net1386));
 sky130_fd_sc_hd__clkbuf_2 wire1387 (.A(_0347_),
    .X(net1387));
 sky130_fd_sc_hd__clkbuf_2 wire1388 (.A(net1389),
    .X(net1388));
 sky130_fd_sc_hd__clkbuf_2 wire1389 (.A(_0346_),
    .X(net1389));
 sky130_fd_sc_hd__clkbuf_2 wire1390 (.A(_0345_),
    .X(net1390));
 sky130_fd_sc_hd__clkbuf_2 wire1391 (.A(_0344_),
    .X(net1391));
 sky130_fd_sc_hd__clkbuf_2 wire1392 (.A(_0343_),
    .X(net1392));
 sky130_fd_sc_hd__buf_2 wire1393 (.A(net1394),
    .X(net1393));
 sky130_fd_sc_hd__clkbuf_2 wire1394 (.A(_0342_),
    .X(net1394));
 sky130_fd_sc_hd__clkbuf_2 wire1395 (.A(net1396),
    .X(net1395));
 sky130_fd_sc_hd__clkbuf_2 wire1396 (.A(_0341_),
    .X(net1396));
 sky130_fd_sc_hd__clkbuf_2 wire1397 (.A(net1398),
    .X(net1397));
 sky130_fd_sc_hd__clkbuf_2 wire1398 (.A(_0340_),
    .X(net1398));
 sky130_fd_sc_hd__clkbuf_2 wire1399 (.A(net1400),
    .X(net1399));
 sky130_fd_sc_hd__clkbuf_2 wire1400 (.A(_0339_),
    .X(net1400));
 sky130_fd_sc_hd__clkbuf_2 wire1401 (.A(_0338_),
    .X(net1401));
 sky130_fd_sc_hd__clkbuf_2 wire1402 (.A(_0337_),
    .X(net1402));
 sky130_fd_sc_hd__clkbuf_2 wire1403 (.A(_0336_),
    .X(net1403));
 sky130_fd_sc_hd__clkbuf_2 wire1404 (.A(_0335_),
    .X(net1404));
 sky130_fd_sc_hd__clkbuf_2 wire1405 (.A(_0327_),
    .X(net1405));
 sky130_fd_sc_hd__clkbuf_2 wire1406 (.A(_0324_),
    .X(net1406));
 sky130_fd_sc_hd__clkbuf_2 wire1407 (.A(_0323_),
    .X(net1407));
 sky130_fd_sc_hd__clkbuf_2 wire1408 (.A(_0322_),
    .X(net1408));
 sky130_fd_sc_hd__clkbuf_2 wire1409 (.A(_0320_),
    .X(net1409));
 sky130_fd_sc_hd__clkbuf_2 wire1410 (.A(_0319_),
    .X(net1410));
 sky130_fd_sc_hd__clkbuf_2 wire1411 (.A(_0317_),
    .X(net1411));
 sky130_fd_sc_hd__clkbuf_2 wire1412 (.A(_0315_),
    .X(net1412));
 sky130_fd_sc_hd__clkbuf_2 wire1413 (.A(_0314_),
    .X(net1413));
 sky130_fd_sc_hd__clkbuf_2 wire1414 (.A(_0313_),
    .X(net1414));
 sky130_fd_sc_hd__clkbuf_2 wire1415 (.A(net1416),
    .X(net1415));
 sky130_fd_sc_hd__clkbuf_2 wire1416 (.A(_0312_),
    .X(net1416));
 sky130_fd_sc_hd__buf_2 wire1417 (.A(net1418),
    .X(net1417));
 sky130_fd_sc_hd__clkbuf_2 wire1418 (.A(_0311_),
    .X(net1418));
 sky130_fd_sc_hd__clkbuf_2 wire1419 (.A(net1420),
    .X(net1419));
 sky130_fd_sc_hd__clkbuf_2 wire1420 (.A(_0308_),
    .X(net1420));
 sky130_fd_sc_hd__clkbuf_2 wire1421 (.A(_0307_),
    .X(net1421));
 sky130_fd_sc_hd__clkbuf_2 wire1422 (.A(net1423),
    .X(net1422));
 sky130_fd_sc_hd__clkbuf_2 wire1423 (.A(_0306_),
    .X(net1423));
 sky130_fd_sc_hd__clkbuf_2 wire1424 (.A(net1425),
    .X(net1424));
 sky130_fd_sc_hd__clkbuf_2 wire1425 (.A(_0305_),
    .X(net1425));
 sky130_fd_sc_hd__buf_2 wire1426 (.A(net1427),
    .X(net1426));
 sky130_fd_sc_hd__clkbuf_2 wire1427 (.A(_0302_),
    .X(net1427));
 sky130_fd_sc_hd__buf_2 wire1428 (.A(net1429),
    .X(net1428));
 sky130_fd_sc_hd__clkbuf_2 wire1429 (.A(_0301_),
    .X(net1429));
 sky130_fd_sc_hd__buf_2 wire1430 (.A(net1431),
    .X(net1430));
 sky130_fd_sc_hd__clkbuf_2 wire1431 (.A(_0300_),
    .X(net1431));
 sky130_fd_sc_hd__buf_2 wire1432 (.A(net1433),
    .X(net1432));
 sky130_fd_sc_hd__clkbuf_2 wire1433 (.A(net1434),
    .X(net1433));
 sky130_fd_sc_hd__clkbuf_2 wire1434 (.A(_0299_),
    .X(net1434));
 sky130_fd_sc_hd__buf_2 wire1435 (.A(net1436),
    .X(net1435));
 sky130_fd_sc_hd__clkbuf_2 wire1436 (.A(net1437),
    .X(net1436));
 sky130_fd_sc_hd__clkbuf_2 wire1437 (.A(_0298_),
    .X(net1437));
 sky130_fd_sc_hd__buf_2 wire1438 (.A(net1439),
    .X(net1438));
 sky130_fd_sc_hd__clkbuf_2 wire1439 (.A(_0297_),
    .X(net1439));
 sky130_fd_sc_hd__clkbuf_2 wire1440 (.A(net1441),
    .X(net1440));
 sky130_fd_sc_hd__clkbuf_2 wire1441 (.A(_0296_),
    .X(net1441));
 sky130_fd_sc_hd__clkbuf_2 wire1442 (.A(_0295_),
    .X(net1442));
 sky130_fd_sc_hd__clkbuf_2 wire1443 (.A(_0282_),
    .X(net1443));
 sky130_fd_sc_hd__clkbuf_2 wire1444 (.A(_0271_),
    .X(net1444));
 sky130_fd_sc_hd__clkbuf_2 wire1445 (.A(_0270_),
    .X(net1445));
 sky130_fd_sc_hd__clkbuf_2 wire1446 (.A(_0269_),
    .X(net1446));
 sky130_fd_sc_hd__buf_2 wire1447 (.A(net1448),
    .X(net1447));
 sky130_fd_sc_hd__clkbuf_2 wire1448 (.A(_0268_),
    .X(net1448));
 sky130_fd_sc_hd__buf_2 wire1449 (.A(net1450),
    .X(net1449));
 sky130_fd_sc_hd__clkbuf_2 wire1450 (.A(_0267_),
    .X(net1450));
 sky130_fd_sc_hd__buf_2 wire1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__clkbuf_2 wire1452 (.A(_0266_),
    .X(net1452));
 sky130_fd_sc_hd__buf_2 wire1453 (.A(net1454),
    .X(net1453));
 sky130_fd_sc_hd__clkbuf_2 wire1454 (.A(net1455),
    .X(net1454));
 sky130_fd_sc_hd__clkbuf_2 wire1455 (.A(_0265_),
    .X(net1455));
 sky130_fd_sc_hd__buf_2 wire1456 (.A(net1457),
    .X(net1456));
 sky130_fd_sc_hd__clkbuf_2 wire1457 (.A(_0264_),
    .X(net1457));
 sky130_fd_sc_hd__buf_4 wire1458 (.A(net1459),
    .X(net1458));
 sky130_fd_sc_hd__clkbuf_2 wire1459 (.A(_0263_),
    .X(net1459));
 sky130_fd_sc_hd__clkbuf_2 wire1460 (.A(net1461),
    .X(net1460));
 sky130_fd_sc_hd__clkbuf_2 wire1461 (.A(_0262_),
    .X(net1461));
 sky130_fd_sc_hd__clkbuf_2 wire1462 (.A(net1463),
    .X(net1462));
 sky130_fd_sc_hd__clkbuf_2 wire1463 (.A(_0261_),
    .X(net1463));
 sky130_fd_sc_hd__buf_2 wire1464 (.A(net1465),
    .X(net1464));
 sky130_fd_sc_hd__clkbuf_2 wire1465 (.A(_0260_),
    .X(net1465));
 sky130_fd_sc_hd__buf_2 wire1466 (.A(net1467),
    .X(net1466));
 sky130_fd_sc_hd__clkbuf_2 wire1467 (.A(net1468),
    .X(net1467));
 sky130_fd_sc_hd__clkbuf_2 wire1468 (.A(_0259_),
    .X(net1468));
 sky130_fd_sc_hd__buf_2 wire1469 (.A(net1470),
    .X(net1469));
 sky130_fd_sc_hd__clkbuf_2 wire1470 (.A(_0258_),
    .X(net1470));
 sky130_fd_sc_hd__buf_2 wire1471 (.A(net1472),
    .X(net1471));
 sky130_fd_sc_hd__clkbuf_2 wire1472 (.A(_0257_),
    .X(net1472));
 sky130_fd_sc_hd__clkbuf_2 wire1473 (.A(net1474),
    .X(net1473));
 sky130_fd_sc_hd__clkbuf_2 wire1474 (.A(_0256_),
    .X(net1474));
 sky130_fd_sc_hd__clkbuf_2 wire1475 (.A(_0255_),
    .X(net1475));
 sky130_fd_sc_hd__clkbuf_2 wire1476 (.A(_0254_),
    .X(net1476));
 sky130_fd_sc_hd__clkbuf_2 wire1477 (.A(_0252_),
    .X(net1477));
 sky130_fd_sc_hd__clkbuf_2 wire1478 (.A(_0251_),
    .X(net1478));
 sky130_fd_sc_hd__clkbuf_2 wire1479 (.A(_0249_),
    .X(net1479));
 sky130_fd_sc_hd__clkbuf_2 wire1480 (.A(net1481),
    .X(net1480));
 sky130_fd_sc_hd__clkbuf_2 wire1481 (.A(_0248_),
    .X(net1481));
 sky130_fd_sc_hd__clkbuf_2 wire1482 (.A(_0247_),
    .X(net1482));
 sky130_fd_sc_hd__buf_2 wire1483 (.A(net1484),
    .X(net1483));
 sky130_fd_sc_hd__clkbuf_2 wire1484 (.A(_0246_),
    .X(net1484));
 sky130_fd_sc_hd__clkbuf_2 wire1485 (.A(_0244_),
    .X(net1485));
 sky130_fd_sc_hd__clkbuf_2 wire1486 (.A(_0243_),
    .X(net1486));
 sky130_fd_sc_hd__clkbuf_2 wire1487 (.A(_0241_),
    .X(net1487));
 sky130_fd_sc_hd__clkbuf_2 wire1488 (.A(_0234_),
    .X(net1488));
 sky130_fd_sc_hd__clkbuf_2 wire1489 (.A(_0230_),
    .X(net1489));
 sky130_fd_sc_hd__clkbuf_2 wire1490 (.A(_0229_),
    .X(net1490));
 sky130_fd_sc_hd__clkbuf_2 wire1491 (.A(_0228_),
    .X(net1491));
 sky130_fd_sc_hd__clkbuf_2 wire1492 (.A(_0227_),
    .X(net1492));
 sky130_fd_sc_hd__clkbuf_2 wire1493 (.A(net1494),
    .X(net1493));
 sky130_fd_sc_hd__clkbuf_2 wire1494 (.A(_0226_),
    .X(net1494));
 sky130_fd_sc_hd__clkbuf_2 wire1495 (.A(_0225_),
    .X(net1495));
 sky130_fd_sc_hd__buf_2 wire1496 (.A(net1497),
    .X(net1496));
 sky130_fd_sc_hd__clkbuf_2 wire1497 (.A(_0223_),
    .X(net1497));
 sky130_fd_sc_hd__clkbuf_2 wire1498 (.A(_0222_),
    .X(net1498));
 sky130_fd_sc_hd__buf_2 wire1499 (.A(net1500),
    .X(net1499));
 sky130_fd_sc_hd__clkbuf_2 wire1500 (.A(_0220_),
    .X(net1500));
 sky130_fd_sc_hd__clkbuf_2 wire1501 (.A(_0219_),
    .X(net1501));
 sky130_fd_sc_hd__clkbuf_2 wire1502 (.A(_0218_),
    .X(net1502));
 sky130_fd_sc_hd__clkbuf_2 wire1503 (.A(net1504),
    .X(net1503));
 sky130_fd_sc_hd__clkbuf_2 wire1504 (.A(_0216_),
    .X(net1504));
 sky130_fd_sc_hd__clkbuf_2 wire1505 (.A(_0215_),
    .X(net1505));
 sky130_fd_sc_hd__clkbuf_2 wire1506 (.A(_0214_),
    .X(net1506));
 sky130_fd_sc_hd__clkbuf_2 wire1507 (.A(_0213_),
    .X(net1507));
 sky130_fd_sc_hd__clkbuf_2 wire1508 (.A(_0212_),
    .X(net1508));
 sky130_fd_sc_hd__clkbuf_2 wire1509 (.A(_0204_),
    .X(net1509));
 sky130_fd_sc_hd__clkbuf_2 wire1510 (.A(_0203_),
    .X(net1510));
 sky130_fd_sc_hd__clkbuf_2 wire1511 (.A(_0202_),
    .X(net1511));
 sky130_fd_sc_hd__clkbuf_2 wire1512 (.A(_0201_),
    .X(net1512));
 sky130_fd_sc_hd__buf_6 wire1513 (.A(net1514),
    .X(net1513));
 sky130_fd_sc_hd__buf_4 wire1514 (.A(net1515),
    .X(net1514));
 sky130_fd_sc_hd__clkbuf_2 wire1515 (.A(_0200_),
    .X(net1515));
 sky130_fd_sc_hd__buf_4 wire1516 (.A(net1517),
    .X(net1516));
 sky130_fd_sc_hd__clkbuf_2 wire1517 (.A(_0199_),
    .X(net1517));
 sky130_fd_sc_hd__buf_4 wire1518 (.A(net1519),
    .X(net1518));
 sky130_fd_sc_hd__clkbuf_2 wire1519 (.A(_0198_),
    .X(net1519));
 sky130_fd_sc_hd__buf_4 wire1520 (.A(net1521),
    .X(net1520));
 sky130_fd_sc_hd__clkbuf_2 wire1521 (.A(_0197_),
    .X(net1521));
 sky130_fd_sc_hd__clkbuf_2 wire1522 (.A(_0196_),
    .X(net1522));
 sky130_fd_sc_hd__clkbuf_2 wire1523 (.A(_0195_),
    .X(net1523));
 sky130_fd_sc_hd__clkbuf_2 wire1524 (.A(_0194_),
    .X(net1524));
 sky130_fd_sc_hd__clkbuf_2 wire1525 (.A(_0193_),
    .X(net1525));
 sky130_fd_sc_hd__clkbuf_2 wire1526 (.A(net1527),
    .X(net1526));
 sky130_fd_sc_hd__clkbuf_2 wire1527 (.A(_0192_),
    .X(net1527));
 sky130_fd_sc_hd__clkbuf_2 wire1528 (.A(net1529),
    .X(net1528));
 sky130_fd_sc_hd__clkbuf_2 wire1529 (.A(_0191_),
    .X(net1529));
 sky130_fd_sc_hd__clkbuf_2 wire1530 (.A(_0190_),
    .X(net1530));
 sky130_fd_sc_hd__clkbuf_2 wire1531 (.A(_0188_),
    .X(net1531));
 sky130_fd_sc_hd__clkbuf_2 wire1532 (.A(_0187_),
    .X(net1532));
 sky130_fd_sc_hd__clkbuf_2 wire1533 (.A(net1534),
    .X(net1533));
 sky130_fd_sc_hd__clkbuf_2 wire1534 (.A(_0186_),
    .X(net1534));
 sky130_fd_sc_hd__clkbuf_2 wire1535 (.A(_0185_),
    .X(net1535));
 sky130_fd_sc_hd__clkbuf_2 wire1536 (.A(_0184_),
    .X(net1536));
 sky130_fd_sc_hd__clkbuf_2 wire1537 (.A(_0183_),
    .X(net1537));
 sky130_fd_sc_hd__clkbuf_2 wire1538 (.A(_0182_),
    .X(net1538));
 sky130_fd_sc_hd__clkbuf_2 wire1539 (.A(_0180_),
    .X(net1539));
 sky130_fd_sc_hd__clkbuf_2 wire1540 (.A(_0175_),
    .X(net1540));
 sky130_fd_sc_hd__clkbuf_2 wire1541 (.A(_0149_),
    .X(net1541));
 sky130_fd_sc_hd__clkbuf_2 wire1542 (.A(_0148_),
    .X(net1542));
 sky130_fd_sc_hd__buf_4 wire1543 (.A(net1544),
    .X(net1543));
 sky130_fd_sc_hd__clkbuf_2 wire1544 (.A(net1545),
    .X(net1544));
 sky130_fd_sc_hd__clkbuf_2 wire1545 (.A(_0140_),
    .X(net1545));
 sky130_fd_sc_hd__clkbuf_2 wire1546 (.A(net1547),
    .X(net1546));
 sky130_fd_sc_hd__clkbuf_2 wire1547 (.A(_0139_),
    .X(net1547));
 sky130_fd_sc_hd__clkbuf_2 wire1548 (.A(_0138_),
    .X(net1548));
 sky130_fd_sc_hd__clkbuf_2 wire1549 (.A(_0137_),
    .X(net1549));
 sky130_fd_sc_hd__clkbuf_2 wire1550 (.A(_0136_),
    .X(net1550));
 sky130_fd_sc_hd__clkbuf_2 wire1551 (.A(_0135_),
    .X(net1551));
 sky130_fd_sc_hd__clkbuf_2 wire1552 (.A(_0115_),
    .X(net1552));
 sky130_fd_sc_hd__clkbuf_2 wire1553 (.A(_0113_),
    .X(net1553));
 sky130_fd_sc_hd__clkbuf_2 wire1554 (.A(_0107_),
    .X(net1554));
 sky130_fd_sc_hd__clkbuf_2 wire1555 (.A(_0105_),
    .X(net1555));
 sky130_fd_sc_hd__clkbuf_2 wire1556 (.A(net1557),
    .X(net1556));
 sky130_fd_sc_hd__clkbuf_2 wire1557 (.A(_0104_),
    .X(net1557));
 sky130_fd_sc_hd__buf_6 wire1558 (.A(net1559),
    .X(net1558));
 sky130_fd_sc_hd__buf_4 wire1559 (.A(net1560),
    .X(net1559));
 sky130_fd_sc_hd__clkbuf_2 wire1560 (.A(_0103_),
    .X(net1560));
 sky130_fd_sc_hd__buf_6 wire1561 (.A(net1562),
    .X(net1561));
 sky130_fd_sc_hd__buf_4 wire1562 (.A(net1563),
    .X(net1562));
 sky130_fd_sc_hd__clkbuf_2 wire1563 (.A(_0102_),
    .X(net1563));
 sky130_fd_sc_hd__buf_2 wire1564 (.A(net1565),
    .X(net1564));
 sky130_fd_sc_hd__clkbuf_2 wire1565 (.A(net1566),
    .X(net1565));
 sky130_fd_sc_hd__clkbuf_2 wire1566 (.A(_0101_),
    .X(net1566));
 sky130_fd_sc_hd__buf_6 wire1567 (.A(net1568),
    .X(net1567));
 sky130_fd_sc_hd__buf_4 wire1568 (.A(net1569),
    .X(net1568));
 sky130_fd_sc_hd__clkbuf_2 wire1569 (.A(_0100_),
    .X(net1569));
 sky130_fd_sc_hd__clkbuf_2 wire1570 (.A(net1571),
    .X(net1570));
 sky130_fd_sc_hd__clkbuf_2 wire1571 (.A(_0099_),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 wire1572 (.A(net1573),
    .X(net1572));
 sky130_fd_sc_hd__clkbuf_2 wire1573 (.A(net1574),
    .X(net1573));
 sky130_fd_sc_hd__clkbuf_2 wire1574 (.A(_0098_),
    .X(net1574));
 sky130_fd_sc_hd__buf_4 wire1575 (.A(net1576),
    .X(net1575));
 sky130_fd_sc_hd__clkbuf_2 wire1576 (.A(_0097_),
    .X(net1576));
 sky130_fd_sc_hd__buf_4 wire1577 (.A(net1578),
    .X(net1577));
 sky130_fd_sc_hd__clkbuf_2 wire1578 (.A(net1579),
    .X(net1578));
 sky130_fd_sc_hd__clkbuf_2 wire1579 (.A(_0096_),
    .X(net1579));
 sky130_fd_sc_hd__buf_2 wire1580 (.A(net1581),
    .X(net1580));
 sky130_fd_sc_hd__clkbuf_2 wire1581 (.A(_0095_),
    .X(net1581));
 sky130_fd_sc_hd__buf_4 wire1582 (.A(net1583),
    .X(net1582));
 sky130_fd_sc_hd__clkbuf_2 wire1583 (.A(net1584),
    .X(net1583));
 sky130_fd_sc_hd__clkbuf_2 wire1584 (.A(_0094_),
    .X(net1584));
 sky130_fd_sc_hd__buf_4 wire1585 (.A(net1586),
    .X(net1585));
 sky130_fd_sc_hd__clkbuf_2 wire1586 (.A(net1587),
    .X(net1586));
 sky130_fd_sc_hd__clkbuf_2 wire1587 (.A(_0093_),
    .X(net1587));
 sky130_fd_sc_hd__buf_6 wire1588 (.A(net1589),
    .X(net1588));
 sky130_fd_sc_hd__buf_4 wire1589 (.A(net1590),
    .X(net1589));
 sky130_fd_sc_hd__clkbuf_2 wire1590 (.A(_0092_),
    .X(net1590));
 sky130_fd_sc_hd__buf_4 wire1591 (.A(net1592),
    .X(net1591));
 sky130_fd_sc_hd__buf_4 wire1592 (.A(net1593),
    .X(net1592));
 sky130_fd_sc_hd__clkbuf_2 wire1593 (.A(_0091_),
    .X(net1593));
 sky130_fd_sc_hd__buf_4 wire1594 (.A(net1595),
    .X(net1594));
 sky130_fd_sc_hd__clkbuf_2 wire1595 (.A(net1596),
    .X(net1595));
 sky130_fd_sc_hd__clkbuf_2 wire1596 (.A(_0090_),
    .X(net1596));
 sky130_fd_sc_hd__buf_6 wire1597 (.A(net1598),
    .X(net1597));
 sky130_fd_sc_hd__buf_4 wire1598 (.A(net1599),
    .X(net1598));
 sky130_fd_sc_hd__clkbuf_2 wire1599 (.A(_0089_),
    .X(net1599));
 sky130_fd_sc_hd__buf_2 wire1600 (.A(net1601),
    .X(net1600));
 sky130_fd_sc_hd__clkbuf_2 wire1601 (.A(_0088_),
    .X(net1601));
 sky130_fd_sc_hd__buf_4 wire1602 (.A(net1603),
    .X(net1602));
 sky130_fd_sc_hd__buf_4 wire1603 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__clkbuf_2 wire1604 (.A(_0087_),
    .X(net1604));
 sky130_fd_sc_hd__buf_4 wire1605 (.A(net1606),
    .X(net1605));
 sky130_fd_sc_hd__clkbuf_2 wire1606 (.A(_0085_),
    .X(net1606));
 sky130_fd_sc_hd__clkbuf_2 wire1607 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__clkbuf_2 wire1608 (.A(_0084_),
    .X(net1608));
 sky130_fd_sc_hd__buf_4 wire1609 (.A(net1610),
    .X(net1609));
 sky130_fd_sc_hd__buf_4 wire1610 (.A(net1611),
    .X(net1610));
 sky130_fd_sc_hd__buf_2 wire1611 (.A(_0083_),
    .X(net1611));
 sky130_fd_sc_hd__buf_2 wire1612 (.A(net1613),
    .X(net1612));
 sky130_fd_sc_hd__clkbuf_2 wire1613 (.A(net1614),
    .X(net1613));
 sky130_fd_sc_hd__clkbuf_2 wire1614 (.A(_0082_),
    .X(net1614));
 sky130_fd_sc_hd__buf_4 wire1615 (.A(net1616),
    .X(net1615));
 sky130_fd_sc_hd__clkbuf_2 wire1616 (.A(_0081_),
    .X(net1616));
 sky130_fd_sc_hd__buf_6 wire1617 (.A(net1618),
    .X(net1617));
 sky130_fd_sc_hd__buf_4 wire1618 (.A(net1619),
    .X(net1618));
 sky130_fd_sc_hd__clkbuf_2 wire1619 (.A(_0080_),
    .X(net1619));
 sky130_fd_sc_hd__buf_2 wire1620 (.A(_0079_),
    .X(net1620));
 sky130_fd_sc_hd__clkbuf_2 wire1621 (.A(net1622),
    .X(net1621));
 sky130_fd_sc_hd__clkbuf_2 wire1622 (.A(_0078_),
    .X(net1622));
 sky130_fd_sc_hd__clkbuf_2 wire1623 (.A(net1624),
    .X(net1623));
 sky130_fd_sc_hd__clkbuf_2 wire1624 (.A(_0077_),
    .X(net1624));
 sky130_fd_sc_hd__buf_4 wire1625 (.A(net1626),
    .X(net1625));
 sky130_fd_sc_hd__clkbuf_4 wire1626 (.A(_0076_),
    .X(net1626));
 sky130_fd_sc_hd__buf_2 wire1627 (.A(net1628),
    .X(net1627));
 sky130_fd_sc_hd__buf_4 wire1628 (.A(_0075_),
    .X(net1628));
 sky130_fd_sc_hd__clkbuf_2 wire1629 (.A(_0074_),
    .X(net1629));
 sky130_fd_sc_hd__clkbuf_2 wire1630 (.A(_0071_),
    .X(net1630));
 sky130_fd_sc_hd__clkbuf_2 wire1631 (.A(_0036_),
    .X(net1631));
 sky130_fd_sc_hd__clkbuf_2 wire1632 (.A(_0031_),
    .X(net1632));
 sky130_fd_sc_hd__clkbuf_2 wire1633 (.A(net99),
    .X(net1633));
 sky130_fd_sc_hd__clkbuf_2 wire1634 (.A(net96),
    .X(net1634));
 sky130_fd_sc_hd__clkbuf_2 wire1635 (.A(net95),
    .X(net1635));
 sky130_fd_sc_hd__clkbuf_2 wire1636 (.A(net91),
    .X(net1636));
 sky130_fd_sc_hd__clkbuf_2 wire1637 (.A(net90),
    .X(net1637));
 sky130_fd_sc_hd__clkbuf_2 wire1638 (.A(net89),
    .X(net1638));
 sky130_fd_sc_hd__clkbuf_2 wire1639 (.A(net88),
    .X(net1639));
 sky130_fd_sc_hd__clkbuf_2 wire1640 (.A(net85),
    .X(net1640));
 sky130_fd_sc_hd__clkbuf_2 wire1641 (.A(net82),
    .X(net1641));
 sky130_fd_sc_hd__clkbuf_2 wire1642 (.A(net81),
    .X(net1642));
 sky130_fd_sc_hd__clkbuf_2 wire1643 (.A(net80),
    .X(net1643));
 sky130_fd_sc_hd__clkbuf_2 wire1644 (.A(net79),
    .X(net1644));
 sky130_fd_sc_hd__clkbuf_2 wire1645 (.A(net69),
    .X(net1645));
 sky130_fd_sc_hd__clkbuf_2 wire1646 (.A(net67),
    .X(net1646));
 sky130_fd_sc_hd__clkbuf_2 wire1647 (.A(net53),
    .X(net1647));
 sky130_fd_sc_hd__clkbuf_2 wire1648 (.A(net51),
    .X(net1648));
 sky130_fd_sc_hd__clkbuf_2 wire1649 (.A(net459),
    .X(net1649));
 sky130_fd_sc_hd__clkbuf_2 wire1650 (.A(net458),
    .X(net1650));
 sky130_fd_sc_hd__clkbuf_2 wire1651 (.A(net452),
    .X(net1651));
 sky130_fd_sc_hd__clkbuf_2 wire1652 (.A(net1653),
    .X(net1652));
 sky130_fd_sc_hd__clkbuf_2 wire1653 (.A(net451),
    .X(net1653));
 sky130_fd_sc_hd__clkbuf_2 wire1654 (.A(net1655),
    .X(net1654));
 sky130_fd_sc_hd__clkbuf_2 wire1655 (.A(net450),
    .X(net1655));
 sky130_fd_sc_hd__buf_2 wire1656 (.A(net1657),
    .X(net1656));
 sky130_fd_sc_hd__clkbuf_2 wire1657 (.A(net449),
    .X(net1657));
 sky130_fd_sc_hd__buf_2 wire1658 (.A(net1659),
    .X(net1658));
 sky130_fd_sc_hd__clkbuf_2 wire1659 (.A(net448),
    .X(net1659));
 sky130_fd_sc_hd__buf_2 wire1660 (.A(net1661),
    .X(net1660));
 sky130_fd_sc_hd__clkbuf_2 wire1661 (.A(net447),
    .X(net1661));
 sky130_fd_sc_hd__buf_2 wire1662 (.A(net1663),
    .X(net1662));
 sky130_fd_sc_hd__clkbuf_2 wire1663 (.A(net1664),
    .X(net1663));
 sky130_fd_sc_hd__clkbuf_2 wire1664 (.A(net446),
    .X(net1664));
 sky130_fd_sc_hd__clkbuf_2 wire1665 (.A(net1666),
    .X(net1665));
 sky130_fd_sc_hd__clkbuf_2 wire1666 (.A(net445),
    .X(net1666));
 sky130_fd_sc_hd__clkbuf_2 wire1667 (.A(net1668),
    .X(net1667));
 sky130_fd_sc_hd__clkbuf_2 wire1668 (.A(net444),
    .X(net1668));
 sky130_fd_sc_hd__clkbuf_2 wire1669 (.A(net443),
    .X(net1669));
 sky130_fd_sc_hd__clkbuf_2 wire1670 (.A(net442),
    .X(net1670));
 sky130_fd_sc_hd__clkbuf_2 wire1671 (.A(net441),
    .X(net1671));
 sky130_fd_sc_hd__clkbuf_2 wire1672 (.A(net44),
    .X(net1672));
 sky130_fd_sc_hd__clkbuf_2 wire1673 (.A(net436),
    .X(net1673));
 sky130_fd_sc_hd__clkbuf_2 wire1674 (.A(net1675),
    .X(net1674));
 sky130_fd_sc_hd__clkbuf_2 wire1675 (.A(net435),
    .X(net1675));
 sky130_fd_sc_hd__clkbuf_2 wire1676 (.A(net1677),
    .X(net1676));
 sky130_fd_sc_hd__clkbuf_2 wire1677 (.A(net434),
    .X(net1677));
 sky130_fd_sc_hd__clkbuf_2 wire1678 (.A(net433),
    .X(net1678));
 sky130_fd_sc_hd__buf_2 wire1679 (.A(net1680),
    .X(net1679));
 sky130_fd_sc_hd__clkbuf_2 wire1680 (.A(net1681),
    .X(net1680));
 sky130_fd_sc_hd__clkbuf_2 wire1681 (.A(net432),
    .X(net1681));
 sky130_fd_sc_hd__clkbuf_2 wire1682 (.A(net431),
    .X(net1682));
 sky130_fd_sc_hd__clkbuf_2 wire1683 (.A(net430),
    .X(net1683));
 sky130_fd_sc_hd__clkbuf_2 wire1684 (.A(net429),
    .X(net1684));
 sky130_fd_sc_hd__clkbuf_2 wire1685 (.A(net1686),
    .X(net1685));
 sky130_fd_sc_hd__clkbuf_2 wire1686 (.A(net428),
    .X(net1686));
 sky130_fd_sc_hd__buf_2 wire1687 (.A(net1688),
    .X(net1687));
 sky130_fd_sc_hd__clkbuf_2 wire1688 (.A(net427),
    .X(net1688));
 sky130_fd_sc_hd__clkbuf_2 wire1689 (.A(net1690),
    .X(net1689));
 sky130_fd_sc_hd__clkbuf_2 wire1690 (.A(net426),
    .X(net1690));
 sky130_fd_sc_hd__clkbuf_2 wire1691 (.A(net424),
    .X(net1691));
 sky130_fd_sc_hd__clkbuf_2 wire1692 (.A(net423),
    .X(net1692));
 sky130_fd_sc_hd__clkbuf_2 wire1693 (.A(net422),
    .X(net1693));
 sky130_fd_sc_hd__buf_2 wire1694 (.A(net1695),
    .X(net1694));
 sky130_fd_sc_hd__clkbuf_2 wire1695 (.A(net1696),
    .X(net1695));
 sky130_fd_sc_hd__clkbuf_2 wire1696 (.A(net421),
    .X(net1696));
 sky130_fd_sc_hd__buf_4 wire1697 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__clkbuf_2 wire1698 (.A(net1699),
    .X(net1698));
 sky130_fd_sc_hd__clkbuf_2 wire1699 (.A(net420),
    .X(net1699));
 sky130_fd_sc_hd__buf_2 wire1700 (.A(net1701),
    .X(net1700));
 sky130_fd_sc_hd__clkbuf_2 wire1701 (.A(net1702),
    .X(net1701));
 sky130_fd_sc_hd__clkbuf_2 wire1702 (.A(net419),
    .X(net1702));
 sky130_fd_sc_hd__buf_6 wire1703 (.A(net1704),
    .X(net1703));
 sky130_fd_sc_hd__buf_6 wire1704 (.A(net1705),
    .X(net1704));
 sky130_fd_sc_hd__buf_4 wire1705 (.A(net1706),
    .X(net1705));
 sky130_fd_sc_hd__clkbuf_2 wire1706 (.A(net1707),
    .X(net1706));
 sky130_fd_sc_hd__clkbuf_2 wire1707 (.A(net418),
    .X(net1707));
 sky130_fd_sc_hd__buf_6 wire1708 (.A(net1709),
    .X(net1708));
 sky130_fd_sc_hd__buf_6 wire1709 (.A(net1710),
    .X(net1709));
 sky130_fd_sc_hd__buf_6 wire1710 (.A(net1711),
    .X(net1710));
 sky130_fd_sc_hd__buf_4 wire1711 (.A(net1712),
    .X(net1711));
 sky130_fd_sc_hd__clkbuf_2 wire1712 (.A(net1713),
    .X(net1712));
 sky130_fd_sc_hd__clkbuf_2 wire1713 (.A(net417),
    .X(net1713));
 sky130_fd_sc_hd__buf_6 wire1714 (.A(net1715),
    .X(net1714));
 sky130_fd_sc_hd__buf_4 wire1715 (.A(net1716),
    .X(net1715));
 sky130_fd_sc_hd__clkbuf_2 wire1716 (.A(net416),
    .X(net1716));
 sky130_fd_sc_hd__buf_6 wire1717 (.A(net1718),
    .X(net1717));
 sky130_fd_sc_hd__buf_6 wire1718 (.A(net1719),
    .X(net1718));
 sky130_fd_sc_hd__buf_4 wire1719 (.A(net1720),
    .X(net1719));
 sky130_fd_sc_hd__clkbuf_2 wire1720 (.A(net415),
    .X(net1720));
 sky130_fd_sc_hd__buf_6 wire1721 (.A(net1722),
    .X(net1721));
 sky130_fd_sc_hd__buf_6 wire1722 (.A(net1723),
    .X(net1722));
 sky130_fd_sc_hd__buf_6 wire1723 (.A(net1724),
    .X(net1723));
 sky130_fd_sc_hd__buf_4 wire1724 (.A(net1725),
    .X(net1724));
 sky130_fd_sc_hd__clkbuf_2 wire1725 (.A(net414),
    .X(net1725));
 sky130_fd_sc_hd__buf_6 wire1726 (.A(net1727),
    .X(net1726));
 sky130_fd_sc_hd__buf_6 wire1727 (.A(net1728),
    .X(net1727));
 sky130_fd_sc_hd__buf_4 wire1728 (.A(net1729),
    .X(net1728));
 sky130_fd_sc_hd__clkbuf_2 wire1729 (.A(net413),
    .X(net1729));
 sky130_fd_sc_hd__buf_6 wire1730 (.A(net1731),
    .X(net1730));
 sky130_fd_sc_hd__buf_6 wire1731 (.A(net1732),
    .X(net1731));
 sky130_fd_sc_hd__buf_4 wire1732 (.A(net1733),
    .X(net1732));
 sky130_fd_sc_hd__clkbuf_2 wire1733 (.A(net412),
    .X(net1733));
 sky130_fd_sc_hd__buf_6 wire1734 (.A(net1735),
    .X(net1734));
 sky130_fd_sc_hd__buf_6 wire1735 (.A(net1736),
    .X(net1735));
 sky130_fd_sc_hd__buf_4 wire1736 (.A(net1737),
    .X(net1736));
 sky130_fd_sc_hd__clkbuf_2 wire1737 (.A(net411),
    .X(net1737));
 sky130_fd_sc_hd__buf_4 wire1738 (.A(net1739),
    .X(net1738));
 sky130_fd_sc_hd__buf_6 wire1739 (.A(net1740),
    .X(net1739));
 sky130_fd_sc_hd__buf_6 wire1740 (.A(net1741),
    .X(net1740));
 sky130_fd_sc_hd__buf_4 wire1741 (.A(net1742),
    .X(net1741));
 sky130_fd_sc_hd__clkbuf_2 wire1742 (.A(net410),
    .X(net1742));
 sky130_fd_sc_hd__clkbuf_2 wire1743 (.A(net41),
    .X(net1743));
 sky130_fd_sc_hd__buf_6 wire1744 (.A(net1745),
    .X(net1744));
 sky130_fd_sc_hd__buf_6 wire1745 (.A(net1746),
    .X(net1745));
 sky130_fd_sc_hd__buf_4 wire1746 (.A(net1747),
    .X(net1746));
 sky130_fd_sc_hd__clkbuf_2 wire1747 (.A(net409),
    .X(net1747));
 sky130_fd_sc_hd__buf_6 wire1748 (.A(net1749),
    .X(net1748));
 sky130_fd_sc_hd__buf_6 wire1749 (.A(net1750),
    .X(net1749));
 sky130_fd_sc_hd__buf_4 wire1750 (.A(net1751),
    .X(net1750));
 sky130_fd_sc_hd__clkbuf_2 wire1751 (.A(net408),
    .X(net1751));
 sky130_fd_sc_hd__buf_6 wire1752 (.A(net1753),
    .X(net1752));
 sky130_fd_sc_hd__buf_6 wire1753 (.A(net1754),
    .X(net1753));
 sky130_fd_sc_hd__buf_4 wire1754 (.A(net1755),
    .X(net1754));
 sky130_fd_sc_hd__clkbuf_2 wire1755 (.A(net1756),
    .X(net1755));
 sky130_fd_sc_hd__clkbuf_2 wire1756 (.A(net407),
    .X(net1756));
 sky130_fd_sc_hd__buf_6 wire1757 (.A(net1758),
    .X(net1757));
 sky130_fd_sc_hd__buf_6 wire1758 (.A(net1759),
    .X(net1758));
 sky130_fd_sc_hd__buf_4 wire1759 (.A(net1760),
    .X(net1759));
 sky130_fd_sc_hd__clkbuf_2 wire1760 (.A(net406),
    .X(net1760));
 sky130_fd_sc_hd__buf_6 wire1761 (.A(net1762),
    .X(net1761));
 sky130_fd_sc_hd__buf_6 wire1762 (.A(net1763),
    .X(net1762));
 sky130_fd_sc_hd__buf_6 wire1763 (.A(net1764),
    .X(net1763));
 sky130_fd_sc_hd__buf_4 wire1764 (.A(net1765),
    .X(net1764));
 sky130_fd_sc_hd__clkbuf_2 wire1765 (.A(net405),
    .X(net1765));
 sky130_fd_sc_hd__buf_6 wire1766 (.A(net1767),
    .X(net1766));
 sky130_fd_sc_hd__buf_6 wire1767 (.A(net1768),
    .X(net1767));
 sky130_fd_sc_hd__buf_4 wire1768 (.A(net1769),
    .X(net1768));
 sky130_fd_sc_hd__clkbuf_2 wire1769 (.A(net1770),
    .X(net1769));
 sky130_fd_sc_hd__clkbuf_2 wire1770 (.A(net404),
    .X(net1770));
 sky130_fd_sc_hd__buf_6 wire1771 (.A(net1772),
    .X(net1771));
 sky130_fd_sc_hd__buf_6 wire1772 (.A(net1773),
    .X(net1772));
 sky130_fd_sc_hd__buf_4 wire1773 (.A(net1774),
    .X(net1773));
 sky130_fd_sc_hd__clkbuf_2 wire1774 (.A(net403),
    .X(net1774));
 sky130_fd_sc_hd__buf_2 wire1775 (.A(net1776),
    .X(net1775));
 sky130_fd_sc_hd__clkbuf_2 wire1776 (.A(net1777),
    .X(net1776));
 sky130_fd_sc_hd__clkbuf_2 wire1777 (.A(net402),
    .X(net1777));
 sky130_fd_sc_hd__buf_4 wire1778 (.A(net1779),
    .X(net1778));
 sky130_fd_sc_hd__buf_6 wire1779 (.A(net1780),
    .X(net1779));
 sky130_fd_sc_hd__buf_6 wire1780 (.A(net1781),
    .X(net1780));
 sky130_fd_sc_hd__buf_4 wire1781 (.A(net1782),
    .X(net1781));
 sky130_fd_sc_hd__clkbuf_2 wire1782 (.A(net401),
    .X(net1782));
 sky130_fd_sc_hd__buf_6 wire1783 (.A(net1784),
    .X(net1783));
 sky130_fd_sc_hd__buf_4 wire1784 (.A(net1785),
    .X(net1784));
 sky130_fd_sc_hd__clkbuf_2 wire1785 (.A(net400),
    .X(net1785));
 sky130_fd_sc_hd__buf_6 wire1786 (.A(net1787),
    .X(net1786));
 sky130_fd_sc_hd__buf_6 wire1787 (.A(net1788),
    .X(net1787));
 sky130_fd_sc_hd__buf_4 wire1788 (.A(net1789),
    .X(net1788));
 sky130_fd_sc_hd__clkbuf_2 wire1789 (.A(net399),
    .X(net1789));
 sky130_fd_sc_hd__buf_6 wire1790 (.A(net1791),
    .X(net1790));
 sky130_fd_sc_hd__buf_6 wire1791 (.A(net1792),
    .X(net1791));
 sky130_fd_sc_hd__buf_4 wire1792 (.A(net1793),
    .X(net1792));
 sky130_fd_sc_hd__clkbuf_2 wire1793 (.A(net398),
    .X(net1793));
 sky130_fd_sc_hd__buf_4 wire1794 (.A(net1795),
    .X(net1794));
 sky130_fd_sc_hd__buf_6 wire1795 (.A(net1796),
    .X(net1795));
 sky130_fd_sc_hd__buf_6 wire1796 (.A(net1797),
    .X(net1796));
 sky130_fd_sc_hd__buf_4 wire1797 (.A(net1798),
    .X(net1797));
 sky130_fd_sc_hd__clkbuf_2 wire1798 (.A(net397),
    .X(net1798));
 sky130_fd_sc_hd__buf_6 wire1799 (.A(net1800),
    .X(net1799));
 sky130_fd_sc_hd__buf_4 wire1800 (.A(net1801),
    .X(net1800));
 sky130_fd_sc_hd__clkbuf_2 wire1801 (.A(net396),
    .X(net1801));
 sky130_fd_sc_hd__buf_4 wire1802 (.A(net1803),
    .X(net1802));
 sky130_fd_sc_hd__buf_6 wire1803 (.A(net1804),
    .X(net1803));
 sky130_fd_sc_hd__buf_6 wire1804 (.A(net1805),
    .X(net1804));
 sky130_fd_sc_hd__buf_4 wire1805 (.A(net1806),
    .X(net1805));
 sky130_fd_sc_hd__clkbuf_2 wire1806 (.A(net395),
    .X(net1806));
 sky130_fd_sc_hd__buf_6 wire1807 (.A(net1808),
    .X(net1807));
 sky130_fd_sc_hd__buf_6 wire1808 (.A(net1809),
    .X(net1808));
 sky130_fd_sc_hd__buf_4 wire1809 (.A(net1810),
    .X(net1809));
 sky130_fd_sc_hd__clkbuf_2 wire1810 (.A(net1811),
    .X(net1810));
 sky130_fd_sc_hd__clkbuf_2 wire1811 (.A(net394),
    .X(net1811));
 sky130_fd_sc_hd__buf_2 wire1812 (.A(net1813),
    .X(net1812));
 sky130_fd_sc_hd__clkbuf_2 wire1813 (.A(net1814),
    .X(net1813));
 sky130_fd_sc_hd__clkbuf_2 wire1814 (.A(net393),
    .X(net1814));
 sky130_fd_sc_hd__buf_6 wire1815 (.A(net1816),
    .X(net1815));
 sky130_fd_sc_hd__buf_4 wire1816 (.A(net1817),
    .X(net1816));
 sky130_fd_sc_hd__clkbuf_2 wire1817 (.A(net392),
    .X(net1817));
 sky130_fd_sc_hd__buf_6 wire1818 (.A(net1819),
    .X(net1818));
 sky130_fd_sc_hd__buf_4 wire1819 (.A(net1820),
    .X(net1819));
 sky130_fd_sc_hd__clkbuf_2 wire1820 (.A(net1821),
    .X(net1820));
 sky130_fd_sc_hd__clkbuf_2 wire1821 (.A(net391),
    .X(net1821));
 sky130_fd_sc_hd__clkbuf_2 wire1822 (.A(net1823),
    .X(net1822));
 sky130_fd_sc_hd__clkbuf_2 wire1823 (.A(net390),
    .X(net1823));
 sky130_fd_sc_hd__clkbuf_2 wire1824 (.A(net1825),
    .X(net1824));
 sky130_fd_sc_hd__clkbuf_2 wire1825 (.A(net389),
    .X(net1825));
 sky130_fd_sc_hd__buf_4 wire1826 (.A(net1827),
    .X(net1826));
 sky130_fd_sc_hd__buf_6 wire1827 (.A(net1828),
    .X(net1827));
 sky130_fd_sc_hd__buf_6 wire1828 (.A(net1829),
    .X(net1828));
 sky130_fd_sc_hd__buf_4 wire1829 (.A(net1830),
    .X(net1829));
 sky130_fd_sc_hd__clkbuf_2 wire1830 (.A(net388),
    .X(net1830));
 sky130_fd_sc_hd__clkbuf_2 wire1831 (.A(net1832),
    .X(net1831));
 sky130_fd_sc_hd__clkbuf_2 wire1832 (.A(net386),
    .X(net1832));
 sky130_fd_sc_hd__clkbuf_2 wire1833 (.A(net1834),
    .X(net1833));
 sky130_fd_sc_hd__clkbuf_2 max_length1834 (.A(net385),
    .X(net1834));
 sky130_fd_sc_hd__clkbuf_2 wire1835 (.A(net384),
    .X(net1835));
 sky130_fd_sc_hd__clkbuf_2 wire1836 (.A(net1837),
    .X(net1836));
 sky130_fd_sc_hd__clkbuf_2 wire1837 (.A(net383),
    .X(net1837));
 sky130_fd_sc_hd__clkbuf_2 wire1838 (.A(net382),
    .X(net1838));
 sky130_fd_sc_hd__clkbuf_2 wire1839 (.A(net381),
    .X(net1839));
 sky130_fd_sc_hd__clkbuf_2 wire1840 (.A(net380),
    .X(net1840));
 sky130_fd_sc_hd__clkbuf_2 wire1841 (.A(net1842),
    .X(net1841));
 sky130_fd_sc_hd__buf_2 wire1842 (.A(net374),
    .X(net1842));
 sky130_fd_sc_hd__buf_6 wire1843 (.A(net1844),
    .X(net1843));
 sky130_fd_sc_hd__clkbuf_2 wire1844 (.A(net373),
    .X(net1844));
 sky130_fd_sc_hd__buf_4 wire1845 (.A(net1846),
    .X(net1845));
 sky130_fd_sc_hd__clkbuf_2 wire1846 (.A(net372),
    .X(net1846));
 sky130_fd_sc_hd__buf_4 wire1847 (.A(net1848),
    .X(net1847));
 sky130_fd_sc_hd__clkbuf_2 wire1848 (.A(net371),
    .X(net1848));
 sky130_fd_sc_hd__buf_4 wire1849 (.A(net1850),
    .X(net1849));
 sky130_fd_sc_hd__clkbuf_2 wire1850 (.A(net370),
    .X(net1850));
 sky130_fd_sc_hd__buf_4 wire1851 (.A(net1852),
    .X(net1851));
 sky130_fd_sc_hd__clkbuf_2 wire1852 (.A(net369),
    .X(net1852));
 sky130_fd_sc_hd__buf_4 wire1853 (.A(net1854),
    .X(net1853));
 sky130_fd_sc_hd__clkbuf_2 wire1854 (.A(net368),
    .X(net1854));
 sky130_fd_sc_hd__buf_4 wire1855 (.A(net1856),
    .X(net1855));
 sky130_fd_sc_hd__clkbuf_2 wire1856 (.A(net367),
    .X(net1856));
 sky130_fd_sc_hd__buf_4 wire1857 (.A(net1858),
    .X(net1857));
 sky130_fd_sc_hd__clkbuf_2 wire1858 (.A(net366),
    .X(net1858));
 sky130_fd_sc_hd__clkbuf_2 wire1859 (.A(net1860),
    .X(net1859));
 sky130_fd_sc_hd__buf_2 wire1860 (.A(net364),
    .X(net1860));
 sky130_fd_sc_hd__buf_4 wire1861 (.A(net1862),
    .X(net1861));
 sky130_fd_sc_hd__clkbuf_2 wire1862 (.A(net363),
    .X(net1862));
 sky130_fd_sc_hd__buf_4 wire1863 (.A(net1864),
    .X(net1863));
 sky130_fd_sc_hd__clkbuf_2 wire1864 (.A(net362),
    .X(net1864));
 sky130_fd_sc_hd__buf_4 wire1865 (.A(net1866),
    .X(net1865));
 sky130_fd_sc_hd__clkbuf_2 wire1866 (.A(net361),
    .X(net1866));
 sky130_fd_sc_hd__buf_2 wire1867 (.A(net360),
    .X(net1867));
 sky130_fd_sc_hd__buf_4 wire1868 (.A(net1869),
    .X(net1868));
 sky130_fd_sc_hd__clkbuf_2 wire1869 (.A(net359),
    .X(net1869));
 sky130_fd_sc_hd__buf_2 wire1870 (.A(net358),
    .X(net1870));
 sky130_fd_sc_hd__buf_2 wire1871 (.A(net357),
    .X(net1871));
 sky130_fd_sc_hd__buf_2 wire1872 (.A(net356),
    .X(net1872));
 sky130_fd_sc_hd__clkbuf_2 wire1873 (.A(net355),
    .X(net1873));
 sky130_fd_sc_hd__buf_2 wire1874 (.A(net353),
    .X(net1874));
 sky130_fd_sc_hd__clkbuf_2 wire1875 (.A(net352),
    .X(net1875));
 sky130_fd_sc_hd__buf_2 wire1876 (.A(net351),
    .X(net1876));
 sky130_fd_sc_hd__clkbuf_2 wire1877 (.A(net1878),
    .X(net1877));
 sky130_fd_sc_hd__buf_2 wire1878 (.A(net350),
    .X(net1878));
 sky130_fd_sc_hd__clkbuf_2 wire1879 (.A(net349),
    .X(net1879));
 sky130_fd_sc_hd__clkbuf_2 wire1880 (.A(net1881),
    .X(net1880));
 sky130_fd_sc_hd__clkbuf_2 max_length1881 (.A(net348),
    .X(net1881));
 sky130_fd_sc_hd__clkbuf_2 wire1882 (.A(net347),
    .X(net1882));
 sky130_fd_sc_hd__clkbuf_2 wire1883 (.A(net347),
    .X(net1883));
 sky130_fd_sc_hd__clkbuf_2 wire1884 (.A(net346),
    .X(net1884));
 sky130_fd_sc_hd__clkbuf_2 wire1885 (.A(net345),
    .X(net1885));
 sky130_fd_sc_hd__buf_2 wire1886 (.A(net344),
    .X(net1886));
 sky130_fd_sc_hd__clkbuf_2 wire1887 (.A(net1888),
    .X(net1887));
 sky130_fd_sc_hd__clkbuf_2 wire1888 (.A(net342),
    .X(net1888));
 sky130_fd_sc_hd__clkbuf_2 max_length1889 (.A(net342),
    .X(net1889));
 sky130_fd_sc_hd__clkbuf_2 wire1890 (.A(net341),
    .X(net1890));
 sky130_fd_sc_hd__clkbuf_2 wire1891 (.A(net340),
    .X(net1891));
 sky130_fd_sc_hd__clkbuf_2 wire1892 (.A(net1893),
    .X(net1892));
 sky130_fd_sc_hd__clkbuf_2 max_length1893 (.A(net340),
    .X(net1893));
 sky130_fd_sc_hd__clkbuf_2 wire1894 (.A(net34),
    .X(net1894));
 sky130_fd_sc_hd__clkbuf_2 wire1895 (.A(net338),
    .X(net1895));
 sky130_fd_sc_hd__clkbuf_2 wire1896 (.A(net1898),
    .X(net1896));
 sky130_fd_sc_hd__clkbuf_2 wire1897 (.A(net337),
    .X(net1897));
 sky130_fd_sc_hd__clkbuf_2 max_length1898 (.A(net337),
    .X(net1898));
 sky130_fd_sc_hd__clkbuf_2 wire1899 (.A(net336),
    .X(net1899));
 sky130_fd_sc_hd__clkbuf_2 wire1900 (.A(net335),
    .X(net1900));
 sky130_fd_sc_hd__clkbuf_2 wire1901 (.A(net334),
    .X(net1901));
 sky130_fd_sc_hd__clkbuf_2 max_length1902 (.A(net334),
    .X(net1902));
 sky130_fd_sc_hd__clkbuf_2 wire1903 (.A(net333),
    .X(net1903));
 sky130_fd_sc_hd__buf_2 wire1904 (.A(net1905),
    .X(net1904));
 sky130_fd_sc_hd__clkbuf_2 wire1905 (.A(net1906),
    .X(net1905));
 sky130_fd_sc_hd__clkbuf_2 max_length1906 (.A(net330),
    .X(net1906));
 sky130_fd_sc_hd__clkbuf_2 wire1907 (.A(net33),
    .X(net1907));
 sky130_fd_sc_hd__buf_2 wire1908 (.A(net1909),
    .X(net1908));
 sky130_fd_sc_hd__clkbuf_2 wire1909 (.A(net329),
    .X(net1909));
 sky130_fd_sc_hd__clkbuf_2 max_length1910 (.A(net329),
    .X(net1910));
 sky130_fd_sc_hd__buf_2 wire1911 (.A(net1912),
    .X(net1911));
 sky130_fd_sc_hd__clkbuf_2 wire1912 (.A(net328),
    .X(net1912));
 sky130_fd_sc_hd__clkbuf_2 wire1913 (.A(net325),
    .X(net1913));
 sky130_fd_sc_hd__clkbuf_2 wire1914 (.A(net1915),
    .X(net1914));
 sky130_fd_sc_hd__clkbuf_2 wire1915 (.A(net325),
    .X(net1915));
 sky130_fd_sc_hd__clkbuf_2 wire1916 (.A(net323),
    .X(net1916));
 sky130_fd_sc_hd__clkbuf_2 wire1917 (.A(net322),
    .X(net1917));
 sky130_fd_sc_hd__clkbuf_2 max_length1918 (.A(net322),
    .X(net1918));
 sky130_fd_sc_hd__clkbuf_2 wire1919 (.A(net32),
    .X(net1919));
 sky130_fd_sc_hd__buf_2 wire1920 (.A(net1921),
    .X(net1920));
 sky130_fd_sc_hd__clkbuf_2 wire1921 (.A(net318),
    .X(net1921));
 sky130_fd_sc_hd__clkbuf_2 wire1922 (.A(net316),
    .X(net1922));
 sky130_fd_sc_hd__clkbuf_2 wire1923 (.A(net31),
    .X(net1923));
 sky130_fd_sc_hd__clkbuf_2 wire1924 (.A(net309),
    .X(net1924));
 sky130_fd_sc_hd__clkbuf_2 max_length1925 (.A(net309),
    .X(net1925));
 sky130_fd_sc_hd__buf_2 wire1926 (.A(net307),
    .X(net1926));
 sky130_fd_sc_hd__clkbuf_2 wire1927 (.A(net306),
    .X(net1927));
 sky130_fd_sc_hd__clkbuf_2 max_length1928 (.A(net306),
    .X(net1928));
 sky130_fd_sc_hd__buf_2 wire1929 (.A(net300),
    .X(net1929));
 sky130_fd_sc_hd__buf_6 wire1930 (.A(net1931),
    .X(net1930));
 sky130_fd_sc_hd__buf_6 wire1931 (.A(net1932),
    .X(net1931));
 sky130_fd_sc_hd__buf_4 wire1932 (.A(net1933),
    .X(net1932));
 sky130_fd_sc_hd__buf_6 wire1933 (.A(net1934),
    .X(net1933));
 sky130_fd_sc_hd__buf_6 wire1934 (.A(net1935),
    .X(net1934));
 sky130_fd_sc_hd__buf_4 wire1935 (.A(net1936),
    .X(net1935));
 sky130_fd_sc_hd__clkbuf_2 wire1936 (.A(net3),
    .X(net1936));
 sky130_fd_sc_hd__clkbuf_2 wire1937 (.A(net297),
    .X(net1937));
 sky130_fd_sc_hd__buf_2 wire1938 (.A(net290),
    .X(net1938));
 sky130_fd_sc_hd__clkbuf_4 wire1939 (.A(net289),
    .X(net1939));
 sky130_fd_sc_hd__clkbuf_2 wire1940 (.A(net288),
    .X(net1940));
 sky130_fd_sc_hd__buf_2 wire1941 (.A(net287),
    .X(net1941));
 sky130_fd_sc_hd__clkbuf_2 wire1942 (.A(net286),
    .X(net1942));
 sky130_fd_sc_hd__clkbuf_2 wire1943 (.A(net285),
    .X(net1943));
 sky130_fd_sc_hd__clkbuf_4 wire1944 (.A(net284),
    .X(net1944));
 sky130_fd_sc_hd__clkbuf_2 wire1945 (.A(net1946),
    .X(net1945));
 sky130_fd_sc_hd__clkbuf_2 wire1946 (.A(net283),
    .X(net1946));
 sky130_fd_sc_hd__clkbuf_2 wire1947 (.A(net281),
    .X(net1947));
 sky130_fd_sc_hd__buf_2 wire1948 (.A(net280),
    .X(net1948));
 sky130_fd_sc_hd__clkbuf_2 wire1949 (.A(net28),
    .X(net1949));
 sky130_fd_sc_hd__buf_2 wire1950 (.A(net279),
    .X(net1950));
 sky130_fd_sc_hd__buf_2 wire1951 (.A(net278),
    .X(net1951));
 sky130_fd_sc_hd__buf_2 wire1952 (.A(net277),
    .X(net1952));
 sky130_fd_sc_hd__clkbuf_2 wire1953 (.A(net1954),
    .X(net1953));
 sky130_fd_sc_hd__clkbuf_2 wire1954 (.A(net276),
    .X(net1954));
 sky130_fd_sc_hd__buf_2 wire1955 (.A(net275),
    .X(net1955));
 sky130_fd_sc_hd__buf_2 wire1956 (.A(net274),
    .X(net1956));
 sky130_fd_sc_hd__buf_2 wire1957 (.A(net273),
    .X(net1957));
 sky130_fd_sc_hd__clkbuf_4 wire1958 (.A(net272),
    .X(net1958));
 sky130_fd_sc_hd__clkbuf_2 wire1959 (.A(net270),
    .X(net1959));
 sky130_fd_sc_hd__clkbuf_2 wire1960 (.A(net27),
    .X(net1960));
 sky130_fd_sc_hd__buf_2 wire1961 (.A(net269),
    .X(net1961));
 sky130_fd_sc_hd__clkbuf_2 wire1962 (.A(net268),
    .X(net1962));
 sky130_fd_sc_hd__clkbuf_2 wire1963 (.A(net1964),
    .X(net1963));
 sky130_fd_sc_hd__clkbuf_2 max_length1964 (.A(net267),
    .X(net1964));
 sky130_fd_sc_hd__clkbuf_2 wire1965 (.A(net1966),
    .X(net1965));
 sky130_fd_sc_hd__clkbuf_2 max_length1966 (.A(net266),
    .X(net1966));
 sky130_fd_sc_hd__clkbuf_2 wire1967 (.A(net265),
    .X(net1967));
 sky130_fd_sc_hd__clkbuf_2 wire1968 (.A(net264),
    .X(net1968));
 sky130_fd_sc_hd__clkbuf_2 wire1969 (.A(net1970),
    .X(net1969));
 sky130_fd_sc_hd__clkbuf_2 wire1970 (.A(net263),
    .X(net1970));
 sky130_fd_sc_hd__clkbuf_2 wire1971 (.A(net262),
    .X(net1971));
 sky130_fd_sc_hd__clkbuf_2 wire1972 (.A(net1973),
    .X(net1972));
 sky130_fd_sc_hd__clkbuf_2 wire1973 (.A(net261),
    .X(net1973));
 sky130_fd_sc_hd__clkbuf_2 wire1974 (.A(net259),
    .X(net1974));
 sky130_fd_sc_hd__buf_2 wire1975 (.A(net1976),
    .X(net1975));
 sky130_fd_sc_hd__clkbuf_2 wire1976 (.A(net245),
    .X(net1976));
 sky130_fd_sc_hd__clkbuf_4 wire1977 (.A(net1978),
    .X(net1977));
 sky130_fd_sc_hd__clkbuf_2 wire1978 (.A(net238),
    .X(net1978));
 sky130_fd_sc_hd__clkbuf_2 wire1979 (.A(net234),
    .X(net1979));
 sky130_fd_sc_hd__clkbuf_2 wire1980 (.A(net233),
    .X(net1980));
 sky130_fd_sc_hd__buf_2 wire1981 (.A(net1982),
    .X(net1981));
 sky130_fd_sc_hd__clkbuf_2 wire1982 (.A(net232),
    .X(net1982));
 sky130_fd_sc_hd__clkbuf_2 wire1983 (.A(net1984),
    .X(net1983));
 sky130_fd_sc_hd__clkbuf_2 wire1984 (.A(net231),
    .X(net1984));
 sky130_fd_sc_hd__clkbuf_2 wire1985 (.A(net1986),
    .X(net1985));
 sky130_fd_sc_hd__clkbuf_2 wire1986 (.A(net230),
    .X(net1986));
 sky130_fd_sc_hd__clkbuf_2 wire1987 (.A(net229),
    .X(net1987));
 sky130_fd_sc_hd__clkbuf_2 wire1988 (.A(net228),
    .X(net1988));
 sky130_fd_sc_hd__clkbuf_2 wire1989 (.A(net227),
    .X(net1989));
 sky130_fd_sc_hd__clkbuf_2 wire1990 (.A(net225),
    .X(net1990));
 sky130_fd_sc_hd__clkbuf_2 wire1991 (.A(net217),
    .X(net1991));
 sky130_fd_sc_hd__clkbuf_2 wire1992 (.A(net216),
    .X(net1992));
 sky130_fd_sc_hd__clkbuf_2 wire1993 (.A(net212),
    .X(net1993));
 sky130_fd_sc_hd__clkbuf_2 wire1994 (.A(net209),
    .X(net1994));
 sky130_fd_sc_hd__clkbuf_2 wire1995 (.A(net208),
    .X(net1995));
 sky130_fd_sc_hd__clkbuf_2 wire1996 (.A(net206),
    .X(net1996));
 sky130_fd_sc_hd__clkbuf_2 wire1997 (.A(net205),
    .X(net1997));
 sky130_fd_sc_hd__clkbuf_2 wire1998 (.A(net202),
    .X(net1998));
 sky130_fd_sc_hd__clkbuf_2 wire1999 (.A(net201),
    .X(net1999));
 sky130_fd_sc_hd__clkbuf_2 wire2000 (.A(net199),
    .X(net2000));
 sky130_fd_sc_hd__clkbuf_2 wire2001 (.A(net197),
    .X(net2001));
 sky130_fd_sc_hd__clkbuf_2 wire2002 (.A(net195),
    .X(net2002));
 sky130_fd_sc_hd__clkbuf_2 wire2003 (.A(net191),
    .X(net2003));
 sky130_fd_sc_hd__clkbuf_2 wire2004 (.A(net188),
    .X(net2004));
 sky130_fd_sc_hd__clkbuf_2 wire2005 (.A(net180),
    .X(net2005));
 sky130_fd_sc_hd__clkbuf_2 wire2006 (.A(net175),
    .X(net2006));
 sky130_fd_sc_hd__clkbuf_2 wire2007 (.A(net17),
    .X(net2007));
 sky130_fd_sc_hd__clkbuf_2 wire2008 (.A(net161),
    .X(net2008));
 sky130_fd_sc_hd__clkbuf_2 wire2009 (.A(net159),
    .X(net2009));
 sky130_fd_sc_hd__clkbuf_2 wire2010 (.A(net158),
    .X(net2010));
 sky130_fd_sc_hd__clkbuf_2 wire2011 (.A(net157),
    .X(net2011));
 sky130_fd_sc_hd__clkbuf_2 wire2012 (.A(net156),
    .X(net2012));
 sky130_fd_sc_hd__clkbuf_2 wire2013 (.A(net2014),
    .X(net2013));
 sky130_fd_sc_hd__clkbuf_2 wire2014 (.A(net155),
    .X(net2014));
 sky130_fd_sc_hd__clkbuf_2 wire2015 (.A(net152),
    .X(net2015));
 sky130_fd_sc_hd__clkbuf_2 wire2016 (.A(net151),
    .X(net2016));
 sky130_fd_sc_hd__buf_2 wire2017 (.A(net2018),
    .X(net2017));
 sky130_fd_sc_hd__clkbuf_2 wire2018 (.A(net149),
    .X(net2018));
 sky130_fd_sc_hd__clkbuf_2 wire2019 (.A(net147),
    .X(net2019));
 sky130_fd_sc_hd__clkbuf_2 wire2020 (.A(net2021),
    .X(net2020));
 sky130_fd_sc_hd__clkbuf_2 wire2021 (.A(net146),
    .X(net2021));
 sky130_fd_sc_hd__clkbuf_2 wire2022 (.A(net145),
    .X(net2022));
 sky130_fd_sc_hd__clkbuf_2 wire2023 (.A(net144),
    .X(net2023));
 sky130_fd_sc_hd__clkbuf_2 wire2024 (.A(net143),
    .X(net2024));
 sky130_fd_sc_hd__clkbuf_2 wire2025 (.A(net142),
    .X(net2025));
 sky130_fd_sc_hd__clkbuf_2 wire2026 (.A(net141),
    .X(net2026));
 sky130_fd_sc_hd__clkbuf_2 wire2027 (.A(net2028),
    .X(net2027));
 sky130_fd_sc_hd__clkbuf_2 wire2028 (.A(net140),
    .X(net2028));
 sky130_fd_sc_hd__clkbuf_2 wire2029 (.A(net118),
    .X(net2029));
 sky130_fd_sc_hd__buf_6 wire2030 (.A(net2031),
    .X(net2030));
 sky130_fd_sc_hd__buf_4 wire2031 (.A(net2032),
    .X(net2031));
 sky130_fd_sc_hd__clkbuf_2 wire2032 (.A(net117),
    .X(net2032));
 sky130_fd_sc_hd__buf_2 wire2033 (.A(net2034),
    .X(net2033));
 sky130_fd_sc_hd__clkbuf_2 wire2034 (.A(net2035),
    .X(net2034));
 sky130_fd_sc_hd__clkbuf_2 wire2035 (.A(net116),
    .X(net2035));
 sky130_fd_sc_hd__buf_2 wire2036 (.A(net2037),
    .X(net2036));
 sky130_fd_sc_hd__clkbuf_2 wire2037 (.A(net115),
    .X(net2037));
 sky130_fd_sc_hd__buf_2 wire2038 (.A(net2039),
    .X(net2038));
 sky130_fd_sc_hd__clkbuf_2 wire2039 (.A(net114),
    .X(net2039));
 sky130_fd_sc_hd__buf_2 wire2040 (.A(net2041),
    .X(net2040));
 sky130_fd_sc_hd__clkbuf_2 wire2041 (.A(net2042),
    .X(net2041));
 sky130_fd_sc_hd__clkbuf_2 wire2042 (.A(net113),
    .X(net2042));
 sky130_fd_sc_hd__buf_2 wire2043 (.A(net2044),
    .X(net2043));
 sky130_fd_sc_hd__clkbuf_2 wire2044 (.A(net2045),
    .X(net2044));
 sky130_fd_sc_hd__clkbuf_2 wire2045 (.A(net112),
    .X(net2045));
 sky130_fd_sc_hd__buf_2 wire2046 (.A(net2047),
    .X(net2046));
 sky130_fd_sc_hd__clkbuf_2 wire2047 (.A(net111),
    .X(net2047));
 sky130_fd_sc_hd__buf_2 wire2048 (.A(net2049),
    .X(net2048));
 sky130_fd_sc_hd__clkbuf_2 wire2049 (.A(net2050),
    .X(net2049));
 sky130_fd_sc_hd__clkbuf_2 wire2050 (.A(net110),
    .X(net2050));
 sky130_fd_sc_hd__clkbuf_2 wire2051 (.A(net108),
    .X(net2051));
 sky130_fd_sc_hd__buf_2 wire2052 (.A(net2053),
    .X(net2052));
 sky130_fd_sc_hd__clkbuf_2 wire2053 (.A(net107),
    .X(net2053));
 sky130_fd_sc_hd__buf_2 wire2054 (.A(net2055),
    .X(net2054));
 sky130_fd_sc_hd__clkbuf_2 wire2055 (.A(net2056),
    .X(net2055));
 sky130_fd_sc_hd__clkbuf_2 wire2056 (.A(net106),
    .X(net2056));
 sky130_fd_sc_hd__buf_2 wire2057 (.A(net2058),
    .X(net2057));
 sky130_fd_sc_hd__clkbuf_2 wire2058 (.A(net105),
    .X(net2058));
 sky130_fd_sc_hd__clkbuf_2 wire2059 (.A(net104),
    .X(net2059));
 sky130_fd_sc_hd__buf_2 wire2060 (.A(net2061),
    .X(net2060));
 sky130_fd_sc_hd__clkbuf_2 wire2061 (.A(net103),
    .X(net2061));
 sky130_fd_sc_hd__clkbuf_2 wire2062 (.A(net102),
    .X(net2062));
 sky130_fd_sc_hd__clkbuf_2 wire2063 (.A(net101),
    .X(net2063));
 sky130_fd_sc_hd__clkbuf_2 wire2064 (.A(net2065),
    .X(net2064));
 sky130_fd_sc_hd__clkbuf_2 wire2065 (.A(net100),
    .X(net2065));
 sky130_fd_sc_hd__buf_6 wire2066 (.A(net2067),
    .X(net2066));
 sky130_fd_sc_hd__buf_4 wire2067 (.A(net2068),
    .X(net2067));
 sky130_fd_sc_hd__clkbuf_2 wire2068 (.A(net2069),
    .X(net2068));
 sky130_fd_sc_hd__clkbuf_2 wire2069 (.A(net1),
    .X(net2069));
 sky130_fd_sc_hd__buf_4 wire2070 (.A(net2071),
    .X(net2070));
 sky130_fd_sc_hd__clkbuf_2 wire2071 (.A(net952),
    .X(net2071));
 sky130_fd_sc_hd__buf_6 wire2072 (.A(net2073),
    .X(net2072));
 sky130_fd_sc_hd__clkbuf_2 wire2073 (.A(net2074),
    .X(net2073));
 sky130_fd_sc_hd__clkbuf_2 wire2074 (.A(net954),
    .X(net2074));
 sky130_fd_sc_hd__buf_2 wire2075 (.A(net2076),
    .X(net2075));
 sky130_fd_sc_hd__clkbuf_2 wire2076 (.A(net2077),
    .X(net2076));
 sky130_fd_sc_hd__clkbuf_2 wire2077 (.A(\mprj_logic1[9] ),
    .X(net2077));
 sky130_fd_sc_hd__buf_6 wire2078 (.A(net2079),
    .X(net2078));
 sky130_fd_sc_hd__buf_4 wire2079 (.A(net2080),
    .X(net2079));
 sky130_fd_sc_hd__clkbuf_2 wire2080 (.A(\mprj_logic1[99] ),
    .X(net2080));
 sky130_fd_sc_hd__buf_2 wire2081 (.A(net2082),
    .X(net2081));
 sky130_fd_sc_hd__clkbuf_2 wire2082 (.A(net2083),
    .X(net2082));
 sky130_fd_sc_hd__clkbuf_2 wire2083 (.A(\mprj_logic1[98] ),
    .X(net2083));
 sky130_fd_sc_hd__buf_2 wire2084 (.A(net2085),
    .X(net2084));
 sky130_fd_sc_hd__clkbuf_2 wire2085 (.A(\mprj_logic1[97] ),
    .X(net2085));
 sky130_fd_sc_hd__buf_4 wire2086 (.A(net2087),
    .X(net2086));
 sky130_fd_sc_hd__buf_4 wire2087 (.A(net2088),
    .X(net2087));
 sky130_fd_sc_hd__clkbuf_2 wire2088 (.A(\mprj_logic1[96] ),
    .X(net2088));
 sky130_fd_sc_hd__buf_6 wire2089 (.A(net2090),
    .X(net2089));
 sky130_fd_sc_hd__buf_4 wire2090 (.A(net2091),
    .X(net2090));
 sky130_fd_sc_hd__clkbuf_2 wire2091 (.A(\mprj_logic1[95] ),
    .X(net2091));
 sky130_fd_sc_hd__buf_6 wire2092 (.A(net2093),
    .X(net2092));
 sky130_fd_sc_hd__buf_4 wire2093 (.A(net2094),
    .X(net2093));
 sky130_fd_sc_hd__clkbuf_2 wire2094 (.A(net2095),
    .X(net2094));
 sky130_fd_sc_hd__clkbuf_2 wire2095 (.A(\mprj_logic1[94] ),
    .X(net2095));
 sky130_fd_sc_hd__buf_6 wire2096 (.A(net2097),
    .X(net2096));
 sky130_fd_sc_hd__buf_4 wire2097 (.A(net2098),
    .X(net2097));
 sky130_fd_sc_hd__clkbuf_2 wire2098 (.A(\mprj_logic1[93] ),
    .X(net2098));
 sky130_fd_sc_hd__buf_6 wire2099 (.A(net2100),
    .X(net2099));
 sky130_fd_sc_hd__buf_4 wire2100 (.A(net2101),
    .X(net2100));
 sky130_fd_sc_hd__clkbuf_2 wire2101 (.A(net2102),
    .X(net2101));
 sky130_fd_sc_hd__clkbuf_2 wire2102 (.A(\mprj_logic1[92] ),
    .X(net2102));
 sky130_fd_sc_hd__buf_2 wire2103 (.A(net2104),
    .X(net2103));
 sky130_fd_sc_hd__clkbuf_2 wire2104 (.A(net2105),
    .X(net2104));
 sky130_fd_sc_hd__clkbuf_2 wire2105 (.A(\mprj_logic1[91] ),
    .X(net2105));
 sky130_fd_sc_hd__buf_2 wire2106 (.A(net2107),
    .X(net2106));
 sky130_fd_sc_hd__clkbuf_2 wire2107 (.A(net2108),
    .X(net2107));
 sky130_fd_sc_hd__clkbuf_2 wire2108 (.A(\mprj_logic1[90] ),
    .X(net2108));
 sky130_fd_sc_hd__buf_2 wire2109 (.A(net2110),
    .X(net2109));
 sky130_fd_sc_hd__clkbuf_2 wire2110 (.A(\mprj_logic1[8] ),
    .X(net2110));
 sky130_fd_sc_hd__buf_6 wire2111 (.A(net2112),
    .X(net2111));
 sky130_fd_sc_hd__buf_4 wire2112 (.A(net2113),
    .X(net2112));
 sky130_fd_sc_hd__clkbuf_2 wire2113 (.A(net2114),
    .X(net2113));
 sky130_fd_sc_hd__clkbuf_2 wire2114 (.A(\mprj_logic1[89] ),
    .X(net2114));
 sky130_fd_sc_hd__buf_6 wire2115 (.A(net2116),
    .X(net2115));
 sky130_fd_sc_hd__buf_4 wire2116 (.A(net2117),
    .X(net2116));
 sky130_fd_sc_hd__clkbuf_2 wire2117 (.A(net2118),
    .X(net2117));
 sky130_fd_sc_hd__clkbuf_2 wire2118 (.A(\mprj_logic1[88] ),
    .X(net2118));
 sky130_fd_sc_hd__buf_6 wire2119 (.A(net2120),
    .X(net2119));
 sky130_fd_sc_hd__buf_4 wire2120 (.A(net2121),
    .X(net2120));
 sky130_fd_sc_hd__clkbuf_2 wire2121 (.A(\mprj_logic1[87] ),
    .X(net2121));
 sky130_fd_sc_hd__buf_2 wire2122 (.A(net2123),
    .X(net2122));
 sky130_fd_sc_hd__clkbuf_2 wire2123 (.A(net2124),
    .X(net2123));
 sky130_fd_sc_hd__clkbuf_2 wire2124 (.A(\mprj_logic1[86] ),
    .X(net2124));
 sky130_fd_sc_hd__buf_6 wire2125 (.A(net2126),
    .X(net2125));
 sky130_fd_sc_hd__buf_4 wire2126 (.A(net2127),
    .X(net2126));
 sky130_fd_sc_hd__clkbuf_2 wire2127 (.A(net2128),
    .X(net2127));
 sky130_fd_sc_hd__clkbuf_2 wire2128 (.A(\mprj_logic1[85] ),
    .X(net2128));
 sky130_fd_sc_hd__buf_6 wire2129 (.A(net2130),
    .X(net2129));
 sky130_fd_sc_hd__buf_4 wire2130 (.A(net2131),
    .X(net2130));
 sky130_fd_sc_hd__clkbuf_2 wire2131 (.A(net2132),
    .X(net2131));
 sky130_fd_sc_hd__clkbuf_2 wire2132 (.A(\mprj_logic1[84] ),
    .X(net2132));
 sky130_fd_sc_hd__buf_6 wire2133 (.A(net2134),
    .X(net2133));
 sky130_fd_sc_hd__buf_4 wire2134 (.A(net2135),
    .X(net2134));
 sky130_fd_sc_hd__clkbuf_2 wire2135 (.A(net2136),
    .X(net2135));
 sky130_fd_sc_hd__clkbuf_2 wire2136 (.A(\mprj_logic1[83] ),
    .X(net2136));
 sky130_fd_sc_hd__buf_6 wire2137 (.A(net2138),
    .X(net2137));
 sky130_fd_sc_hd__buf_4 wire2138 (.A(net2139),
    .X(net2138));
 sky130_fd_sc_hd__clkbuf_2 wire2139 (.A(\mprj_logic1[82] ),
    .X(net2139));
 sky130_fd_sc_hd__buf_6 wire2140 (.A(net2141),
    .X(net2140));
 sky130_fd_sc_hd__buf_6 wire2141 (.A(net2142),
    .X(net2141));
 sky130_fd_sc_hd__buf_4 wire2142 (.A(net2143),
    .X(net2142));
 sky130_fd_sc_hd__clkbuf_2 wire2143 (.A(\mprj_logic1[81] ),
    .X(net2143));
 sky130_fd_sc_hd__buf_6 wire2144 (.A(net2145),
    .X(net2144));
 sky130_fd_sc_hd__buf_4 wire2145 (.A(net2146),
    .X(net2145));
 sky130_fd_sc_hd__clkbuf_2 wire2146 (.A(net2147),
    .X(net2146));
 sky130_fd_sc_hd__clkbuf_2 wire2147 (.A(\mprj_logic1[80] ),
    .X(net2147));
 sky130_fd_sc_hd__buf_2 wire2148 (.A(net2149),
    .X(net2148));
 sky130_fd_sc_hd__clkbuf_2 wire2149 (.A(\mprj_logic1[7] ),
    .X(net2149));
 sky130_fd_sc_hd__buf_6 wire2150 (.A(net2151),
    .X(net2150));
 sky130_fd_sc_hd__buf_4 wire2151 (.A(net2152),
    .X(net2151));
 sky130_fd_sc_hd__clkbuf_2 wire2152 (.A(\mprj_logic1[79] ),
    .X(net2152));
 sky130_fd_sc_hd__buf_6 wire2153 (.A(net2154),
    .X(net2153));
 sky130_fd_sc_hd__buf_4 wire2154 (.A(net2155),
    .X(net2154));
 sky130_fd_sc_hd__clkbuf_2 wire2155 (.A(\mprj_logic1[78] ),
    .X(net2155));
 sky130_fd_sc_hd__buf_6 wire2156 (.A(net2157),
    .X(net2156));
 sky130_fd_sc_hd__buf_4 wire2157 (.A(net2158),
    .X(net2157));
 sky130_fd_sc_hd__clkbuf_2 wire2158 (.A(\mprj_logic1[77] ),
    .X(net2158));
 sky130_fd_sc_hd__buf_4 wire2159 (.A(net2160),
    .X(net2159));
 sky130_fd_sc_hd__clkbuf_2 wire2160 (.A(net2161),
    .X(net2160));
 sky130_fd_sc_hd__clkbuf_2 wire2161 (.A(\mprj_logic1[76] ),
    .X(net2161));
 sky130_fd_sc_hd__buf_6 wire2162 (.A(net2163),
    .X(net2162));
 sky130_fd_sc_hd__buf_4 wire2163 (.A(net2164),
    .X(net2163));
 sky130_fd_sc_hd__clkbuf_2 wire2164 (.A(\mprj_logic1[75] ),
    .X(net2164));
 sky130_fd_sc_hd__buf_6 wire2165 (.A(net2166),
    .X(net2165));
 sky130_fd_sc_hd__buf_4 wire2166 (.A(net2167),
    .X(net2166));
 sky130_fd_sc_hd__clkbuf_2 wire2167 (.A(\mprj_logic1[74] ),
    .X(net2167));
 sky130_fd_sc_hd__clkbuf_2 wire2168 (.A(\mprj_logic1[73] ),
    .X(net2168));
 sky130_fd_sc_hd__clkbuf_2 wire2169 (.A(\mprj_logic1[72] ),
    .X(net2169));
 sky130_fd_sc_hd__clkbuf_2 wire2170 (.A(net2171),
    .X(net2170));
 sky130_fd_sc_hd__clkbuf_2 wire2171 (.A(\mprj_logic1[71] ),
    .X(net2171));
 sky130_fd_sc_hd__buf_2 wire2172 (.A(net2173),
    .X(net2172));
 sky130_fd_sc_hd__clkbuf_2 wire2173 (.A(\mprj_logic1[70] ),
    .X(net2173));
 sky130_fd_sc_hd__buf_2 wire2174 (.A(net2175),
    .X(net2174));
 sky130_fd_sc_hd__clkbuf_2 wire2175 (.A(\mprj_logic1[6] ),
    .X(net2175));
 sky130_fd_sc_hd__buf_6 wire2176 (.A(net2177),
    .X(net2176));
 sky130_fd_sc_hd__buf_4 wire2177 (.A(net2178),
    .X(net2177));
 sky130_fd_sc_hd__clkbuf_2 wire2178 (.A(net2179),
    .X(net2178));
 sky130_fd_sc_hd__clkbuf_2 wire2179 (.A(\mprj_logic1[69] ),
    .X(net2179));
 sky130_fd_sc_hd__buf_2 wire2180 (.A(net2181),
    .X(net2180));
 sky130_fd_sc_hd__clkbuf_2 wire2181 (.A(\mprj_logic1[68] ),
    .X(net2181));
 sky130_fd_sc_hd__buf_2 wire2182 (.A(net2183),
    .X(net2182));
 sky130_fd_sc_hd__clkbuf_2 wire2183 (.A(net2184),
    .X(net2183));
 sky130_fd_sc_hd__clkbuf_2 wire2184 (.A(\mprj_logic1[67] ),
    .X(net2184));
 sky130_fd_sc_hd__buf_2 wire2185 (.A(net2186),
    .X(net2185));
 sky130_fd_sc_hd__clkbuf_2 wire2186 (.A(net2187),
    .X(net2186));
 sky130_fd_sc_hd__clkbuf_2 wire2187 (.A(\mprj_logic1[66] ),
    .X(net2187));
 sky130_fd_sc_hd__clkbuf_2 wire2188 (.A(\mprj_logic1[65] ),
    .X(net2188));
 sky130_fd_sc_hd__clkbuf_2 wire2189 (.A(\mprj_logic1[64] ),
    .X(net2189));
 sky130_fd_sc_hd__clkbuf_2 wire2190 (.A(\mprj_logic1[63] ),
    .X(net2190));
 sky130_fd_sc_hd__clkbuf_2 wire2191 (.A(net2192),
    .X(net2191));
 sky130_fd_sc_hd__clkbuf_2 wire2192 (.A(\mprj_logic1[62] ),
    .X(net2192));
 sky130_fd_sc_hd__clkbuf_2 wire2193 (.A(\mprj_logic1[61] ),
    .X(net2193));
 sky130_fd_sc_hd__clkbuf_2 wire2194 (.A(\mprj_logic1[60] ),
    .X(net2194));
 sky130_fd_sc_hd__clkbuf_2 wire2195 (.A(\mprj_logic1[5] ),
    .X(net2195));
 sky130_fd_sc_hd__clkbuf_2 wire2196 (.A(net2197),
    .X(net2196));
 sky130_fd_sc_hd__clkbuf_2 wire2197 (.A(\mprj_logic1[59] ),
    .X(net2197));
 sky130_fd_sc_hd__clkbuf_2 wire2198 (.A(\mprj_logic1[58] ),
    .X(net2198));
 sky130_fd_sc_hd__clkbuf_2 wire2199 (.A(\mprj_logic1[56] ),
    .X(net2199));
 sky130_fd_sc_hd__buf_2 wire2200 (.A(net2201),
    .X(net2200));
 sky130_fd_sc_hd__clkbuf_2 wire2201 (.A(\mprj_logic1[55] ),
    .X(net2201));
 sky130_fd_sc_hd__clkbuf_2 wire2202 (.A(net2203),
    .X(net2202));
 sky130_fd_sc_hd__clkbuf_2 wire2203 (.A(\mprj_logic1[54] ),
    .X(net2203));
 sky130_fd_sc_hd__clkbuf_2 wire2204 (.A(net2205),
    .X(net2204));
 sky130_fd_sc_hd__clkbuf_2 wire2205 (.A(\mprj_logic1[53] ),
    .X(net2205));
 sky130_fd_sc_hd__clkbuf_2 wire2206 (.A(\mprj_logic1[52] ),
    .X(net2206));
 sky130_fd_sc_hd__clkbuf_2 wire2207 (.A(\mprj_logic1[51] ),
    .X(net2207));
 sky130_fd_sc_hd__clkbuf_2 wire2208 (.A(\mprj_logic1[4] ),
    .X(net2208));
 sky130_fd_sc_hd__clkbuf_2 wire2209 (.A(\mprj_logic1[49] ),
    .X(net2209));
 sky130_fd_sc_hd__buf_6 wire2210 (.A(net2211),
    .X(net2210));
 sky130_fd_sc_hd__buf_4 wire2211 (.A(net2212),
    .X(net2211));
 sky130_fd_sc_hd__clkbuf_2 wire2212 (.A(net2213),
    .X(net2212));
 sky130_fd_sc_hd__clkbuf_2 wire2213 (.A(\mprj_logic1[462] ),
    .X(net2213));
 sky130_fd_sc_hd__buf_6 wire2214 (.A(net2215),
    .X(net2214));
 sky130_fd_sc_hd__buf_6 wire2215 (.A(net2216),
    .X(net2215));
 sky130_fd_sc_hd__buf_4 wire2216 (.A(net2217),
    .X(net2216));
 sky130_fd_sc_hd__clkbuf_2 wire2217 (.A(net951),
    .X(net2217));
 sky130_fd_sc_hd__buf_6 wire2218 (.A(net2219),
    .X(net2218));
 sky130_fd_sc_hd__buf_4 wire2219 (.A(net2220),
    .X(net2219));
 sky130_fd_sc_hd__clkbuf_2 wire2220 (.A(\mprj_logic1[460] ),
    .X(net2220));
 sky130_fd_sc_hd__buf_6 wire2221 (.A(net2222),
    .X(net2221));
 sky130_fd_sc_hd__buf_4 wire2222 (.A(net2223),
    .X(net2222));
 sky130_fd_sc_hd__clkbuf_2 wire2223 (.A(net2224),
    .X(net2223));
 sky130_fd_sc_hd__clkbuf_2 wire2224 (.A(\mprj_logic1[459] ),
    .X(net2224));
 sky130_fd_sc_hd__buf_6 wire2225 (.A(net2226),
    .X(net2225));
 sky130_fd_sc_hd__buf_4 wire2226 (.A(net2227),
    .X(net2226));
 sky130_fd_sc_hd__clkbuf_2 wire2227 (.A(net2228),
    .X(net2227));
 sky130_fd_sc_hd__clkbuf_2 wire2228 (.A(\mprj_logic1[458] ),
    .X(net2228));
 sky130_fd_sc_hd__buf_2 wire2229 (.A(net2230),
    .X(net2229));
 sky130_fd_sc_hd__clkbuf_2 wire2230 (.A(\mprj_logic1[457] ),
    .X(net2230));
 sky130_fd_sc_hd__buf_6 wire2231 (.A(net2232),
    .X(net2231));
 sky130_fd_sc_hd__buf_4 wire2232 (.A(net2233),
    .X(net2232));
 sky130_fd_sc_hd__clkbuf_2 wire2233 (.A(\mprj_logic1[456] ),
    .X(net2233));
 sky130_fd_sc_hd__buf_4 wire2234 (.A(net2235),
    .X(net2234));
 sky130_fd_sc_hd__clkbuf_2 wire2235 (.A(net2236),
    .X(net2235));
 sky130_fd_sc_hd__clkbuf_2 wire2236 (.A(\mprj_logic1[455] ),
    .X(net2236));
 sky130_fd_sc_hd__buf_6 wire2237 (.A(net2238),
    .X(net2237));
 sky130_fd_sc_hd__buf_4 wire2238 (.A(net2239),
    .X(net2238));
 sky130_fd_sc_hd__clkbuf_2 wire2239 (.A(\mprj_logic1[454] ),
    .X(net2239));
 sky130_fd_sc_hd__buf_6 wire2240 (.A(net2241),
    .X(net2240));
 sky130_fd_sc_hd__buf_4 wire2241 (.A(net2242),
    .X(net2241));
 sky130_fd_sc_hd__clkbuf_2 wire2242 (.A(\mprj_logic1[453] ),
    .X(net2242));
 sky130_fd_sc_hd__buf_6 wire2243 (.A(net2244),
    .X(net2243));
 sky130_fd_sc_hd__buf_4 wire2244 (.A(net2245),
    .X(net2244));
 sky130_fd_sc_hd__clkbuf_2 wire2245 (.A(\mprj_logic1[452] ),
    .X(net2245));
 sky130_fd_sc_hd__buf_6 wire2246 (.A(net2247),
    .X(net2246));
 sky130_fd_sc_hd__buf_4 wire2247 (.A(net2248),
    .X(net2247));
 sky130_fd_sc_hd__clkbuf_2 wire2248 (.A(\mprj_logic1[451] ),
    .X(net2248));
 sky130_fd_sc_hd__buf_6 wire2249 (.A(net2250),
    .X(net2249));
 sky130_fd_sc_hd__buf_6 wire2250 (.A(net2251),
    .X(net2250));
 sky130_fd_sc_hd__buf_4 wire2251 (.A(net2252),
    .X(net2251));
 sky130_fd_sc_hd__clkbuf_2 wire2252 (.A(\mprj_logic1[450] ),
    .X(net2252));
 sky130_fd_sc_hd__clkbuf_2 wire2253 (.A(\mprj_logic1[44] ),
    .X(net2253));
 sky130_fd_sc_hd__buf_2 wire2254 (.A(net2255),
    .X(net2254));
 sky130_fd_sc_hd__clkbuf_2 wire2255 (.A(\mprj_logic1[449] ),
    .X(net2255));
 sky130_fd_sc_hd__buf_6 wire2256 (.A(net2257),
    .X(net2256));
 sky130_fd_sc_hd__buf_4 wire2257 (.A(net2258),
    .X(net2257));
 sky130_fd_sc_hd__clkbuf_2 wire2258 (.A(\mprj_logic1[448] ),
    .X(net2258));
 sky130_fd_sc_hd__buf_2 wire2259 (.A(net2260),
    .X(net2259));
 sky130_fd_sc_hd__clkbuf_2 wire2260 (.A(net2261),
    .X(net2260));
 sky130_fd_sc_hd__clkbuf_2 wire2261 (.A(\mprj_logic1[447] ),
    .X(net2261));
 sky130_fd_sc_hd__buf_2 wire2262 (.A(net2263),
    .X(net2262));
 sky130_fd_sc_hd__clkbuf_2 wire2263 (.A(\mprj_logic1[446] ),
    .X(net2263));
 sky130_fd_sc_hd__buf_6 wire2264 (.A(net2265),
    .X(net2264));
 sky130_fd_sc_hd__buf_6 wire2265 (.A(net2266),
    .X(net2265));
 sky130_fd_sc_hd__buf_4 wire2266 (.A(net2267),
    .X(net2266));
 sky130_fd_sc_hd__clkbuf_2 wire2267 (.A(\mprj_logic1[445] ),
    .X(net2267));
 sky130_fd_sc_hd__buf_2 wire2268 (.A(net2269),
    .X(net2268));
 sky130_fd_sc_hd__clkbuf_2 wire2269 (.A(\mprj_logic1[444] ),
    .X(net2269));
 sky130_fd_sc_hd__buf_6 wire2270 (.A(net2271),
    .X(net2270));
 sky130_fd_sc_hd__buf_4 wire2271 (.A(net2272),
    .X(net2271));
 sky130_fd_sc_hd__clkbuf_2 wire2272 (.A(\mprj_logic1[443] ),
    .X(net2272));
 sky130_fd_sc_hd__buf_6 wire2273 (.A(net2274),
    .X(net2273));
 sky130_fd_sc_hd__buf_4 wire2274 (.A(net2275),
    .X(net2274));
 sky130_fd_sc_hd__clkbuf_2 wire2275 (.A(\mprj_logic1[442] ),
    .X(net2275));
 sky130_fd_sc_hd__buf_6 wire2276 (.A(net2277),
    .X(net2276));
 sky130_fd_sc_hd__buf_4 wire2277 (.A(net2278),
    .X(net2277));
 sky130_fd_sc_hd__clkbuf_2 wire2278 (.A(\mprj_logic1[441] ),
    .X(net2278));
 sky130_fd_sc_hd__buf_2 wire2279 (.A(net2280),
    .X(net2279));
 sky130_fd_sc_hd__clkbuf_2 wire2280 (.A(\mprj_logic1[440] ),
    .X(net2280));
 sky130_fd_sc_hd__buf_6 wire2281 (.A(net2282),
    .X(net2281));
 sky130_fd_sc_hd__buf_4 wire2282 (.A(net2283),
    .X(net2282));
 sky130_fd_sc_hd__clkbuf_2 wire2283 (.A(\mprj_logic1[439] ),
    .X(net2283));
 sky130_fd_sc_hd__buf_2 wire2284 (.A(net2285),
    .X(net2284));
 sky130_fd_sc_hd__clkbuf_2 wire2285 (.A(net2286),
    .X(net2285));
 sky130_fd_sc_hd__clkbuf_2 wire2286 (.A(\mprj_logic1[438] ),
    .X(net2286));
 sky130_fd_sc_hd__buf_6 wire2287 (.A(net2288),
    .X(net2287));
 sky130_fd_sc_hd__buf_4 wire2288 (.A(net2289),
    .X(net2288));
 sky130_fd_sc_hd__clkbuf_2 wire2289 (.A(\mprj_logic1[437] ),
    .X(net2289));
 sky130_fd_sc_hd__buf_2 wire2290 (.A(net2291),
    .X(net2290));
 sky130_fd_sc_hd__clkbuf_2 wire2291 (.A(\mprj_logic1[436] ),
    .X(net2291));
 sky130_fd_sc_hd__clkbuf_2 wire2292 (.A(\mprj_logic1[435] ),
    .X(net2292));
 sky130_fd_sc_hd__clkbuf_2 wire2293 (.A(\mprj_logic1[434] ),
    .X(net2293));
 sky130_fd_sc_hd__clkbuf_2 wire2294 (.A(\mprj_logic1[432] ),
    .X(net2294));
 sky130_fd_sc_hd__clkbuf_2 wire2295 (.A(\mprj_logic1[430] ),
    .X(net2295));
 sky130_fd_sc_hd__clkbuf_2 wire2296 (.A(\mprj_logic1[429] ),
    .X(net2296));
 sky130_fd_sc_hd__clkbuf_2 wire2297 (.A(\mprj_logic1[428] ),
    .X(net2297));
 sky130_fd_sc_hd__clkbuf_2 wire2298 (.A(\mprj_logic1[427] ),
    .X(net2298));
 sky130_fd_sc_hd__clkbuf_2 wire2299 (.A(\mprj_logic1[426] ),
    .X(net2299));
 sky130_fd_sc_hd__clkbuf_2 wire2300 (.A(\mprj_logic1[425] ),
    .X(net2300));
 sky130_fd_sc_hd__clkbuf_2 wire2301 (.A(\mprj_logic1[424] ),
    .X(net2301));
 sky130_fd_sc_hd__clkbuf_2 wire2302 (.A(\mprj_logic1[423] ),
    .X(net2302));
 sky130_fd_sc_hd__clkbuf_2 wire2303 (.A(\mprj_logic1[422] ),
    .X(net2303));
 sky130_fd_sc_hd__clkbuf_2 wire2304 (.A(\mprj_logic1[421] ),
    .X(net2304));
 sky130_fd_sc_hd__clkbuf_2 wire2305 (.A(\mprj_logic1[419] ),
    .X(net2305));
 sky130_fd_sc_hd__clkbuf_2 wire2306 (.A(\mprj_logic1[418] ),
    .X(net2306));
 sky130_fd_sc_hd__buf_4 wire2307 (.A(net2308),
    .X(net2307));
 sky130_fd_sc_hd__clkbuf_2 wire2308 (.A(net2309),
    .X(net2308));
 sky130_fd_sc_hd__clkbuf_2 wire2309 (.A(\mprj_logic1[417] ),
    .X(net2309));
 sky130_fd_sc_hd__clkbuf_2 wire2310 (.A(\mprj_logic1[416] ),
    .X(net2310));
 sky130_fd_sc_hd__clkbuf_2 wire2311 (.A(\mprj_logic1[415] ),
    .X(net2311));
 sky130_fd_sc_hd__clkbuf_2 wire2312 (.A(\mprj_logic1[414] ),
    .X(net2312));
 sky130_fd_sc_hd__clkbuf_2 wire2313 (.A(\mprj_logic1[413] ),
    .X(net2313));
 sky130_fd_sc_hd__buf_2 wire2314 (.A(net2315),
    .X(net2314));
 sky130_fd_sc_hd__clkbuf_2 wire2315 (.A(net2316),
    .X(net2315));
 sky130_fd_sc_hd__clkbuf_2 wire2316 (.A(\mprj_logic1[410] ),
    .X(net2316));
 sky130_fd_sc_hd__clkbuf_2 wire2317 (.A(\mprj_logic1[409] ),
    .X(net2317));
 sky130_fd_sc_hd__clkbuf_2 wire2318 (.A(\mprj_logic1[408] ),
    .X(net2318));
 sky130_fd_sc_hd__clkbuf_2 wire2319 (.A(\mprj_logic1[407] ),
    .X(net2319));
 sky130_fd_sc_hd__clkbuf_2 wire2320 (.A(\mprj_logic1[406] ),
    .X(net2320));
 sky130_fd_sc_hd__buf_2 wire2321 (.A(net2322),
    .X(net2321));
 sky130_fd_sc_hd__clkbuf_2 wire2322 (.A(\mprj_logic1[405] ),
    .X(net2322));
 sky130_fd_sc_hd__clkbuf_2 wire2323 (.A(net2324),
    .X(net2323));
 sky130_fd_sc_hd__clkbuf_2 wire2324 (.A(\mprj_logic1[404] ),
    .X(net2324));
 sky130_fd_sc_hd__clkbuf_2 wire2325 (.A(net2326),
    .X(net2325));
 sky130_fd_sc_hd__clkbuf_2 wire2326 (.A(\mprj_logic1[403] ),
    .X(net2326));
 sky130_fd_sc_hd__clkbuf_2 wire2327 (.A(\mprj_logic1[402] ),
    .X(net2327));
 sky130_fd_sc_hd__clkbuf_2 wire2328 (.A(\mprj_logic1[401] ),
    .X(net2328));
 sky130_fd_sc_hd__clkbuf_2 wire2329 (.A(\mprj_logic1[400] ),
    .X(net2329));
 sky130_fd_sc_hd__clkbuf_2 wire2330 (.A(\mprj_logic1[391] ),
    .X(net2330));
 sky130_fd_sc_hd__clkbuf_2 wire2331 (.A(\mprj_logic1[390] ),
    .X(net2331));
 sky130_fd_sc_hd__clkbuf_2 wire2332 (.A(\mprj_logic1[387] ),
    .X(net2332));
 sky130_fd_sc_hd__clkbuf_2 wire2333 (.A(\mprj_logic1[386] ),
    .X(net2333));
 sky130_fd_sc_hd__clkbuf_2 wire2334 (.A(\mprj_logic1[384] ),
    .X(net2334));
 sky130_fd_sc_hd__clkbuf_2 wire2335 (.A(\mprj_logic1[383] ),
    .X(net2335));
 sky130_fd_sc_hd__clkbuf_2 wire2336 (.A(\mprj_logic1[382] ),
    .X(net2336));
 sky130_fd_sc_hd__clkbuf_2 wire2337 (.A(\mprj_logic1[381] ),
    .X(net2337));
 sky130_fd_sc_hd__clkbuf_2 wire2338 (.A(\mprj_logic1[380] ),
    .X(net2338));
 sky130_fd_sc_hd__clkbuf_2 wire2339 (.A(\mprj_logic1[378] ),
    .X(net2339));
 sky130_fd_sc_hd__clkbuf_2 wire2340 (.A(\mprj_logic1[377] ),
    .X(net2340));
 sky130_fd_sc_hd__clkbuf_2 wire2341 (.A(\mprj_logic1[376] ),
    .X(net2341));
 sky130_fd_sc_hd__clkbuf_2 wire2342 (.A(\mprj_logic1[375] ),
    .X(net2342));
 sky130_fd_sc_hd__clkbuf_2 wire2343 (.A(\mprj_logic1[374] ),
    .X(net2343));
 sky130_fd_sc_hd__clkbuf_2 wire2344 (.A(\mprj_logic1[373] ),
    .X(net2344));
 sky130_fd_sc_hd__clkbuf_2 wire2345 (.A(\mprj_logic1[372] ),
    .X(net2345));
 sky130_fd_sc_hd__clkbuf_2 wire2346 (.A(\mprj_logic1[371] ),
    .X(net2346));
 sky130_fd_sc_hd__clkbuf_2 wire2347 (.A(\mprj_logic1[370] ),
    .X(net2347));
 sky130_fd_sc_hd__clkbuf_2 wire2348 (.A(\mprj_logic1[369] ),
    .X(net2348));
 sky130_fd_sc_hd__clkbuf_2 wire2349 (.A(net2350),
    .X(net2349));
 sky130_fd_sc_hd__clkbuf_2 wire2350 (.A(\mprj_logic1[368] ),
    .X(net2350));
 sky130_fd_sc_hd__clkbuf_2 wire2351 (.A(\mprj_logic1[366] ),
    .X(net2351));
 sky130_fd_sc_hd__clkbuf_2 wire2352 (.A(net2353),
    .X(net2352));
 sky130_fd_sc_hd__clkbuf_2 wire2353 (.A(\mprj_logic1[365] ),
    .X(net2353));
 sky130_fd_sc_hd__clkbuf_2 wire2354 (.A(\mprj_logic1[364] ),
    .X(net2354));
 sky130_fd_sc_hd__clkbuf_2 wire2355 (.A(net2356),
    .X(net2355));
 sky130_fd_sc_hd__clkbuf_2 wire2356 (.A(\mprj_logic1[363] ),
    .X(net2356));
 sky130_fd_sc_hd__clkbuf_2 wire2357 (.A(\mprj_logic1[362] ),
    .X(net2357));
 sky130_fd_sc_hd__clkbuf_2 wire2358 (.A(\mprj_logic1[361] ),
    .X(net2358));
 sky130_fd_sc_hd__clkbuf_2 wire2359 (.A(net2360),
    .X(net2359));
 sky130_fd_sc_hd__clkbuf_2 wire2360 (.A(\mprj_logic1[360] ),
    .X(net2360));
 sky130_fd_sc_hd__clkbuf_2 wire2361 (.A(net2362),
    .X(net2361));
 sky130_fd_sc_hd__clkbuf_2 wire2362 (.A(\mprj_logic1[359] ),
    .X(net2362));
 sky130_fd_sc_hd__buf_2 wire2363 (.A(net2364),
    .X(net2363));
 sky130_fd_sc_hd__clkbuf_2 wire2364 (.A(\mprj_logic1[358] ),
    .X(net2364));
 sky130_fd_sc_hd__clkbuf_2 wire2365 (.A(\mprj_logic1[357] ),
    .X(net2365));
 sky130_fd_sc_hd__buf_2 wire2366 (.A(net2367),
    .X(net2366));
 sky130_fd_sc_hd__clkbuf_2 wire2367 (.A(\mprj_logic1[356] ),
    .X(net2367));
 sky130_fd_sc_hd__clkbuf_2 wire2368 (.A(net2369),
    .X(net2368));
 sky130_fd_sc_hd__clkbuf_2 wire2369 (.A(\mprj_logic1[355] ),
    .X(net2369));
 sky130_fd_sc_hd__clkbuf_2 wire2370 (.A(net2371),
    .X(net2370));
 sky130_fd_sc_hd__clkbuf_2 wire2371 (.A(\mprj_logic1[354] ),
    .X(net2371));
 sky130_fd_sc_hd__buf_2 wire2372 (.A(net2373),
    .X(net2372));
 sky130_fd_sc_hd__clkbuf_2 wire2373 (.A(net2374),
    .X(net2373));
 sky130_fd_sc_hd__clkbuf_2 wire2374 (.A(\mprj_logic1[353] ),
    .X(net2374));
 sky130_fd_sc_hd__buf_2 wire2375 (.A(net2376),
    .X(net2375));
 sky130_fd_sc_hd__clkbuf_2 wire2376 (.A(\mprj_logic1[352] ),
    .X(net2376));
 sky130_fd_sc_hd__clkbuf_2 wire2377 (.A(\mprj_logic1[351] ),
    .X(net2377));
 sky130_fd_sc_hd__buf_2 wire2378 (.A(net2379),
    .X(net2378));
 sky130_fd_sc_hd__clkbuf_2 wire2379 (.A(\mprj_logic1[350] ),
    .X(net2379));
 sky130_fd_sc_hd__buf_2 wire2380 (.A(net2381),
    .X(net2380));
 sky130_fd_sc_hd__clkbuf_2 wire2381 (.A(\mprj_logic1[349] ),
    .X(net2381));
 sky130_fd_sc_hd__buf_2 wire2382 (.A(net2383),
    .X(net2382));
 sky130_fd_sc_hd__clkbuf_2 wire2383 (.A(\mprj_logic1[348] ),
    .X(net2383));
 sky130_fd_sc_hd__clkbuf_2 wire2384 (.A(net2385),
    .X(net2384));
 sky130_fd_sc_hd__clkbuf_2 wire2385 (.A(\mprj_logic1[347] ),
    .X(net2385));
 sky130_fd_sc_hd__clkbuf_2 wire2386 (.A(net2387),
    .X(net2386));
 sky130_fd_sc_hd__clkbuf_2 wire2387 (.A(\mprj_logic1[346] ),
    .X(net2387));
 sky130_fd_sc_hd__buf_2 wire2388 (.A(net2389),
    .X(net2388));
 sky130_fd_sc_hd__clkbuf_2 wire2389 (.A(\mprj_logic1[345] ),
    .X(net2389));
 sky130_fd_sc_hd__buf_2 wire2390 (.A(net2391),
    .X(net2390));
 sky130_fd_sc_hd__clkbuf_2 wire2391 (.A(\mprj_logic1[344] ),
    .X(net2391));
 sky130_fd_sc_hd__buf_6 wire2392 (.A(net2393),
    .X(net2392));
 sky130_fd_sc_hd__buf_4 wire2393 (.A(net2394),
    .X(net2393));
 sky130_fd_sc_hd__clkbuf_2 wire2394 (.A(net2395),
    .X(net2394));
 sky130_fd_sc_hd__clkbuf_2 wire2395 (.A(\mprj_logic1[343] ),
    .X(net2395));
 sky130_fd_sc_hd__buf_2 wire2396 (.A(net2397),
    .X(net2396));
 sky130_fd_sc_hd__clkbuf_2 wire2397 (.A(net2398),
    .X(net2397));
 sky130_fd_sc_hd__clkbuf_2 wire2398 (.A(\mprj_logic1[342] ),
    .X(net2398));
 sky130_fd_sc_hd__buf_2 wire2399 (.A(net2400),
    .X(net2399));
 sky130_fd_sc_hd__clkbuf_2 wire2400 (.A(net2401),
    .X(net2400));
 sky130_fd_sc_hd__clkbuf_2 wire2401 (.A(\mprj_logic1[341] ),
    .X(net2401));
 sky130_fd_sc_hd__clkbuf_2 wire2402 (.A(\mprj_logic1[340] ),
    .X(net2402));
 sky130_fd_sc_hd__clkbuf_2 wire2403 (.A(\mprj_logic1[339] ),
    .X(net2403));
 sky130_fd_sc_hd__clkbuf_2 wire2404 (.A(\mprj_logic1[338] ),
    .X(net2404));
 sky130_fd_sc_hd__buf_2 wire2405 (.A(net2406),
    .X(net2405));
 sky130_fd_sc_hd__clkbuf_2 wire2406 (.A(\mprj_logic1[337] ),
    .X(net2406));
 sky130_fd_sc_hd__clkbuf_2 wire2407 (.A(\mprj_logic1[336] ),
    .X(net2407));
 sky130_fd_sc_hd__clkbuf_2 wire2408 (.A(net2409),
    .X(net2408));
 sky130_fd_sc_hd__clkbuf_2 wire2409 (.A(\mprj_logic1[335] ),
    .X(net2409));
 sky130_fd_sc_hd__buf_2 wire2410 (.A(net2411),
    .X(net2410));
 sky130_fd_sc_hd__clkbuf_2 wire2411 (.A(net2412),
    .X(net2411));
 sky130_fd_sc_hd__clkbuf_2 wire2412 (.A(\mprj_logic1[334] ),
    .X(net2412));
 sky130_fd_sc_hd__buf_2 wire2413 (.A(net2414),
    .X(net2413));
 sky130_fd_sc_hd__clkbuf_2 wire2414 (.A(\mprj_logic1[333] ),
    .X(net2414));
 sky130_fd_sc_hd__buf_2 wire2415 (.A(net2416),
    .X(net2415));
 sky130_fd_sc_hd__clkbuf_2 wire2416 (.A(\mprj_logic1[332] ),
    .X(net2416));
 sky130_fd_sc_hd__buf_6 wire2417 (.A(net2418),
    .X(net2417));
 sky130_fd_sc_hd__buf_4 wire2418 (.A(net2419),
    .X(net2418));
 sky130_fd_sc_hd__clkbuf_2 wire2419 (.A(\mprj_logic1[331] ),
    .X(net2419));
 sky130_fd_sc_hd__buf_2 wire2420 (.A(net2421),
    .X(net2420));
 sky130_fd_sc_hd__clkbuf_2 wire2421 (.A(\mprj_logic1[330] ),
    .X(net2421));
 sky130_fd_sc_hd__buf_6 wire2422 (.A(net2423),
    .X(net2422));
 sky130_fd_sc_hd__buf_6 wire2423 (.A(net2424),
    .X(net2423));
 sky130_fd_sc_hd__buf_4 wire2424 (.A(net2425),
    .X(net2424));
 sky130_fd_sc_hd__clkbuf_2 wire2425 (.A(net2426),
    .X(net2425));
 sky130_fd_sc_hd__clkbuf_2 wire2426 (.A(\mprj_logic1[329] ),
    .X(net2426));
 sky130_fd_sc_hd__buf_6 wire2427 (.A(net2428),
    .X(net2427));
 sky130_fd_sc_hd__buf_6 wire2428 (.A(net2429),
    .X(net2428));
 sky130_fd_sc_hd__buf_4 wire2429 (.A(net2430),
    .X(net2429));
 sky130_fd_sc_hd__clkbuf_2 wire2430 (.A(\mprj_logic1[328] ),
    .X(net2430));
 sky130_fd_sc_hd__buf_6 wire2431 (.A(net2432),
    .X(net2431));
 sky130_fd_sc_hd__buf_6 wire2432 (.A(net2433),
    .X(net2432));
 sky130_fd_sc_hd__buf_4 wire2433 (.A(net2434),
    .X(net2433));
 sky130_fd_sc_hd__clkbuf_2 wire2434 (.A(\mprj_logic1[327] ),
    .X(net2434));
 sky130_fd_sc_hd__buf_6 wire2435 (.A(net2436),
    .X(net2435));
 sky130_fd_sc_hd__buf_4 wire2436 (.A(net2437),
    .X(net2436));
 sky130_fd_sc_hd__clkbuf_2 wire2437 (.A(net2438),
    .X(net2437));
 sky130_fd_sc_hd__clkbuf_2 wire2438 (.A(\mprj_logic1[326] ),
    .X(net2438));
 sky130_fd_sc_hd__buf_6 wire2439 (.A(net2440),
    .X(net2439));
 sky130_fd_sc_hd__buf_6 wire2440 (.A(net2441),
    .X(net2440));
 sky130_fd_sc_hd__buf_4 wire2441 (.A(net2442),
    .X(net2441));
 sky130_fd_sc_hd__clkbuf_2 wire2442 (.A(\mprj_logic1[325] ),
    .X(net2442));
 sky130_fd_sc_hd__buf_6 wire2443 (.A(net2444),
    .X(net2443));
 sky130_fd_sc_hd__buf_6 wire2444 (.A(net2445),
    .X(net2444));
 sky130_fd_sc_hd__buf_4 wire2445 (.A(net2446),
    .X(net2445));
 sky130_fd_sc_hd__clkbuf_2 wire2446 (.A(\mprj_logic1[324] ),
    .X(net2446));
 sky130_fd_sc_hd__buf_6 wire2447 (.A(net2448),
    .X(net2447));
 sky130_fd_sc_hd__buf_4 wire2448 (.A(net2449),
    .X(net2448));
 sky130_fd_sc_hd__clkbuf_2 wire2449 (.A(net2450),
    .X(net2449));
 sky130_fd_sc_hd__clkbuf_2 wire2450 (.A(\mprj_logic1[323] ),
    .X(net2450));
 sky130_fd_sc_hd__buf_6 wire2451 (.A(net2452),
    .X(net2451));
 sky130_fd_sc_hd__buf_6 wire2452 (.A(net2453),
    .X(net2452));
 sky130_fd_sc_hd__buf_4 wire2453 (.A(net2454),
    .X(net2453));
 sky130_fd_sc_hd__clkbuf_2 wire2454 (.A(\mprj_logic1[322] ),
    .X(net2454));
 sky130_fd_sc_hd__buf_6 wire2455 (.A(net2456),
    .X(net2455));
 sky130_fd_sc_hd__buf_6 wire2456 (.A(net2457),
    .X(net2456));
 sky130_fd_sc_hd__buf_4 wire2457 (.A(net2458),
    .X(net2457));
 sky130_fd_sc_hd__clkbuf_2 wire2458 (.A(\mprj_logic1[321] ),
    .X(net2458));
 sky130_fd_sc_hd__buf_6 wire2459 (.A(net2460),
    .X(net2459));
 sky130_fd_sc_hd__buf_4 wire2460 (.A(net2461),
    .X(net2460));
 sky130_fd_sc_hd__clkbuf_2 wire2461 (.A(\mprj_logic1[320] ),
    .X(net2461));
 sky130_fd_sc_hd__clkbuf_2 wire2462 (.A(\mprj_logic1[31] ),
    .X(net2462));
 sky130_fd_sc_hd__buf_6 wire2463 (.A(net2464),
    .X(net2463));
 sky130_fd_sc_hd__buf_4 wire2464 (.A(net2465),
    .X(net2464));
 sky130_fd_sc_hd__clkbuf_2 wire2465 (.A(\mprj_logic1[319] ),
    .X(net2465));
 sky130_fd_sc_hd__buf_6 wire2466 (.A(net2467),
    .X(net2466));
 sky130_fd_sc_hd__buf_4 wire2467 (.A(net2468),
    .X(net2467));
 sky130_fd_sc_hd__clkbuf_2 wire2468 (.A(\mprj_logic1[318] ),
    .X(net2468));
 sky130_fd_sc_hd__buf_6 wire2469 (.A(net2470),
    .X(net2469));
 sky130_fd_sc_hd__buf_4 wire2470 (.A(net2471),
    .X(net2470));
 sky130_fd_sc_hd__clkbuf_2 wire2471 (.A(net2472),
    .X(net2471));
 sky130_fd_sc_hd__clkbuf_2 wire2472 (.A(\mprj_logic1[317] ),
    .X(net2472));
 sky130_fd_sc_hd__buf_6 wire2473 (.A(net2474),
    .X(net2473));
 sky130_fd_sc_hd__buf_6 wire2474 (.A(net2475),
    .X(net2474));
 sky130_fd_sc_hd__buf_4 wire2475 (.A(net2476),
    .X(net2475));
 sky130_fd_sc_hd__clkbuf_2 wire2476 (.A(\mprj_logic1[316] ),
    .X(net2476));
 sky130_fd_sc_hd__buf_2 wire2477 (.A(net2478),
    .X(net2477));
 sky130_fd_sc_hd__clkbuf_2 wire2478 (.A(net2479),
    .X(net2478));
 sky130_fd_sc_hd__clkbuf_2 wire2479 (.A(\mprj_logic1[315] ),
    .X(net2479));
 sky130_fd_sc_hd__buf_2 wire2480 (.A(net2481),
    .X(net2480));
 sky130_fd_sc_hd__clkbuf_2 wire2481 (.A(\mprj_logic1[314] ),
    .X(net2481));
 sky130_fd_sc_hd__buf_2 wire2482 (.A(net2483),
    .X(net2482));
 sky130_fd_sc_hd__clkbuf_2 wire2483 (.A(net2484),
    .X(net2483));
 sky130_fd_sc_hd__clkbuf_2 wire2484 (.A(\mprj_logic1[313] ),
    .X(net2484));
 sky130_fd_sc_hd__buf_6 wire2485 (.A(net2486),
    .X(net2485));
 sky130_fd_sc_hd__buf_6 wire2486 (.A(net2487),
    .X(net2486));
 sky130_fd_sc_hd__buf_4 wire2487 (.A(net2488),
    .X(net2487));
 sky130_fd_sc_hd__clkbuf_2 wire2488 (.A(\mprj_logic1[312] ),
    .X(net2488));
 sky130_fd_sc_hd__buf_6 wire2489 (.A(net2490),
    .X(net2489));
 sky130_fd_sc_hd__buf_4 wire2490 (.A(net2491),
    .X(net2490));
 sky130_fd_sc_hd__clkbuf_2 wire2491 (.A(\mprj_logic1[311] ),
    .X(net2491));
 sky130_fd_sc_hd__buf_6 wire2492 (.A(net2493),
    .X(net2492));
 sky130_fd_sc_hd__buf_4 wire2493 (.A(net2494),
    .X(net2493));
 sky130_fd_sc_hd__clkbuf_2 wire2494 (.A(\mprj_logic1[310] ),
    .X(net2494));
 sky130_fd_sc_hd__buf_6 wire2495 (.A(net2496),
    .X(net2495));
 sky130_fd_sc_hd__buf_4 wire2496 (.A(net2497),
    .X(net2496));
 sky130_fd_sc_hd__clkbuf_2 wire2497 (.A(\mprj_logic1[309] ),
    .X(net2497));
 sky130_fd_sc_hd__buf_4 wire2498 (.A(net2499),
    .X(net2498));
 sky130_fd_sc_hd__clkbuf_2 wire2499 (.A(net2500),
    .X(net2499));
 sky130_fd_sc_hd__clkbuf_2 wire2500 (.A(\mprj_logic1[308] ),
    .X(net2500));
 sky130_fd_sc_hd__buf_2 wire2501 (.A(net2502),
    .X(net2501));
 sky130_fd_sc_hd__clkbuf_2 wire2502 (.A(net2503),
    .X(net2502));
 sky130_fd_sc_hd__clkbuf_2 wire2503 (.A(\mprj_logic1[307] ),
    .X(net2503));
 sky130_fd_sc_hd__buf_2 wire2504 (.A(net2505),
    .X(net2504));
 sky130_fd_sc_hd__clkbuf_2 wire2505 (.A(\mprj_logic1[306] ),
    .X(net2505));
 sky130_fd_sc_hd__buf_2 wire2506 (.A(net2507),
    .X(net2506));
 sky130_fd_sc_hd__clkbuf_2 wire2507 (.A(net2508),
    .X(net2507));
 sky130_fd_sc_hd__clkbuf_2 wire2508 (.A(\mprj_logic1[305] ),
    .X(net2508));
 sky130_fd_sc_hd__buf_6 wire2509 (.A(net2510),
    .X(net2509));
 sky130_fd_sc_hd__buf_4 wire2510 (.A(net2511),
    .X(net2510));
 sky130_fd_sc_hd__clkbuf_2 wire2511 (.A(\mprj_logic1[304] ),
    .X(net2511));
 sky130_fd_sc_hd__buf_6 wire2512 (.A(net2513),
    .X(net2512));
 sky130_fd_sc_hd__buf_4 wire2513 (.A(net2514),
    .X(net2513));
 sky130_fd_sc_hd__clkbuf_2 wire2514 (.A(\mprj_logic1[303] ),
    .X(net2514));
 sky130_fd_sc_hd__buf_6 wire2515 (.A(net2516),
    .X(net2515));
 sky130_fd_sc_hd__buf_4 wire2516 (.A(net2517),
    .X(net2516));
 sky130_fd_sc_hd__clkbuf_2 wire2517 (.A(\mprj_logic1[302] ),
    .X(net2517));
 sky130_fd_sc_hd__buf_2 wire2518 (.A(net2519),
    .X(net2518));
 sky130_fd_sc_hd__clkbuf_2 wire2519 (.A(net2520),
    .X(net2519));
 sky130_fd_sc_hd__clkbuf_2 wire2520 (.A(\mprj_logic1[301] ),
    .X(net2520));
 sky130_fd_sc_hd__buf_2 wire2521 (.A(net2522),
    .X(net2521));
 sky130_fd_sc_hd__clkbuf_2 wire2522 (.A(net2523),
    .X(net2522));
 sky130_fd_sc_hd__clkbuf_2 wire2523 (.A(\mprj_logic1[300] ),
    .X(net2523));
 sky130_fd_sc_hd__buf_6 wire2524 (.A(net2525),
    .X(net2524));
 sky130_fd_sc_hd__buf_6 wire2525 (.A(net2526),
    .X(net2525));
 sky130_fd_sc_hd__buf_4 wire2526 (.A(net2527),
    .X(net2526));
 sky130_fd_sc_hd__clkbuf_2 wire2527 (.A(net2528),
    .X(net2527));
 sky130_fd_sc_hd__clkbuf_2 wire2528 (.A(\mprj_logic1[2] ),
    .X(net2528));
 sky130_fd_sc_hd__buf_2 wire2529 (.A(net2530),
    .X(net2529));
 sky130_fd_sc_hd__clkbuf_2 wire2530 (.A(\mprj_logic1[299] ),
    .X(net2530));
 sky130_fd_sc_hd__buf_2 wire2531 (.A(net2532),
    .X(net2531));
 sky130_fd_sc_hd__clkbuf_2 wire2532 (.A(net2533),
    .X(net2532));
 sky130_fd_sc_hd__clkbuf_2 wire2533 (.A(\mprj_logic1[298] ),
    .X(net2533));
 sky130_fd_sc_hd__buf_6 wire2534 (.A(net2535),
    .X(net2534));
 sky130_fd_sc_hd__buf_4 wire2535 (.A(net2536),
    .X(net2535));
 sky130_fd_sc_hd__clkbuf_2 wire2536 (.A(\mprj_logic1[297] ),
    .X(net2536));
 sky130_fd_sc_hd__buf_2 wire2537 (.A(net2538),
    .X(net2537));
 sky130_fd_sc_hd__clkbuf_2 wire2538 (.A(\mprj_logic1[296] ),
    .X(net2538));
 sky130_fd_sc_hd__clkbuf_2 wire2539 (.A(net2540),
    .X(net2539));
 sky130_fd_sc_hd__clkbuf_2 wire2540 (.A(\mprj_logic1[295] ),
    .X(net2540));
 sky130_fd_sc_hd__clkbuf_2 wire2541 (.A(\mprj_logic1[293] ),
    .X(net2541));
 sky130_fd_sc_hd__clkbuf_2 wire2542 (.A(\mprj_logic1[292] ),
    .X(net2542));
 sky130_fd_sc_hd__clkbuf_2 wire2543 (.A(\mprj_logic1[291] ),
    .X(net2543));
 sky130_fd_sc_hd__buf_6 wire2544 (.A(net2545),
    .X(net2544));
 sky130_fd_sc_hd__buf_4 wire2545 (.A(net2546),
    .X(net2545));
 sky130_fd_sc_hd__clkbuf_2 wire2546 (.A(\mprj_logic1[290] ),
    .X(net2546));
 sky130_fd_sc_hd__clkbuf_2 wire2547 (.A(\mprj_logic1[28] ),
    .X(net2547));
 sky130_fd_sc_hd__buf_6 wire2548 (.A(net2549),
    .X(net2548));
 sky130_fd_sc_hd__buf_4 wire2549 (.A(net2550),
    .X(net2549));
 sky130_fd_sc_hd__clkbuf_2 wire2550 (.A(\mprj_logic1[289] ),
    .X(net2550));
 sky130_fd_sc_hd__buf_6 wire2551 (.A(net2552),
    .X(net2551));
 sky130_fd_sc_hd__buf_4 wire2552 (.A(net2553),
    .X(net2552));
 sky130_fd_sc_hd__clkbuf_2 wire2553 (.A(net2554),
    .X(net2553));
 sky130_fd_sc_hd__clkbuf_2 wire2554 (.A(\mprj_logic1[288] ),
    .X(net2554));
 sky130_fd_sc_hd__buf_2 wire2555 (.A(net2556),
    .X(net2555));
 sky130_fd_sc_hd__clkbuf_2 wire2556 (.A(net2557),
    .X(net2556));
 sky130_fd_sc_hd__clkbuf_2 wire2557 (.A(\mprj_logic1[287] ),
    .X(net2557));
 sky130_fd_sc_hd__buf_6 wire2558 (.A(net2559),
    .X(net2558));
 sky130_fd_sc_hd__buf_4 wire2559 (.A(net2560),
    .X(net2559));
 sky130_fd_sc_hd__clkbuf_2 wire2560 (.A(\mprj_logic1[286] ),
    .X(net2560));
 sky130_fd_sc_hd__buf_6 wire2561 (.A(net2562),
    .X(net2561));
 sky130_fd_sc_hd__buf_4 wire2562 (.A(net2563),
    .X(net2562));
 sky130_fd_sc_hd__clkbuf_2 wire2563 (.A(\mprj_logic1[285] ),
    .X(net2563));
 sky130_fd_sc_hd__buf_6 wire2564 (.A(net2565),
    .X(net2564));
 sky130_fd_sc_hd__buf_4 wire2565 (.A(net2566),
    .X(net2565));
 sky130_fd_sc_hd__clkbuf_2 wire2566 (.A(net2567),
    .X(net2566));
 sky130_fd_sc_hd__clkbuf_2 wire2567 (.A(\mprj_logic1[284] ),
    .X(net2567));
 sky130_fd_sc_hd__buf_2 wire2568 (.A(net2569),
    .X(net2568));
 sky130_fd_sc_hd__clkbuf_2 wire2569 (.A(\mprj_logic1[283] ),
    .X(net2569));
 sky130_fd_sc_hd__buf_6 wire2570 (.A(net2571),
    .X(net2570));
 sky130_fd_sc_hd__buf_4 wire2571 (.A(net2572),
    .X(net2571));
 sky130_fd_sc_hd__clkbuf_2 wire2572 (.A(\mprj_logic1[282] ),
    .X(net2572));
 sky130_fd_sc_hd__buf_2 wire2573 (.A(net2574),
    .X(net2573));
 sky130_fd_sc_hd__clkbuf_2 wire2574 (.A(\mprj_logic1[281] ),
    .X(net2574));
 sky130_fd_sc_hd__buf_2 wire2575 (.A(net2576),
    .X(net2575));
 sky130_fd_sc_hd__clkbuf_2 wire2576 (.A(net2577),
    .X(net2576));
 sky130_fd_sc_hd__clkbuf_2 wire2577 (.A(\mprj_logic1[280] ),
    .X(net2577));
 sky130_fd_sc_hd__buf_2 wire2578 (.A(net2579),
    .X(net2578));
 sky130_fd_sc_hd__clkbuf_2 wire2579 (.A(net2580),
    .X(net2579));
 sky130_fd_sc_hd__clkbuf_2 wire2580 (.A(\mprj_logic1[279] ),
    .X(net2580));
 sky130_fd_sc_hd__buf_2 wire2581 (.A(net2582),
    .X(net2581));
 sky130_fd_sc_hd__clkbuf_2 wire2582 (.A(net2583),
    .X(net2582));
 sky130_fd_sc_hd__clkbuf_2 wire2583 (.A(\mprj_logic1[278] ),
    .X(net2583));
 sky130_fd_sc_hd__buf_2 wire2584 (.A(net2585),
    .X(net2584));
 sky130_fd_sc_hd__clkbuf_2 wire2585 (.A(\mprj_logic1[277] ),
    .X(net2585));
 sky130_fd_sc_hd__buf_2 wire2586 (.A(net2587),
    .X(net2586));
 sky130_fd_sc_hd__clkbuf_2 wire2587 (.A(\mprj_logic1[276] ),
    .X(net2587));
 sky130_fd_sc_hd__clkbuf_2 wire2588 (.A(\mprj_logic1[275] ),
    .X(net2588));
 sky130_fd_sc_hd__clkbuf_2 wire2589 (.A(net2590),
    .X(net2589));
 sky130_fd_sc_hd__clkbuf_2 wire2590 (.A(\mprj_logic1[274] ),
    .X(net2590));
 sky130_fd_sc_hd__clkbuf_2 wire2591 (.A(net2592),
    .X(net2591));
 sky130_fd_sc_hd__clkbuf_2 wire2592 (.A(\mprj_logic1[273] ),
    .X(net2592));
 sky130_fd_sc_hd__clkbuf_2 wire2593 (.A(\mprj_logic1[272] ),
    .X(net2593));
 sky130_fd_sc_hd__clkbuf_2 wire2594 (.A(\mprj_logic1[271] ),
    .X(net2594));
 sky130_fd_sc_hd__clkbuf_2 wire2595 (.A(net2596),
    .X(net2595));
 sky130_fd_sc_hd__clkbuf_2 wire2596 (.A(\mprj_logic1[270] ),
    .X(net2596));
 sky130_fd_sc_hd__clkbuf_2 wire2597 (.A(\mprj_logic1[26] ),
    .X(net2597));
 sky130_fd_sc_hd__clkbuf_2 wire2598 (.A(\mprj_logic1[268] ),
    .X(net2598));
 sky130_fd_sc_hd__clkbuf_2 wire2599 (.A(\mprj_logic1[266] ),
    .X(net2599));
 sky130_fd_sc_hd__clkbuf_2 wire2600 (.A(\mprj_logic1[261] ),
    .X(net2600));
 sky130_fd_sc_hd__clkbuf_2 wire2601 (.A(\mprj_logic1[259] ),
    .X(net2601));
 sky130_fd_sc_hd__clkbuf_2 wire2602 (.A(\mprj_logic1[257] ),
    .X(net2602));
 sky130_fd_sc_hd__clkbuf_2 wire2603 (.A(\mprj_logic1[255] ),
    .X(net2603));
 sky130_fd_sc_hd__clkbuf_2 wire2604 (.A(\mprj_logic1[254] ),
    .X(net2604));
 sky130_fd_sc_hd__clkbuf_2 wire2605 (.A(\mprj_logic1[252] ),
    .X(net2605));
 sky130_fd_sc_hd__clkbuf_2 wire2606 (.A(\mprj_logic1[250] ),
    .X(net2606));
 sky130_fd_sc_hd__clkbuf_2 wire2607 (.A(\mprj_logic1[248] ),
    .X(net2607));
 sky130_fd_sc_hd__clkbuf_2 wire2608 (.A(\mprj_logic1[243] ),
    .X(net2608));
 sky130_fd_sc_hd__clkbuf_2 wire2609 (.A(\mprj_logic1[238] ),
    .X(net2609));
 sky130_fd_sc_hd__clkbuf_2 wire2610 (.A(\mprj_logic1[236] ),
    .X(net2610));
 sky130_fd_sc_hd__clkbuf_2 wire2611 (.A(\mprj_logic1[235] ),
    .X(net2611));
 sky130_fd_sc_hd__clkbuf_2 wire2612 (.A(\mprj_logic1[234] ),
    .X(net2612));
 sky130_fd_sc_hd__clkbuf_2 wire2613 (.A(net2614),
    .X(net2613));
 sky130_fd_sc_hd__clkbuf_2 wire2614 (.A(\mprj_logic1[233] ),
    .X(net2614));
 sky130_fd_sc_hd__clkbuf_2 wire2615 (.A(\mprj_logic1[232] ),
    .X(net2615));
 sky130_fd_sc_hd__clkbuf_2 wire2616 (.A(\mprj_logic1[231] ),
    .X(net2616));
 sky130_fd_sc_hd__clkbuf_2 wire2617 (.A(\mprj_logic1[230] ),
    .X(net2617));
 sky130_fd_sc_hd__buf_2 wire2618 (.A(net2619),
    .X(net2618));
 sky130_fd_sc_hd__clkbuf_2 wire2619 (.A(\mprj_logic1[229] ),
    .X(net2619));
 sky130_fd_sc_hd__buf_2 wire2620 (.A(net2621),
    .X(net2620));
 sky130_fd_sc_hd__clkbuf_2 wire2621 (.A(\mprj_logic1[227] ),
    .X(net2621));
 sky130_fd_sc_hd__clkbuf_2 wire2622 (.A(\mprj_logic1[226] ),
    .X(net2622));
 sky130_fd_sc_hd__buf_2 wire2623 (.A(net2624),
    .X(net2623));
 sky130_fd_sc_hd__clkbuf_2 wire2624 (.A(net2625),
    .X(net2624));
 sky130_fd_sc_hd__clkbuf_2 wire2625 (.A(\mprj_logic1[225] ),
    .X(net2625));
 sky130_fd_sc_hd__clkbuf_2 wire2626 (.A(\mprj_logic1[224] ),
    .X(net2626));
 sky130_fd_sc_hd__clkbuf_2 wire2627 (.A(\mprj_logic1[223] ),
    .X(net2627));
 sky130_fd_sc_hd__buf_2 wire2628 (.A(net2629),
    .X(net2628));
 sky130_fd_sc_hd__clkbuf_2 wire2629 (.A(\mprj_logic1[222] ),
    .X(net2629));
 sky130_fd_sc_hd__clkbuf_2 wire2630 (.A(net2631),
    .X(net2630));
 sky130_fd_sc_hd__clkbuf_2 wire2631 (.A(\mprj_logic1[221] ),
    .X(net2631));
 sky130_fd_sc_hd__buf_2 wire2632 (.A(net2633),
    .X(net2632));
 sky130_fd_sc_hd__clkbuf_2 wire2633 (.A(net2634),
    .X(net2633));
 sky130_fd_sc_hd__clkbuf_2 wire2634 (.A(\mprj_logic1[220] ),
    .X(net2634));
 sky130_fd_sc_hd__clkbuf_2 wire2635 (.A(\mprj_logic1[21] ),
    .X(net2635));
 sky130_fd_sc_hd__buf_2 wire2636 (.A(net2637),
    .X(net2636));
 sky130_fd_sc_hd__clkbuf_2 wire2637 (.A(\mprj_logic1[219] ),
    .X(net2637));
 sky130_fd_sc_hd__buf_2 wire2638 (.A(net2639),
    .X(net2638));
 sky130_fd_sc_hd__clkbuf_2 wire2639 (.A(\mprj_logic1[218] ),
    .X(net2639));
 sky130_fd_sc_hd__clkbuf_2 wire2640 (.A(net2641),
    .X(net2640));
 sky130_fd_sc_hd__clkbuf_2 wire2641 (.A(\mprj_logic1[217] ),
    .X(net2641));
 sky130_fd_sc_hd__buf_2 wire2642 (.A(net2643),
    .X(net2642));
 sky130_fd_sc_hd__clkbuf_2 wire2643 (.A(net2644),
    .X(net2643));
 sky130_fd_sc_hd__clkbuf_2 wire2644 (.A(\mprj_logic1[216] ),
    .X(net2644));
 sky130_fd_sc_hd__buf_2 wire2645 (.A(net2646),
    .X(net2645));
 sky130_fd_sc_hd__clkbuf_2 wire2646 (.A(net2647),
    .X(net2646));
 sky130_fd_sc_hd__clkbuf_2 wire2647 (.A(\mprj_logic1[215] ),
    .X(net2647));
 sky130_fd_sc_hd__clkbuf_2 wire2648 (.A(\mprj_logic1[214] ),
    .X(net2648));
 sky130_fd_sc_hd__buf_2 wire2649 (.A(net2650),
    .X(net2649));
 sky130_fd_sc_hd__clkbuf_2 wire2650 (.A(\mprj_logic1[213] ),
    .X(net2650));
 sky130_fd_sc_hd__buf_2 wire2651 (.A(net2652),
    .X(net2651));
 sky130_fd_sc_hd__clkbuf_2 wire2652 (.A(net2653),
    .X(net2652));
 sky130_fd_sc_hd__clkbuf_2 wire2653 (.A(\mprj_logic1[212] ),
    .X(net2653));
 sky130_fd_sc_hd__buf_6 wire2654 (.A(net2655),
    .X(net2654));
 sky130_fd_sc_hd__buf_4 wire2655 (.A(net2656),
    .X(net2655));
 sky130_fd_sc_hd__clkbuf_2 wire2656 (.A(\mprj_logic1[211] ),
    .X(net2656));
 sky130_fd_sc_hd__buf_2 wire2657 (.A(net2658),
    .X(net2657));
 sky130_fd_sc_hd__clkbuf_2 wire2658 (.A(\mprj_logic1[210] ),
    .X(net2658));
 sky130_fd_sc_hd__buf_2 wire2659 (.A(net2660),
    .X(net2659));
 sky130_fd_sc_hd__clkbuf_2 wire2660 (.A(\mprj_logic1[209] ),
    .X(net2660));
 sky130_fd_sc_hd__buf_4 wire2661 (.A(net2662),
    .X(net2661));
 sky130_fd_sc_hd__clkbuf_2 wire2662 (.A(net2663),
    .X(net2662));
 sky130_fd_sc_hd__clkbuf_2 wire2663 (.A(\mprj_logic1[208] ),
    .X(net2663));
 sky130_fd_sc_hd__buf_6 wire2664 (.A(net2665),
    .X(net2664));
 sky130_fd_sc_hd__buf_4 wire2665 (.A(net2666),
    .X(net2665));
 sky130_fd_sc_hd__clkbuf_2 wire2666 (.A(\mprj_logic1[207] ),
    .X(net2666));
 sky130_fd_sc_hd__buf_2 wire2667 (.A(net2668),
    .X(net2667));
 sky130_fd_sc_hd__clkbuf_2 wire2668 (.A(\mprj_logic1[206] ),
    .X(net2668));
 sky130_fd_sc_hd__buf_6 wire2669 (.A(net2670),
    .X(net2669));
 sky130_fd_sc_hd__buf_4 wire2670 (.A(net2671),
    .X(net2670));
 sky130_fd_sc_hd__clkbuf_2 wire2671 (.A(\mprj_logic1[205] ),
    .X(net2671));
 sky130_fd_sc_hd__buf_6 wire2672 (.A(net2673),
    .X(net2672));
 sky130_fd_sc_hd__buf_4 wire2673 (.A(net2674),
    .X(net2673));
 sky130_fd_sc_hd__clkbuf_2 wire2674 (.A(\mprj_logic1[204] ),
    .X(net2674));
 sky130_fd_sc_hd__buf_6 wire2675 (.A(net2676),
    .X(net2675));
 sky130_fd_sc_hd__buf_4 wire2676 (.A(net2677),
    .X(net2676));
 sky130_fd_sc_hd__clkbuf_2 wire2677 (.A(\mprj_logic1[203] ),
    .X(net2677));
 sky130_fd_sc_hd__buf_2 wire2678 (.A(net2679),
    .X(net2678));
 sky130_fd_sc_hd__clkbuf_2 wire2679 (.A(\mprj_logic1[202] ),
    .X(net2679));
 sky130_fd_sc_hd__buf_6 wire2680 (.A(net2681),
    .X(net2680));
 sky130_fd_sc_hd__buf_4 wire2681 (.A(net2682),
    .X(net2681));
 sky130_fd_sc_hd__clkbuf_2 wire2682 (.A(\mprj_logic1[201] ),
    .X(net2682));
 sky130_fd_sc_hd__buf_6 wire2683 (.A(net2684),
    .X(net2683));
 sky130_fd_sc_hd__buf_6 wire2684 (.A(net2685),
    .X(net2684));
 sky130_fd_sc_hd__buf_4 wire2685 (.A(net2686),
    .X(net2685));
 sky130_fd_sc_hd__clkbuf_2 wire2686 (.A(\mprj_logic1[200] ),
    .X(net2686));
 sky130_fd_sc_hd__buf_6 wire2687 (.A(net2688),
    .X(net2687));
 sky130_fd_sc_hd__buf_4 wire2688 (.A(net2689),
    .X(net2688));
 sky130_fd_sc_hd__clkbuf_2 wire2689 (.A(net2690),
    .X(net2689));
 sky130_fd_sc_hd__clkbuf_2 wire2690 (.A(\mprj_logic1[199] ),
    .X(net2690));
 sky130_fd_sc_hd__buf_6 wire2691 (.A(net2692),
    .X(net2691));
 sky130_fd_sc_hd__buf_4 wire2692 (.A(net2693),
    .X(net2692));
 sky130_fd_sc_hd__clkbuf_2 wire2693 (.A(net2694),
    .X(net2693));
 sky130_fd_sc_hd__clkbuf_2 wire2694 (.A(\mprj_logic1[198] ),
    .X(net2694));
 sky130_fd_sc_hd__buf_6 wire2695 (.A(net2696),
    .X(net2695));
 sky130_fd_sc_hd__buf_4 wire2696 (.A(net2697),
    .X(net2696));
 sky130_fd_sc_hd__clkbuf_2 wire2697 (.A(\mprj_logic1[197] ),
    .X(net2697));
 sky130_fd_sc_hd__buf_4 wire2698 (.A(net2699),
    .X(net2698));
 sky130_fd_sc_hd__buf_4 wire2699 (.A(net2700),
    .X(net2699));
 sky130_fd_sc_hd__clkbuf_2 wire2700 (.A(\mprj_logic1[196] ),
    .X(net2700));
 sky130_fd_sc_hd__buf_6 wire2701 (.A(net2702),
    .X(net2701));
 sky130_fd_sc_hd__buf_6 wire2702 (.A(net2703),
    .X(net2702));
 sky130_fd_sc_hd__buf_4 wire2703 (.A(net2704),
    .X(net2703));
 sky130_fd_sc_hd__clkbuf_2 wire2704 (.A(\mprj_logic1[195] ),
    .X(net2704));
 sky130_fd_sc_hd__buf_2 wire2705 (.A(net2706),
    .X(net2705));
 sky130_fd_sc_hd__clkbuf_2 wire2706 (.A(net2707),
    .X(net2706));
 sky130_fd_sc_hd__clkbuf_2 wire2707 (.A(\mprj_logic1[194] ),
    .X(net2707));
 sky130_fd_sc_hd__buf_6 wire2708 (.A(net2709),
    .X(net2708));
 sky130_fd_sc_hd__buf_4 wire2709 (.A(net2710),
    .X(net2709));
 sky130_fd_sc_hd__clkbuf_2 wire2710 (.A(\mprj_logic1[193] ),
    .X(net2710));
 sky130_fd_sc_hd__buf_6 wire2711 (.A(net2712),
    .X(net2711));
 sky130_fd_sc_hd__buf_4 wire2712 (.A(net2713),
    .X(net2712));
 sky130_fd_sc_hd__clkbuf_2 wire2713 (.A(\mprj_logic1[192] ),
    .X(net2713));
 sky130_fd_sc_hd__buf_2 wire2714 (.A(net2715),
    .X(net2714));
 sky130_fd_sc_hd__clkbuf_2 wire2715 (.A(\mprj_logic1[191] ),
    .X(net2715));
 sky130_fd_sc_hd__buf_6 wire2716 (.A(net2717),
    .X(net2716));
 sky130_fd_sc_hd__buf_4 wire2717 (.A(net2718),
    .X(net2717));
 sky130_fd_sc_hd__clkbuf_2 wire2718 (.A(\mprj_logic1[190] ),
    .X(net2718));
 sky130_fd_sc_hd__buf_2 wire2719 (.A(net2720),
    .X(net2719));
 sky130_fd_sc_hd__clkbuf_2 wire2720 (.A(net2721),
    .X(net2720));
 sky130_fd_sc_hd__clkbuf_2 wire2721 (.A(\mprj_logic1[189] ),
    .X(net2721));
 sky130_fd_sc_hd__buf_2 wire2722 (.A(net2723),
    .X(net2722));
 sky130_fd_sc_hd__clkbuf_2 wire2723 (.A(net2724),
    .X(net2723));
 sky130_fd_sc_hd__clkbuf_2 wire2724 (.A(\mprj_logic1[188] ),
    .X(net2724));
 sky130_fd_sc_hd__buf_2 wire2725 (.A(net2726),
    .X(net2725));
 sky130_fd_sc_hd__clkbuf_2 wire2726 (.A(\mprj_logic1[187] ),
    .X(net2726));
 sky130_fd_sc_hd__buf_2 wire2727 (.A(net2728),
    .X(net2727));
 sky130_fd_sc_hd__clkbuf_2 wire2728 (.A(\mprj_logic1[186] ),
    .X(net2728));
 sky130_fd_sc_hd__buf_6 wire2729 (.A(net2730),
    .X(net2729));
 sky130_fd_sc_hd__buf_4 wire2730 (.A(net2731),
    .X(net2730));
 sky130_fd_sc_hd__clkbuf_2 wire2731 (.A(\mprj_logic1[185] ),
    .X(net2731));
 sky130_fd_sc_hd__buf_2 wire2732 (.A(net2733),
    .X(net2732));
 sky130_fd_sc_hd__clkbuf_2 wire2733 (.A(\mprj_logic1[184] ),
    .X(net2733));
 sky130_fd_sc_hd__buf_2 wire2734 (.A(net2735),
    .X(net2734));
 sky130_fd_sc_hd__clkbuf_2 wire2735 (.A(\mprj_logic1[183] ),
    .X(net2735));
 sky130_fd_sc_hd__buf_2 wire2736 (.A(net2737),
    .X(net2736));
 sky130_fd_sc_hd__clkbuf_2 wire2737 (.A(net2738),
    .X(net2737));
 sky130_fd_sc_hd__clkbuf_2 wire2738 (.A(\mprj_logic1[182] ),
    .X(net2738));
 sky130_fd_sc_hd__clkbuf_2 wire2739 (.A(net2740),
    .X(net2739));
 sky130_fd_sc_hd__clkbuf_2 wire2740 (.A(\mprj_logic1[181] ),
    .X(net2740));
 sky130_fd_sc_hd__clkbuf_2 wire2741 (.A(\mprj_logic1[180] ),
    .X(net2741));
 sky130_fd_sc_hd__clkbuf_2 wire2742 (.A(\mprj_logic1[17] ),
    .X(net2742));
 sky130_fd_sc_hd__clkbuf_2 wire2743 (.A(net2744),
    .X(net2743));
 sky130_fd_sc_hd__clkbuf_2 wire2744 (.A(\mprj_logic1[179] ),
    .X(net2744));
 sky130_fd_sc_hd__clkbuf_2 wire2745 (.A(\mprj_logic1[178] ),
    .X(net2745));
 sky130_fd_sc_hd__buf_2 wire2746 (.A(net2747),
    .X(net2746));
 sky130_fd_sc_hd__clkbuf_2 wire2747 (.A(\mprj_logic1[177] ),
    .X(net2747));
 sky130_fd_sc_hd__clkbuf_2 wire2748 (.A(net2749),
    .X(net2748));
 sky130_fd_sc_hd__clkbuf_2 wire2749 (.A(\mprj_logic1[176] ),
    .X(net2749));
 sky130_fd_sc_hd__clkbuf_2 wire2750 (.A(\mprj_logic1[175] ),
    .X(net2750));
 sky130_fd_sc_hd__clkbuf_2 wire2751 (.A(net2752),
    .X(net2751));
 sky130_fd_sc_hd__clkbuf_2 wire2752 (.A(\mprj_logic1[174] ),
    .X(net2752));
 sky130_fd_sc_hd__clkbuf_2 wire2753 (.A(\mprj_logic1[173] ),
    .X(net2753));
 sky130_fd_sc_hd__clkbuf_2 wire2754 (.A(\mprj_logic1[172] ),
    .X(net2754));
 sky130_fd_sc_hd__clkbuf_2 wire2755 (.A(\mprj_logic1[171] ),
    .X(net2755));
 sky130_fd_sc_hd__clkbuf_2 wire2756 (.A(\mprj_logic1[170] ),
    .X(net2756));
 sky130_fd_sc_hd__clkbuf_2 wire2757 (.A(net2758),
    .X(net2757));
 sky130_fd_sc_hd__clkbuf_2 wire2758 (.A(\mprj_logic1[169] ),
    .X(net2758));
 sky130_fd_sc_hd__clkbuf_2 wire2759 (.A(\mprj_logic1[168] ),
    .X(net2759));
 sky130_fd_sc_hd__clkbuf_2 wire2760 (.A(\mprj_logic1[166] ),
    .X(net2760));
 sky130_fd_sc_hd__clkbuf_2 wire2761 (.A(\mprj_logic1[165] ),
    .X(net2761));
 sky130_fd_sc_hd__clkbuf_2 wire2762 (.A(\mprj_logic1[164] ),
    .X(net2762));
 sky130_fd_sc_hd__clkbuf_2 wire2763 (.A(\mprj_logic1[163] ),
    .X(net2763));
 sky130_fd_sc_hd__buf_2 wire2764 (.A(net2765),
    .X(net2764));
 sky130_fd_sc_hd__clkbuf_2 wire2765 (.A(net2766),
    .X(net2765));
 sky130_fd_sc_hd__clkbuf_2 wire2766 (.A(\mprj_logic1[162] ),
    .X(net2766));
 sky130_fd_sc_hd__buf_6 wire2767 (.A(net2768),
    .X(net2767));
 sky130_fd_sc_hd__buf_6 wire2768 (.A(net2769),
    .X(net2768));
 sky130_fd_sc_hd__buf_4 wire2769 (.A(net2770),
    .X(net2769));
 sky130_fd_sc_hd__clkbuf_2 wire2770 (.A(net2771),
    .X(net2770));
 sky130_fd_sc_hd__clkbuf_2 wire2771 (.A(\mprj_logic1[161] ),
    .X(net2771));
 sky130_fd_sc_hd__buf_6 wire2772 (.A(net2773),
    .X(net2772));
 sky130_fd_sc_hd__buf_6 wire2773 (.A(net2774),
    .X(net2773));
 sky130_fd_sc_hd__buf_4 wire2774 (.A(net2775),
    .X(net2774));
 sky130_fd_sc_hd__clkbuf_2 wire2775 (.A(\mprj_logic1[160] ),
    .X(net2775));
 sky130_fd_sc_hd__buf_6 wire2776 (.A(net2777),
    .X(net2776));
 sky130_fd_sc_hd__buf_6 wire2777 (.A(net2778),
    .X(net2777));
 sky130_fd_sc_hd__buf_4 wire2778 (.A(net2779),
    .X(net2778));
 sky130_fd_sc_hd__clkbuf_2 wire2779 (.A(\mprj_logic1[159] ),
    .X(net2779));
 sky130_fd_sc_hd__buf_6 wire2780 (.A(net2781),
    .X(net2780));
 sky130_fd_sc_hd__buf_4 wire2781 (.A(net2782),
    .X(net2781));
 sky130_fd_sc_hd__clkbuf_2 wire2782 (.A(\mprj_logic1[158] ),
    .X(net2782));
 sky130_fd_sc_hd__buf_6 wire2783 (.A(net2784),
    .X(net2783));
 sky130_fd_sc_hd__buf_6 wire2784 (.A(net2785),
    .X(net2784));
 sky130_fd_sc_hd__buf_4 wire2785 (.A(net2786),
    .X(net2785));
 sky130_fd_sc_hd__clkbuf_2 wire2786 (.A(\mprj_logic1[157] ),
    .X(net2786));
 sky130_fd_sc_hd__buf_6 wire2787 (.A(net2788),
    .X(net2787));
 sky130_fd_sc_hd__buf_6 wire2788 (.A(net2789),
    .X(net2788));
 sky130_fd_sc_hd__buf_4 wire2789 (.A(net2790),
    .X(net2789));
 sky130_fd_sc_hd__clkbuf_2 wire2790 (.A(\mprj_logic1[156] ),
    .X(net2790));
 sky130_fd_sc_hd__buf_6 wire2791 (.A(net2792),
    .X(net2791));
 sky130_fd_sc_hd__buf_4 wire2792 (.A(net2793),
    .X(net2792));
 sky130_fd_sc_hd__clkbuf_2 wire2793 (.A(net2794),
    .X(net2793));
 sky130_fd_sc_hd__clkbuf_2 wire2794 (.A(\mprj_logic1[155] ),
    .X(net2794));
 sky130_fd_sc_hd__buf_6 wire2795 (.A(net2796),
    .X(net2795));
 sky130_fd_sc_hd__buf_4 wire2796 (.A(net2797),
    .X(net2796));
 sky130_fd_sc_hd__clkbuf_2 wire2797 (.A(net2798),
    .X(net2797));
 sky130_fd_sc_hd__clkbuf_2 wire2798 (.A(\mprj_logic1[154] ),
    .X(net2798));
 sky130_fd_sc_hd__clkbuf_2 wire2799 (.A(net2800),
    .X(net2799));
 sky130_fd_sc_hd__clkbuf_2 wire2800 (.A(\mprj_logic1[153] ),
    .X(net2800));
 sky130_fd_sc_hd__buf_6 wire2801 (.A(net2802),
    .X(net2801));
 sky130_fd_sc_hd__buf_4 wire2802 (.A(net2803),
    .X(net2802));
 sky130_fd_sc_hd__clkbuf_2 wire2803 (.A(\mprj_logic1[152] ),
    .X(net2803));
 sky130_fd_sc_hd__buf_6 wire2804 (.A(net2805),
    .X(net2804));
 sky130_fd_sc_hd__buf_4 wire2805 (.A(net2806),
    .X(net2805));
 sky130_fd_sc_hd__clkbuf_2 wire2806 (.A(\mprj_logic1[151] ),
    .X(net2806));
 sky130_fd_sc_hd__buf_6 wire2807 (.A(net2808),
    .X(net2807));
 sky130_fd_sc_hd__buf_4 wire2808 (.A(net2809),
    .X(net2808));
 sky130_fd_sc_hd__clkbuf_2 wire2809 (.A(\mprj_logic1[150] ),
    .X(net2809));
 sky130_fd_sc_hd__clkbuf_2 wire2810 (.A(\mprj_logic1[14] ),
    .X(net2810));
 sky130_fd_sc_hd__clkbuf_2 wire2811 (.A(net2812),
    .X(net2811));
 sky130_fd_sc_hd__clkbuf_2 wire2812 (.A(\mprj_logic1[149] ),
    .X(net2812));
 sky130_fd_sc_hd__buf_6 wire2813 (.A(net2814),
    .X(net2813));
 sky130_fd_sc_hd__buf_4 wire2814 (.A(net2815),
    .X(net2814));
 sky130_fd_sc_hd__clkbuf_2 wire2815 (.A(\mprj_logic1[148] ),
    .X(net2815));
 sky130_fd_sc_hd__clkbuf_2 wire2816 (.A(net2817),
    .X(net2816));
 sky130_fd_sc_hd__clkbuf_2 wire2817 (.A(\mprj_logic1[147] ),
    .X(net2817));
 sky130_fd_sc_hd__clkbuf_2 wire2818 (.A(net2819),
    .X(net2818));
 sky130_fd_sc_hd__clkbuf_2 wire2819 (.A(\mprj_logic1[146] ),
    .X(net2819));
 sky130_fd_sc_hd__buf_2 wire2820 (.A(net2821),
    .X(net2820));
 sky130_fd_sc_hd__clkbuf_2 wire2821 (.A(\mprj_logic1[145] ),
    .X(net2821));
 sky130_fd_sc_hd__buf_2 wire2822 (.A(net2823),
    .X(net2822));
 sky130_fd_sc_hd__clkbuf_2 wire2823 (.A(\mprj_logic1[144] ),
    .X(net2823));
 sky130_fd_sc_hd__clkbuf_2 wire2824 (.A(\mprj_logic1[143] ),
    .X(net2824));
 sky130_fd_sc_hd__clkbuf_2 wire2825 (.A(net2826),
    .X(net2825));
 sky130_fd_sc_hd__clkbuf_2 wire2826 (.A(\mprj_logic1[142] ),
    .X(net2826));
 sky130_fd_sc_hd__clkbuf_2 wire2827 (.A(\mprj_logic1[141] ),
    .X(net2827));
 sky130_fd_sc_hd__clkbuf_2 wire2828 (.A(\mprj_logic1[134] ),
    .X(net2828));
 sky130_fd_sc_hd__clkbuf_2 wire2829 (.A(\mprj_logic1[12] ),
    .X(net2829));
 sky130_fd_sc_hd__clkbuf_2 wire2830 (.A(\mprj_logic1[128] ),
    .X(net2830));
 sky130_fd_sc_hd__clkbuf_2 wire2831 (.A(\mprj_logic1[127] ),
    .X(net2831));
 sky130_fd_sc_hd__clkbuf_2 wire2832 (.A(\mprj_logic1[126] ),
    .X(net2832));
 sky130_fd_sc_hd__clkbuf_2 wire2833 (.A(\mprj_logic1[121] ),
    .X(net2833));
 sky130_fd_sc_hd__clkbuf_2 wire2834 (.A(\mprj_logic1[117] ),
    .X(net2834));
 sky130_fd_sc_hd__clkbuf_2 wire2835 (.A(\mprj_logic1[115] ),
    .X(net2835));
 sky130_fd_sc_hd__clkbuf_2 wire2836 (.A(\mprj_logic1[114] ),
    .X(net2836));
 sky130_fd_sc_hd__clkbuf_2 wire2837 (.A(\mprj_logic1[10] ),
    .X(net2837));
 sky130_fd_sc_hd__clkbuf_2 wire2838 (.A(\mprj_logic1[107] ),
    .X(net2838));
 sky130_fd_sc_hd__clkbuf_2 wire2839 (.A(\mprj_logic1[106] ),
    .X(net2839));
 sky130_fd_sc_hd__clkbuf_2 wire2840 (.A(\mprj_logic1[105] ),
    .X(net2840));
 sky130_fd_sc_hd__clkbuf_2 wire2841 (.A(\mprj_logic1[104] ),
    .X(net2841));
 sky130_fd_sc_hd__clkbuf_2 wire2842 (.A(net2843),
    .X(net2842));
 sky130_fd_sc_hd__clkbuf_2 wire2843 (.A(\mprj_logic1[103] ),
    .X(net2843));
 sky130_fd_sc_hd__clkbuf_2 wire2844 (.A(\mprj_logic1[102] ),
    .X(net2844));
 sky130_fd_sc_hd__clkbuf_2 wire2845 (.A(net2846),
    .X(net2845));
 sky130_fd_sc_hd__clkbuf_2 wire2846 (.A(\mprj_logic1[101] ),
    .X(net2846));
 sky130_fd_sc_hd__clkbuf_2 wire2847 (.A(\mprj_logic1[100] ),
    .X(net2847));
 sky130_fd_sc_hd__clkbuf_2 wire2848 (.A(net2849),
    .X(net2848));
 sky130_fd_sc_hd__clkbuf_2 wire2849 (.A(\mprj_logic1[0] ),
    .X(net2849));
 sky130_fd_sc_hd__buf_6 wire2850 (.A(net2851),
    .X(net2850));
 sky130_fd_sc_hd__buf_4 wire2851 (.A(net2852),
    .X(net2851));
 sky130_fd_sc_hd__buf_6 wire2852 (.A(net2853),
    .X(net2852));
 sky130_fd_sc_hd__buf_6 wire2853 (.A(net2854),
    .X(net2853));
 sky130_fd_sc_hd__buf_4 wire2854 (.A(net2855),
    .X(net2854));
 sky130_fd_sc_hd__clkbuf_2 wire2855 (.A(net953),
    .X(net2855));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__A (.DIODE(_0018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0658__A (.DIODE(_0024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0662__A (.DIODE(_0026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A (.DIODE(_0030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A (.DIODE(_0032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0676__A (.DIODE(_0033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0680__A (.DIODE(_0035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A (.DIODE(_0044_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0706__A (.DIODE(_0048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A (.DIODE(_0050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0718__A (.DIODE(_0054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A (.DIODE(_0060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__A (.DIODE(_0068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A (.DIODE(_0072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__A (.DIODE(_0073_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1628_A (.DIODE(_0075_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1626_A (.DIODE(_0076_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1620_A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1619_A (.DIODE(_0080_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1616_A (.DIODE(_0081_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1611_A (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1606_A (.DIODE(_0085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__A (.DIODE(_0086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1604_A (.DIODE(_0087_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1601_A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1599_A (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1593_A (.DIODE(_0091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1590_A (.DIODE(_0092_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1581_A (.DIODE(_0095_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1576_A (.DIODE(_0097_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1569_A (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1563_A (.DIODE(_0102_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1560_A (.DIODE(_0103_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1555_A (.DIODE(_0105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__A (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A (.DIODE(_0109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A (.DIODE(_0112_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1553_A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1552_A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0844__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__A (.DIODE(_0126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__A (.DIODE(_0132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A (.DIODE(_0133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1551_A (.DIODE(_0135_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1550_A (.DIODE(_0136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1549_A (.DIODE(_0137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1548_A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0894__A (.DIODE(_0142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0896__A (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__A (.DIODE(_0145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A (.DIODE(_0146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0904__A (.DIODE(_0147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(_0150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0912__A (.DIODE(_0151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__A (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A (.DIODE(_0154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0920__A (.DIODE(_0155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A (.DIODE(_0156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (.DIODE(_0158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0928__A (.DIODE(_0159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0932__A (.DIODE(_0161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0934__A (.DIODE(_0162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0936__A (.DIODE(_0163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A (.DIODE(_0164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A (.DIODE(_0165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0942__A (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1540_A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0972__A (.DIODE(_0181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1536_A (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1535_A (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1530_A (.DIODE(_0190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1525_A (.DIODE(_0193_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1524_A (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1523_A (.DIODE(_0195_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1522_A (.DIODE(_0196_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1521_A (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1519_A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1515_A (.DIODE(_0200_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1512_A (.DIODE(_0201_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1511_A (.DIODE(_0202_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1510_A (.DIODE(_0203_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1509_A (.DIODE(_0204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__A (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__A (.DIODE(_0207_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1508_A (.DIODE(_0212_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1505_A (.DIODE(_0215_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1504_A (.DIODE(_0216_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1501_A (.DIODE(_0219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1500_A (.DIODE(_0220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__A (.DIODE(_0221_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1498_A (.DIODE(_0222_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1497_A (.DIODE(_0223_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1495_A (.DIODE(_0225_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1492_A (.DIODE(_0227_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1490_A (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1489_A (.DIODE(_0230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__A (.DIODE(_0231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A (.DIODE(_0232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A (.DIODE(_0233_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1488_A (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__A (.DIODE(_0235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A (.DIODE(_0238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A (.DIODE(_0239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A (.DIODE(_0240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A (.DIODE(_0242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A (.DIODE(_0245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1484_A (.DIODE(_0246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1482_A (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1481_A (.DIODE(_0248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A (.DIODE(_0250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1477_A (.DIODE(_0252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1476_A (.DIODE(_0254_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1472_A (.DIODE(_0257_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1470_A (.DIODE(_0258_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1465_A (.DIODE(_0260_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1463_A (.DIODE(_0261_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1461_A (.DIODE(_0262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1459_A (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1452_A (.DIODE(_0266_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1450_A (.DIODE(_0267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1448_A (.DIODE(_0268_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1446_A (.DIODE(_0269_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1444_A (.DIODE(_0271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A (.DIODE(_0272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A (.DIODE(_0273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A (.DIODE(_0276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__A (.DIODE(_0278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__A (.DIODE(_0279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (.DIODE(_0283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A (.DIODE(_0284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A (.DIODE(_0289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A (.DIODE(_0290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__A (.DIODE(_0291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A (.DIODE(_0292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__A (.DIODE(_0293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A (.DIODE(_0294_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1439_A (.DIODE(_0297_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1431_A (.DIODE(_0300_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1429_A (.DIODE(_0301_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1427_A (.DIODE(_0302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A (.DIODE(_0304_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1423_A (.DIODE(_0306_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1421_A (.DIODE(_0307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__A (.DIODE(_0310_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1418_A (.DIODE(_0311_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1414_A (.DIODE(_0313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1413_A (.DIODE(_0314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__A (.DIODE(_0316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__A (.DIODE(_0318_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1410_A (.DIODE(_0319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__A (.DIODE(_0321_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1406_A (.DIODE(_0324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A (.DIODE(_0325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__A (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1405_A (.DIODE(_0327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A (.DIODE(_0328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__A (.DIODE(_0329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__A (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__A (.DIODE(_0332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__A (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A (.DIODE(_0334_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1404_A (.DIODE(_0335_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1403_A (.DIODE(_0336_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1401_A (.DIODE(_0338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1394_A (.DIODE(_0342_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1392_A (.DIODE(_0343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1391_A (.DIODE(_0344_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1390_A (.DIODE(_0345_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1389_A (.DIODE(_0346_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1387_A (.DIODE(_0347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1386_A (.DIODE(_0348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1385_A (.DIODE(_0349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1382_A (.DIODE(_0351_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1381_A (.DIODE(_0352_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1374_A (.DIODE(_0357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__A (.DIODE(_0359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1334__A (.DIODE(_0362_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1368_A (.DIODE(_0363_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1367_A (.DIODE(_0364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1366_A (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1365_A (.DIODE(_0366_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1364_A (.DIODE(_0367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__A (.DIODE(_0368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1362_A (.DIODE(_0370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__A (.DIODE(_0373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A (.DIODE(_0376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1366__A (.DIODE(_0378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A (.DIODE(_0381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__A (.DIODE(_0382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1354_A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__A (.DIODE(_0387_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1350_A (.DIODE(_0388_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1348_A (.DIODE(_0389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__A (.DIODE(_0390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1347_A (.DIODE(_0391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1394__A (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1343_A (.DIODE(_0394_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1341_A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A (.DIODE(_0397_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1338_A (.DIODE(_0398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__A (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__A (.DIODE(_0401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A (.DIODE(_0402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__A (.DIODE(_0403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1418__A (.DIODE(_0404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__A (.DIODE(_0405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__A (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1430__A (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1436__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__A (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1442__A (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1448__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1333_A (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1330_A (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1329_A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__A (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__A (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__A (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__A (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__A (.DIODE(_0458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (.DIODE(_0459_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(caravel_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(caravel_clk2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(caravel_rstn));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[100]_B  (.DIODE(\la_data_in_enable[100] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[101]_B  (.DIODE(\la_data_in_enable[101] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[103]_B  (.DIODE(\la_data_in_enable[103] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[104]_B  (.DIODE(\la_data_in_enable[104] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[12]_B  (.DIODE(\la_data_in_enable[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[55]_B  (.DIODE(\la_data_in_enable[55] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[56]_B  (.DIODE(\la_data_in_enable[56] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[57]_B  (.DIODE(\la_data_in_enable[57] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[58]_B  (.DIODE(\la_data_in_enable[58] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[59]_B  (.DIODE(\la_data_in_enable[59] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[60]_B  (.DIODE(\la_data_in_enable[60] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[71]_B  (.DIODE(\la_data_in_enable[71] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[75]_B  (.DIODE(\la_data_in_enable[75] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[84]_B  (.DIODE(\la_data_in_enable[84] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[88]_B  (.DIODE(\la_data_in_enable[88] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[93]_B  (.DIODE(\la_data_in_enable[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1086_A (.DIODE(\la_data_in_mprj_bar[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1083_A (.DIODE(\la_data_in_mprj_bar[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__A (.DIODE(\la_data_in_mprj_bar[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0552__A (.DIODE(\la_data_in_mprj_bar[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0553__A (.DIODE(\la_data_in_mprj_bar[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0555__A (.DIODE(\la_data_in_mprj_bar[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0557__A (.DIODE(\la_data_in_mprj_bar[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0562__A (.DIODE(\la_data_in_mprj_bar[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0568__A (.DIODE(\la_data_in_mprj_bar[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0474__A (.DIODE(\la_data_in_mprj_bar[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0476__A (.DIODE(\la_data_in_mprj_bar[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0477__A (.DIODE(\la_data_in_mprj_bar[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0479__A (.DIODE(\la_data_in_mprj_bar[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0481__A (.DIODE(\la_data_in_mprj_bar[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0484__A (.DIODE(\la_data_in_mprj_bar[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A (.DIODE(\la_data_in_mprj_bar[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0485__A (.DIODE(\la_data_in_mprj_bar[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0487__A (.DIODE(\la_data_in_mprj_bar[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0492__A (.DIODE(\la_data_in_mprj_bar[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0494__A (.DIODE(\la_data_in_mprj_bar[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0495__A (.DIODE(\la_data_in_mprj_bar[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0497__A (.DIODE(\la_data_in_mprj_bar[52] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0499__A (.DIODE(\la_data_in_mprj_bar[54] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0501__A (.DIODE(\la_data_in_mprj_bar[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0502__A (.DIODE(\la_data_in_mprj_bar[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0503__A (.DIODE(\la_data_in_mprj_bar[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0504__A (.DIODE(\la_data_in_mprj_bar[59] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0505__A (.DIODE(\la_data_in_mprj_bar[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0506__A (.DIODE(\la_data_in_mprj_bar[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0507__A (.DIODE(\la_data_in_mprj_bar[62] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0508__A (.DIODE(\la_data_in_mprj_bar[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0510__A (.DIODE(\la_data_in_mprj_bar[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0511__A (.DIODE(\la_data_in_mprj_bar[66] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0512__A (.DIODE(\la_data_in_mprj_bar[67] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0513__A (.DIODE(\la_data_in_mprj_bar[68] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0514__A (.DIODE(\la_data_in_mprj_bar[69] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1078_A (.DIODE(\la_data_in_mprj_bar[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1074_A (.DIODE(\la_data_in_mprj_bar[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1069_A (.DIODE(\la_data_in_mprj_bar[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1062_A (.DIODE(\la_data_in_mprj_bar[78] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1060_A (.DIODE(\la_data_in_mprj_bar[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1058_A (.DIODE(\la_data_in_mprj_bar[80] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1055_A (.DIODE(\la_data_in_mprj_bar[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1052_A (.DIODE(\la_data_in_mprj_bar[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1050_A (.DIODE(\la_data_in_mprj_bar[83] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1045_A (.DIODE(\la_data_in_mprj_bar[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1035_A (.DIODE(\la_data_in_mprj_bar[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1034_A (.DIODE(\la_data_in_mprj_bar[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1031_A (.DIODE(\la_data_in_mprj_bar[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1029_A (.DIODE(\la_data_in_mprj_bar[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1025_A (.DIODE(\la_data_in_mprj_bar[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1018_A (.DIODE(\la_data_in_mprj_bar[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1016_A (.DIODE(\la_data_in_mprj_bar[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1014_A (.DIODE(\la_data_in_mprj_bar[99] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[0]_A  (.DIODE(la_data_out_core[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[100]_A  (.DIODE(la_data_out_core[100]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[101]_A  (.DIODE(la_data_out_core[101]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[102]_A  (.DIODE(la_data_out_core[102]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[103]_A  (.DIODE(la_data_out_core[103]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[104]_A  (.DIODE(la_data_out_core[104]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[105]_A  (.DIODE(la_data_out_core[105]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[106]_A  (.DIODE(la_data_out_core[106]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[107]_A  (.DIODE(la_data_out_core[107]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[108]_A  (.DIODE(la_data_out_core[108]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[109]_A  (.DIODE(la_data_out_core[109]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[10]_A  (.DIODE(la_data_out_core[10]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[110]_A  (.DIODE(la_data_out_core[110]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[111]_A  (.DIODE(la_data_out_core[111]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[112]_A  (.DIODE(la_data_out_core[112]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[113]_A  (.DIODE(la_data_out_core[113]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[114]_A  (.DIODE(la_data_out_core[114]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[115]_A  (.DIODE(la_data_out_core[115]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[116]_A  (.DIODE(la_data_out_core[116]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[117]_A  (.DIODE(la_data_out_core[117]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[118]_A  (.DIODE(la_data_out_core[118]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[119]_A  (.DIODE(la_data_out_core[119]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[11]_A  (.DIODE(la_data_out_core[11]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[120]_A  (.DIODE(la_data_out_core[120]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[121]_A  (.DIODE(la_data_out_core[121]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[122]_A  (.DIODE(la_data_out_core[122]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[123]_A  (.DIODE(la_data_out_core[123]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[124]_A  (.DIODE(la_data_out_core[124]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[125]_A  (.DIODE(la_data_out_core[125]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[126]_A  (.DIODE(la_data_out_core[126]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[127]_A  (.DIODE(la_data_out_core[127]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[12]_A  (.DIODE(la_data_out_core[12]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[13]_A  (.DIODE(la_data_out_core[13]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[14]_A  (.DIODE(la_data_out_core[14]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[15]_A  (.DIODE(la_data_out_core[15]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[16]_A  (.DIODE(la_data_out_core[16]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[17]_A  (.DIODE(la_data_out_core[17]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[18]_A  (.DIODE(la_data_out_core[18]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[19]_A  (.DIODE(la_data_out_core[19]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[1]_A  (.DIODE(la_data_out_core[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[20]_A  (.DIODE(la_data_out_core[20]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[21]_A  (.DIODE(la_data_out_core[21]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[22]_A  (.DIODE(la_data_out_core[22]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[23]_A  (.DIODE(la_data_out_core[23]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[24]_A  (.DIODE(la_data_out_core[24]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[25]_A  (.DIODE(la_data_out_core[25]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[26]_A  (.DIODE(la_data_out_core[26]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[27]_A  (.DIODE(la_data_out_core[27]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[28]_A  (.DIODE(la_data_out_core[28]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[29]_A  (.DIODE(la_data_out_core[29]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[2]_A  (.DIODE(la_data_out_core[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[30]_A  (.DIODE(la_data_out_core[30]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[31]_A  (.DIODE(la_data_out_core[31]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[32]_A  (.DIODE(la_data_out_core[32]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[33]_A  (.DIODE(la_data_out_core[33]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[34]_A  (.DIODE(la_data_out_core[34]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[35]_A  (.DIODE(la_data_out_core[35]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[36]_A  (.DIODE(la_data_out_core[36]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[37]_A  (.DIODE(la_data_out_core[37]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[38]_A  (.DIODE(la_data_out_core[38]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[39]_A  (.DIODE(la_data_out_core[39]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[3]_A  (.DIODE(la_data_out_core[3]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[40]_A  (.DIODE(la_data_out_core[40]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[41]_A  (.DIODE(la_data_out_core[41]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[42]_A  (.DIODE(la_data_out_core[42]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[43]_A  (.DIODE(la_data_out_core[43]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[44]_A  (.DIODE(la_data_out_core[44]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[45]_A  (.DIODE(la_data_out_core[45]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[46]_A  (.DIODE(la_data_out_core[46]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[47]_A  (.DIODE(la_data_out_core[47]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[48]_A  (.DIODE(la_data_out_core[48]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[49]_A  (.DIODE(la_data_out_core[49]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[4]_A  (.DIODE(la_data_out_core[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[50]_A  (.DIODE(la_data_out_core[50]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[51]_A  (.DIODE(la_data_out_core[51]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[52]_A  (.DIODE(la_data_out_core[52]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[53]_A  (.DIODE(la_data_out_core[53]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[54]_A  (.DIODE(la_data_out_core[54]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[55]_A  (.DIODE(la_data_out_core[55]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[56]_A  (.DIODE(la_data_out_core[56]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[57]_A  (.DIODE(la_data_out_core[57]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[58]_A  (.DIODE(la_data_out_core[58]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[59]_A  (.DIODE(la_data_out_core[59]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[5]_A  (.DIODE(la_data_out_core[5]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[60]_A  (.DIODE(la_data_out_core[60]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[61]_A  (.DIODE(la_data_out_core[61]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[62]_A  (.DIODE(la_data_out_core[62]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[63]_A  (.DIODE(la_data_out_core[63]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[64]_A  (.DIODE(la_data_out_core[64]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[65]_A  (.DIODE(la_data_out_core[65]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[66]_A  (.DIODE(la_data_out_core[66]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[67]_A  (.DIODE(la_data_out_core[67]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[68]_A  (.DIODE(la_data_out_core[68]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[69]_A  (.DIODE(la_data_out_core[69]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[6]_A  (.DIODE(la_data_out_core[6]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[70]_A  (.DIODE(la_data_out_core[70]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[71]_A  (.DIODE(la_data_out_core[71]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[72]_A  (.DIODE(la_data_out_core[72]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[73]_A  (.DIODE(la_data_out_core[73]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[74]_A  (.DIODE(la_data_out_core[74]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[75]_A  (.DIODE(la_data_out_core[75]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[76]_A  (.DIODE(la_data_out_core[76]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[77]_A  (.DIODE(la_data_out_core[77]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[78]_A  (.DIODE(la_data_out_core[78]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[79]_A  (.DIODE(la_data_out_core[79]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[7]_A  (.DIODE(la_data_out_core[7]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[80]_A  (.DIODE(la_data_out_core[80]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[81]_A  (.DIODE(la_data_out_core[81]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[82]_A  (.DIODE(la_data_out_core[82]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[83]_A  (.DIODE(la_data_out_core[83]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[84]_A  (.DIODE(la_data_out_core[84]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[85]_A  (.DIODE(la_data_out_core[85]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[86]_A  (.DIODE(la_data_out_core[86]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[87]_A  (.DIODE(la_data_out_core[87]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[88]_A  (.DIODE(la_data_out_core[88]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[89]_A  (.DIODE(la_data_out_core[89]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[8]_A  (.DIODE(la_data_out_core[8]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[90]_A  (.DIODE(la_data_out_core[90]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[91]_A  (.DIODE(la_data_out_core[91]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[92]_A  (.DIODE(la_data_out_core[92]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[93]_A  (.DIODE(la_data_out_core[93]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[94]_A  (.DIODE(la_data_out_core[94]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[95]_A  (.DIODE(la_data_out_core[95]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[96]_A  (.DIODE(la_data_out_core[96]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[97]_A  (.DIODE(la_data_out_core[97]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[98]_A  (.DIODE(la_data_out_core[98]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[99]_A  (.DIODE(la_data_out_core[99]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[9]_A  (.DIODE(la_data_out_core[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(la_data_out_mprj[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(la_data_out_mprj[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(la_data_out_mprj[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(la_data_out_mprj[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(la_data_out_mprj[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(la_data_out_mprj[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(la_data_out_mprj[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(la_data_out_mprj[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(la_data_out_mprj[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(la_data_out_mprj[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(la_data_out_mprj[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(la_data_out_mprj[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(la_data_out_mprj[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(la_data_out_mprj[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(la_data_out_mprj[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(la_data_out_mprj[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(la_data_out_mprj[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(la_data_out_mprj[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(la_data_out_mprj[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(la_data_out_mprj[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(la_data_out_mprj[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(la_data_out_mprj[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(la_data_out_mprj[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(la_data_out_mprj[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(la_data_out_mprj[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(la_data_out_mprj[122]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(la_data_out_mprj[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(la_data_out_mprj[124]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(la_data_out_mprj[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(la_data_out_mprj[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(la_data_out_mprj[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(la_data_out_mprj[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(la_data_out_mprj[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(la_data_out_mprj[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(la_data_out_mprj[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(la_data_out_mprj[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(la_data_out_mprj[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(la_data_out_mprj[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(la_data_out_mprj[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(la_data_out_mprj[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(la_data_out_mprj[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(la_data_out_mprj[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(la_data_out_mprj[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(la_data_out_mprj[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(la_data_out_mprj[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(la_data_out_mprj[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(la_data_out_mprj[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(la_data_out_mprj[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(la_data_out_mprj[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(la_data_out_mprj[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(la_data_out_mprj[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(la_data_out_mprj[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(la_data_out_mprj[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(la_data_out_mprj[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(la_data_out_mprj[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(la_data_out_mprj[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(la_data_out_mprj[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(la_data_out_mprj[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(la_data_out_mprj[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(la_data_out_mprj[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(la_data_out_mprj[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(la_data_out_mprj[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(la_data_out_mprj[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(la_data_out_mprj[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(la_data_out_mprj[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(la_data_out_mprj[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(la_data_out_mprj[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(la_data_out_mprj[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(la_data_out_mprj[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(la_data_out_mprj[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(la_data_out_mprj[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(la_data_out_mprj[49]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(la_data_out_mprj[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(la_data_out_mprj[50]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(la_data_out_mprj[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(la_data_out_mprj[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(la_data_out_mprj[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(la_data_out_mprj[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(la_data_out_mprj[55]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(la_data_out_mprj[56]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(la_data_out_mprj[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(la_data_out_mprj[58]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(la_data_out_mprj[59]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(la_data_out_mprj[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(la_data_out_mprj[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(la_data_out_mprj[61]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(la_data_out_mprj[62]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(la_data_out_mprj[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(la_data_out_mprj[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(la_data_out_mprj[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(la_data_out_mprj[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(la_data_out_mprj[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(la_data_out_mprj[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(la_data_out_mprj[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(la_data_out_mprj[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(la_data_out_mprj[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(la_data_out_mprj[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(la_data_out_mprj[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(la_data_out_mprj[73]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(la_data_out_mprj[74]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(la_data_out_mprj[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(la_data_out_mprj[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(la_data_out_mprj[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(la_data_out_mprj[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(la_data_out_mprj[79]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(la_data_out_mprj[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(la_data_out_mprj[80]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(la_data_out_mprj[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(la_data_out_mprj[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(la_data_out_mprj[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(la_data_out_mprj[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(la_data_out_mprj[85]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(la_data_out_mprj[86]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(la_data_out_mprj[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(la_data_out_mprj[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(la_data_out_mprj[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(la_data_out_mprj[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(la_data_out_mprj[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(la_data_out_mprj[91]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(la_data_out_mprj[92]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(la_data_out_mprj[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(la_data_out_mprj[94]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(la_data_out_mprj[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(la_data_out_mprj[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(la_data_out_mprj[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(la_data_out_mprj[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(la_data_out_mprj[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(la_data_out_mprj[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(la_iena_mprj[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(la_iena_mprj[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(la_iena_mprj[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(la_iena_mprj[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(la_iena_mprj[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(la_iena_mprj[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(la_iena_mprj[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(la_iena_mprj[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(la_iena_mprj[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(la_iena_mprj[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(la_iena_mprj[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(la_iena_mprj[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(la_iena_mprj[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(la_iena_mprj[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(la_iena_mprj[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(la_iena_mprj[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(la_iena_mprj[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(la_iena_mprj[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(la_iena_mprj[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(la_iena_mprj[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(la_iena_mprj[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(la_iena_mprj[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(la_iena_mprj[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(la_iena_mprj[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(la_iena_mprj[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(la_iena_mprj[122]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(la_iena_mprj[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(la_iena_mprj[124]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(la_iena_mprj[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(la_iena_mprj[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(la_iena_mprj[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(la_iena_mprj[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(la_iena_mprj[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(la_iena_mprj[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(la_iena_mprj[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(la_iena_mprj[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(la_iena_mprj[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(la_iena_mprj[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(la_iena_mprj[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(la_iena_mprj[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(la_iena_mprj[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(la_iena_mprj[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(la_iena_mprj[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(la_iena_mprj[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(la_iena_mprj[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(la_iena_mprj[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(la_iena_mprj[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(la_iena_mprj[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(la_iena_mprj[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(la_iena_mprj[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(la_iena_mprj[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(la_iena_mprj[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(la_iena_mprj[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(la_iena_mprj[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(la_iena_mprj[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(la_iena_mprj[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(la_iena_mprj[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(la_iena_mprj[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(la_iena_mprj[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(la_iena_mprj[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(la_iena_mprj[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(la_iena_mprj[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(la_iena_mprj[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(la_iena_mprj[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(la_iena_mprj[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(la_iena_mprj[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(la_iena_mprj[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input199_A (.DIODE(la_iena_mprj[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input200_A (.DIODE(la_iena_mprj[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input201_A (.DIODE(la_iena_mprj[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input202_A (.DIODE(la_iena_mprj[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input203_A (.DIODE(la_iena_mprj[49]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input204_A (.DIODE(la_iena_mprj[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input205_A (.DIODE(la_iena_mprj[50]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input206_A (.DIODE(la_iena_mprj[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input207_A (.DIODE(la_iena_mprj[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input208_A (.DIODE(la_iena_mprj[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input209_A (.DIODE(la_iena_mprj[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input210_A (.DIODE(la_iena_mprj[55]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input211_A (.DIODE(la_iena_mprj[56]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input212_A (.DIODE(la_iena_mprj[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input213_A (.DIODE(la_iena_mprj[58]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input214_A (.DIODE(la_iena_mprj[59]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input215_A (.DIODE(la_iena_mprj[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input216_A (.DIODE(la_iena_mprj[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input217_A (.DIODE(la_iena_mprj[61]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input218_A (.DIODE(la_iena_mprj[62]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input219_A (.DIODE(la_iena_mprj[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input220_A (.DIODE(la_iena_mprj[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input221_A (.DIODE(la_iena_mprj[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input222_A (.DIODE(la_iena_mprj[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input223_A (.DIODE(la_iena_mprj[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input224_A (.DIODE(la_iena_mprj[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input225_A (.DIODE(la_iena_mprj[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input226_A (.DIODE(la_iena_mprj[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input227_A (.DIODE(la_iena_mprj[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input228_A (.DIODE(la_iena_mprj[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input229_A (.DIODE(la_iena_mprj[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input230_A (.DIODE(la_iena_mprj[73]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input231_A (.DIODE(la_iena_mprj[74]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input232_A (.DIODE(la_iena_mprj[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input233_A (.DIODE(la_iena_mprj[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input234_A (.DIODE(la_iena_mprj[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input235_A (.DIODE(la_iena_mprj[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input236_A (.DIODE(la_iena_mprj[79]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input237_A (.DIODE(la_iena_mprj[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input238_A (.DIODE(la_iena_mprj[80]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input239_A (.DIODE(la_iena_mprj[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input240_A (.DIODE(la_iena_mprj[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input241_A (.DIODE(la_iena_mprj[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input242_A (.DIODE(la_iena_mprj[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input243_A (.DIODE(la_iena_mprj[85]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input244_A (.DIODE(la_iena_mprj[86]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input245_A (.DIODE(la_iena_mprj[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input246_A (.DIODE(la_iena_mprj[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input247_A (.DIODE(la_iena_mprj[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input248_A (.DIODE(la_iena_mprj[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input249_A (.DIODE(la_iena_mprj[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input250_A (.DIODE(la_iena_mprj[91]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input251_A (.DIODE(la_iena_mprj[92]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input252_A (.DIODE(la_iena_mprj[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input253_A (.DIODE(la_iena_mprj[94]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input254_A (.DIODE(la_iena_mprj[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input255_A (.DIODE(la_iena_mprj[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input256_A (.DIODE(la_iena_mprj[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input257_A (.DIODE(la_iena_mprj[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input258_A (.DIODE(la_iena_mprj[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input259_A (.DIODE(la_iena_mprj[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input260_A (.DIODE(la_oenb_mprj[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input261_A (.DIODE(la_oenb_mprj[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input262_A (.DIODE(la_oenb_mprj[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input263_A (.DIODE(la_oenb_mprj[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input264_A (.DIODE(la_oenb_mprj[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input265_A (.DIODE(la_oenb_mprj[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input266_A (.DIODE(la_oenb_mprj[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input267_A (.DIODE(la_oenb_mprj[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input268_A (.DIODE(la_oenb_mprj[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input269_A (.DIODE(la_oenb_mprj[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input270_A (.DIODE(la_oenb_mprj[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input271_A (.DIODE(la_oenb_mprj[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input272_A (.DIODE(la_oenb_mprj[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input273_A (.DIODE(la_oenb_mprj[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input274_A (.DIODE(la_oenb_mprj[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input275_A (.DIODE(la_oenb_mprj[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input276_A (.DIODE(la_oenb_mprj[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input277_A (.DIODE(la_oenb_mprj[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input278_A (.DIODE(la_oenb_mprj[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input279_A (.DIODE(la_oenb_mprj[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input280_A (.DIODE(la_oenb_mprj[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input281_A (.DIODE(la_oenb_mprj[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input282_A (.DIODE(la_oenb_mprj[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input283_A (.DIODE(la_oenb_mprj[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input284_A (.DIODE(la_oenb_mprj[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input285_A (.DIODE(la_oenb_mprj[122]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input286_A (.DIODE(la_oenb_mprj[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input287_A (.DIODE(la_oenb_mprj[124]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input288_A (.DIODE(la_oenb_mprj[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input289_A (.DIODE(la_oenb_mprj[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input290_A (.DIODE(la_oenb_mprj[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input291_A (.DIODE(la_oenb_mprj[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input292_A (.DIODE(la_oenb_mprj[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input293_A (.DIODE(la_oenb_mprj[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input294_A (.DIODE(la_oenb_mprj[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input295_A (.DIODE(la_oenb_mprj[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input296_A (.DIODE(la_oenb_mprj[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input297_A (.DIODE(la_oenb_mprj[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input298_A (.DIODE(la_oenb_mprj[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input299_A (.DIODE(la_oenb_mprj[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input300_A (.DIODE(la_oenb_mprj[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input301_A (.DIODE(la_oenb_mprj[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input302_A (.DIODE(la_oenb_mprj[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input303_A (.DIODE(la_oenb_mprj[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input304_A (.DIODE(la_oenb_mprj[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input305_A (.DIODE(la_oenb_mprj[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input306_A (.DIODE(la_oenb_mprj[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input307_A (.DIODE(la_oenb_mprj[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input308_A (.DIODE(la_oenb_mprj[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input309_A (.DIODE(la_oenb_mprj[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input310_A (.DIODE(la_oenb_mprj[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input311_A (.DIODE(la_oenb_mprj[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input312_A (.DIODE(la_oenb_mprj[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input313_A (.DIODE(la_oenb_mprj[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input314_A (.DIODE(la_oenb_mprj[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input315_A (.DIODE(la_oenb_mprj[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input316_A (.DIODE(la_oenb_mprj[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input317_A (.DIODE(la_oenb_mprj[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input318_A (.DIODE(la_oenb_mprj[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input319_A (.DIODE(la_oenb_mprj[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input320_A (.DIODE(la_oenb_mprj[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input321_A (.DIODE(la_oenb_mprj[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input322_A (.DIODE(la_oenb_mprj[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input323_A (.DIODE(la_oenb_mprj[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input324_A (.DIODE(la_oenb_mprj[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input325_A (.DIODE(la_oenb_mprj[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input326_A (.DIODE(la_oenb_mprj[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input327_A (.DIODE(la_oenb_mprj[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input328_A (.DIODE(la_oenb_mprj[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input329_A (.DIODE(la_oenb_mprj[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input330_A (.DIODE(la_oenb_mprj[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input331_A (.DIODE(la_oenb_mprj[49]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input332_A (.DIODE(la_oenb_mprj[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input333_A (.DIODE(la_oenb_mprj[50]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input334_A (.DIODE(la_oenb_mprj[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input335_A (.DIODE(la_oenb_mprj[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input336_A (.DIODE(la_oenb_mprj[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input337_A (.DIODE(la_oenb_mprj[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input338_A (.DIODE(la_oenb_mprj[55]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input339_A (.DIODE(la_oenb_mprj[56]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input340_A (.DIODE(la_oenb_mprj[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input341_A (.DIODE(la_oenb_mprj[58]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input342_A (.DIODE(la_oenb_mprj[59]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input343_A (.DIODE(la_oenb_mprj[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input344_A (.DIODE(la_oenb_mprj[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input345_A (.DIODE(la_oenb_mprj[61]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input346_A (.DIODE(la_oenb_mprj[62]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input347_A (.DIODE(la_oenb_mprj[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input348_A (.DIODE(la_oenb_mprj[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input349_A (.DIODE(la_oenb_mprj[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input350_A (.DIODE(la_oenb_mprj[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input351_A (.DIODE(la_oenb_mprj[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input352_A (.DIODE(la_oenb_mprj[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input353_A (.DIODE(la_oenb_mprj[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input354_A (.DIODE(la_oenb_mprj[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input355_A (.DIODE(la_oenb_mprj[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input356_A (.DIODE(la_oenb_mprj[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input357_A (.DIODE(la_oenb_mprj[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input358_A (.DIODE(la_oenb_mprj[73]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input359_A (.DIODE(la_oenb_mprj[74]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input360_A (.DIODE(la_oenb_mprj[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input361_A (.DIODE(la_oenb_mprj[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input362_A (.DIODE(la_oenb_mprj[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input363_A (.DIODE(la_oenb_mprj[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input364_A (.DIODE(la_oenb_mprj[79]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input365_A (.DIODE(la_oenb_mprj[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input366_A (.DIODE(la_oenb_mprj[80]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input367_A (.DIODE(la_oenb_mprj[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input368_A (.DIODE(la_oenb_mprj[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input369_A (.DIODE(la_oenb_mprj[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input370_A (.DIODE(la_oenb_mprj[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input371_A (.DIODE(la_oenb_mprj[85]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input372_A (.DIODE(la_oenb_mprj[86]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input373_A (.DIODE(la_oenb_mprj[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input374_A (.DIODE(la_oenb_mprj[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input375_A (.DIODE(la_oenb_mprj[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input376_A (.DIODE(la_oenb_mprj[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input377_A (.DIODE(la_oenb_mprj[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input378_A (.DIODE(la_oenb_mprj[91]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input379_A (.DIODE(la_oenb_mprj[92]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input380_A (.DIODE(la_oenb_mprj[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input381_A (.DIODE(la_oenb_mprj[94]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input382_A (.DIODE(la_oenb_mprj[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input383_A (.DIODE(la_oenb_mprj[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input384_A (.DIODE(la_oenb_mprj[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input385_A (.DIODE(la_oenb_mprj[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input386_A (.DIODE(la_oenb_mprj[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input387_A (.DIODE(la_oenb_mprj[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_user_wb_ack_gate_A (.DIODE(mprj_ack_i_user));
 sky130_fd_sc_hd__diode_2 ANTENNA_input388_A (.DIODE(mprj_adr_o_core[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input389_A (.DIODE(mprj_adr_o_core[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input390_A (.DIODE(mprj_adr_o_core[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input391_A (.DIODE(mprj_adr_o_core[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input392_A (.DIODE(mprj_adr_o_core[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input393_A (.DIODE(mprj_adr_o_core[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input394_A (.DIODE(mprj_adr_o_core[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input395_A (.DIODE(mprj_adr_o_core[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input396_A (.DIODE(mprj_adr_o_core[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input397_A (.DIODE(mprj_adr_o_core[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input398_A (.DIODE(mprj_adr_o_core[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input399_A (.DIODE(mprj_adr_o_core[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input400_A (.DIODE(mprj_adr_o_core[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input401_A (.DIODE(mprj_adr_o_core[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input402_A (.DIODE(mprj_adr_o_core[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input403_A (.DIODE(mprj_adr_o_core[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input404_A (.DIODE(mprj_adr_o_core[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input405_A (.DIODE(mprj_adr_o_core[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input406_A (.DIODE(mprj_adr_o_core[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input407_A (.DIODE(mprj_adr_o_core[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input408_A (.DIODE(mprj_adr_o_core[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input409_A (.DIODE(mprj_adr_o_core[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input410_A (.DIODE(mprj_adr_o_core[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input411_A (.DIODE(mprj_adr_o_core[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input412_A (.DIODE(mprj_adr_o_core[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input413_A (.DIODE(mprj_adr_o_core[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input414_A (.DIODE(mprj_adr_o_core[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input415_A (.DIODE(mprj_adr_o_core[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input416_A (.DIODE(mprj_adr_o_core[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input417_A (.DIODE(mprj_adr_o_core[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input418_A (.DIODE(mprj_adr_o_core[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input419_A (.DIODE(mprj_adr_o_core[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input420_A (.DIODE(mprj_cyc_o_core));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__A (.DIODE(\mprj_dat_i_core_bar[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0592__A (.DIODE(\mprj_dat_i_core_bar[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__A (.DIODE(\mprj_dat_i_core_bar[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__A (.DIODE(\mprj_dat_i_core_bar[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__A (.DIODE(\mprj_dat_i_core_bar[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__A (.DIODE(\mprj_dat_i_core_bar[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__A (.DIODE(\mprj_dat_i_core_bar[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[0]_A  (.DIODE(mprj_dat_i_user[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[10]_A  (.DIODE(mprj_dat_i_user[10]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[11]_A  (.DIODE(mprj_dat_i_user[11]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[12]_A  (.DIODE(mprj_dat_i_user[12]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[13]_A  (.DIODE(mprj_dat_i_user[13]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[14]_A  (.DIODE(mprj_dat_i_user[14]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[15]_A  (.DIODE(mprj_dat_i_user[15]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[16]_A  (.DIODE(mprj_dat_i_user[16]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[17]_A  (.DIODE(mprj_dat_i_user[17]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[18]_A  (.DIODE(mprj_dat_i_user[18]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[19]_A  (.DIODE(mprj_dat_i_user[19]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[1]_A  (.DIODE(mprj_dat_i_user[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[20]_A  (.DIODE(mprj_dat_i_user[20]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[21]_A  (.DIODE(mprj_dat_i_user[21]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[22]_A  (.DIODE(mprj_dat_i_user[22]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[23]_A  (.DIODE(mprj_dat_i_user[23]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[24]_A  (.DIODE(mprj_dat_i_user[24]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[25]_A  (.DIODE(mprj_dat_i_user[25]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[26]_A  (.DIODE(mprj_dat_i_user[26]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[27]_A  (.DIODE(mprj_dat_i_user[27]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[28]_A  (.DIODE(mprj_dat_i_user[28]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[29]_A  (.DIODE(mprj_dat_i_user[29]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[2]_A  (.DIODE(mprj_dat_i_user[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[30]_A  (.DIODE(mprj_dat_i_user[30]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[31]_A  (.DIODE(mprj_dat_i_user[31]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[3]_A  (.DIODE(mprj_dat_i_user[3]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[4]_A  (.DIODE(mprj_dat_i_user[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[5]_A  (.DIODE(mprj_dat_i_user[5]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[6]_A  (.DIODE(mprj_dat_i_user[6]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[7]_A  (.DIODE(mprj_dat_i_user[7]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[8]_A  (.DIODE(mprj_dat_i_user[8]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[9]_A  (.DIODE(mprj_dat_i_user[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input421_A (.DIODE(mprj_dat_o_core[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input422_A (.DIODE(mprj_dat_o_core[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input423_A (.DIODE(mprj_dat_o_core[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input424_A (.DIODE(mprj_dat_o_core[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input425_A (.DIODE(mprj_dat_o_core[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input426_A (.DIODE(mprj_dat_o_core[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input427_A (.DIODE(mprj_dat_o_core[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input428_A (.DIODE(mprj_dat_o_core[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input429_A (.DIODE(mprj_dat_o_core[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input430_A (.DIODE(mprj_dat_o_core[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input431_A (.DIODE(mprj_dat_o_core[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input432_A (.DIODE(mprj_dat_o_core[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input433_A (.DIODE(mprj_dat_o_core[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input434_A (.DIODE(mprj_dat_o_core[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input435_A (.DIODE(mprj_dat_o_core[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input436_A (.DIODE(mprj_dat_o_core[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input437_A (.DIODE(mprj_dat_o_core[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input438_A (.DIODE(mprj_dat_o_core[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input439_A (.DIODE(mprj_dat_o_core[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input440_A (.DIODE(mprj_dat_o_core[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input441_A (.DIODE(mprj_dat_o_core[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input442_A (.DIODE(mprj_dat_o_core[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input443_A (.DIODE(mprj_dat_o_core[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input444_A (.DIODE(mprj_dat_o_core[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input445_A (.DIODE(mprj_dat_o_core[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input446_A (.DIODE(mprj_dat_o_core[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input447_A (.DIODE(mprj_dat_o_core[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input448_A (.DIODE(mprj_dat_o_core[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input449_A (.DIODE(mprj_dat_o_core[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input450_A (.DIODE(mprj_dat_o_core[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input451_A (.DIODE(mprj_dat_o_core[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input452_A (.DIODE(mprj_dat_o_core[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input453_A (.DIODE(mprj_iena_wb));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2847_A (.DIODE(\mprj_logic1[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2844_A (.DIODE(\mprj_logic1[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2838_A (.DIODE(\mprj_logic1[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__B (.DIODE(\mprj_logic1[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__B (.DIODE(\mprj_logic1[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2837_A (.DIODE(\mprj_logic1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__B (.DIODE(\mprj_logic1[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__B (.DIODE(\mprj_logic1[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__B (.DIODE(\mprj_logic1[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2836_A (.DIODE(\mprj_logic1[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2835_A (.DIODE(\mprj_logic1[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__B (.DIODE(\mprj_logic1[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2834_A (.DIODE(\mprj_logic1[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__B (.DIODE(\mprj_logic1[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__B (.DIODE(\mprj_logic1[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__A (.DIODE(\mprj_logic1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__B (.DIODE(\mprj_logic1[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__B (.DIODE(\mprj_logic1[122] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__B (.DIODE(\mprj_logic1[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__B (.DIODE(\mprj_logic1[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2832_A (.DIODE(\mprj_logic1[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2830_A (.DIODE(\mprj_logic1[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__B (.DIODE(\mprj_logic1[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2829_A (.DIODE(\mprj_logic1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__B (.DIODE(\mprj_logic1[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__B (.DIODE(\mprj_logic1[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__B (.DIODE(\mprj_logic1[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__B (.DIODE(\mprj_logic1[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__B (.DIODE(\mprj_logic1[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__B (.DIODE(\mprj_logic1[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__B (.DIODE(\mprj_logic1[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__B (.DIODE(\mprj_logic1[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__B (.DIODE(\mprj_logic1[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A (.DIODE(\mprj_logic1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__B (.DIODE(\mprj_logic1[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2827_A (.DIODE(\mprj_logic1[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2826_A (.DIODE(\mprj_logic1[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2824_A (.DIODE(\mprj_logic1[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2823_A (.DIODE(\mprj_logic1[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2821_A (.DIODE(\mprj_logic1[145] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2819_A (.DIODE(\mprj_logic1[146] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2815_A (.DIODE(\mprj_logic1[148] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2812_A (.DIODE(\mprj_logic1[149] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2809_A (.DIODE(\mprj_logic1[150] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2806_A (.DIODE(\mprj_logic1[151] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2803_A (.DIODE(\mprj_logic1[152] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2790_A (.DIODE(\mprj_logic1[156] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2782_A (.DIODE(\mprj_logic1[158] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2779_A (.DIODE(\mprj_logic1[159] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__A (.DIODE(\mprj_logic1[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2775_A (.DIODE(\mprj_logic1[160] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2763_A (.DIODE(\mprj_logic1[163] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2761_A (.DIODE(\mprj_logic1[165] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2760_A (.DIODE(\mprj_logic1[166] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__B (.DIODE(\mprj_logic1[167] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2759_A (.DIODE(\mprj_logic1[168] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2755_A (.DIODE(\mprj_logic1[171] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2754_A (.DIODE(\mprj_logic1[172] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2753_A (.DIODE(\mprj_logic1[173] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2750_A (.DIODE(\mprj_logic1[175] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2747_A (.DIODE(\mprj_logic1[177] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2745_A (.DIODE(\mprj_logic1[178] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2742_A (.DIODE(\mprj_logic1[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2735_A (.DIODE(\mprj_logic1[183] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2733_A (.DIODE(\mprj_logic1[184] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2731_A (.DIODE(\mprj_logic1[185] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2728_A (.DIODE(\mprj_logic1[186] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2726_A (.DIODE(\mprj_logic1[187] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__A (.DIODE(\mprj_logic1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2718_A (.DIODE(\mprj_logic1[190] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2715_A (.DIODE(\mprj_logic1[191] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2713_A (.DIODE(\mprj_logic1[192] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2710_A (.DIODE(\mprj_logic1[193] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2704_A (.DIODE(\mprj_logic1[195] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2700_A (.DIODE(\mprj_logic1[196] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2697_A (.DIODE(\mprj_logic1[197] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__A (.DIODE(\mprj_logic1[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A (.DIODE(\mprj_logic1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2686_A (.DIODE(\mprj_logic1[200] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2682_A (.DIODE(\mprj_logic1[201] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2679_A (.DIODE(\mprj_logic1[202] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2677_A (.DIODE(\mprj_logic1[203] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2674_A (.DIODE(\mprj_logic1[204] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2671_A (.DIODE(\mprj_logic1[205] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2668_A (.DIODE(\mprj_logic1[206] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2666_A (.DIODE(\mprj_logic1[207] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2663_A (.DIODE(\mprj_logic1[208] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2660_A (.DIODE(\mprj_logic1[209] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__A (.DIODE(\mprj_logic1[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2658_A (.DIODE(\mprj_logic1[210] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2656_A (.DIODE(\mprj_logic1[211] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2650_A (.DIODE(\mprj_logic1[213] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2648_A (.DIODE(\mprj_logic1[214] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2641_A (.DIODE(\mprj_logic1[217] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2639_A (.DIODE(\mprj_logic1[218] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2637_A (.DIODE(\mprj_logic1[219] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2629_A (.DIODE(\mprj_logic1[222] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2627_A (.DIODE(\mprj_logic1[223] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2626_A (.DIODE(\mprj_logic1[224] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2622_A (.DIODE(\mprj_logic1[226] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2621_A (.DIODE(\mprj_logic1[227] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2619_A (.DIODE(\mprj_logic1[229] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2617_A (.DIODE(\mprj_logic1[230] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2615_A (.DIODE(\mprj_logic1[232] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2612_A (.DIODE(\mprj_logic1[234] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2611_A (.DIODE(\mprj_logic1[235] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__B (.DIODE(\mprj_logic1[237] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2609_A (.DIODE(\mprj_logic1[238] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__B (.DIODE(\mprj_logic1[239] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__B (.DIODE(\mprj_logic1[240] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__B (.DIODE(\mprj_logic1[241] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__B (.DIODE(\mprj_logic1[242] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2608_A (.DIODE(\mprj_logic1[243] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__B (.DIODE(\mprj_logic1[244] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__B (.DIODE(\mprj_logic1[245] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1363__B (.DIODE(\mprj_logic1[246] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__B (.DIODE(\mprj_logic1[247] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2607_A (.DIODE(\mprj_logic1[248] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__B (.DIODE(\mprj_logic1[249] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__A (.DIODE(\mprj_logic1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2606_A (.DIODE(\mprj_logic1[250] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2605_A (.DIODE(\mprj_logic1[252] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2604_A (.DIODE(\mprj_logic1[254] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__B (.DIODE(\mprj_logic1[256] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2602_A (.DIODE(\mprj_logic1[257] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__B (.DIODE(\mprj_logic1[258] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__A (.DIODE(\mprj_logic1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__B (.DIODE(\mprj_logic1[260] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2600_A (.DIODE(\mprj_logic1[261] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__B (.DIODE(\mprj_logic1[262] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__B (.DIODE(\mprj_logic1[263] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__B (.DIODE(\mprj_logic1[264] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B (.DIODE(\mprj_logic1[265] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2599_A (.DIODE(\mprj_logic1[266] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__B (.DIODE(\mprj_logic1[267] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2598_A (.DIODE(\mprj_logic1[268] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__B (.DIODE(\mprj_logic1[269] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2594_A (.DIODE(\mprj_logic1[271] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2593_A (.DIODE(\mprj_logic1[272] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2588_A (.DIODE(\mprj_logic1[275] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2587_A (.DIODE(\mprj_logic1[276] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2585_A (.DIODE(\mprj_logic1[277] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2574_A (.DIODE(\mprj_logic1[281] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2572_A (.DIODE(\mprj_logic1[282] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2569_A (.DIODE(\mprj_logic1[283] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2563_A (.DIODE(\mprj_logic1[285] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2560_A (.DIODE(\mprj_logic1[286] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2550_A (.DIODE(\mprj_logic1[289] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2546_A (.DIODE(\mprj_logic1[290] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2543_A (.DIODE(\mprj_logic1[291] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2541_A (.DIODE(\mprj_logic1[293] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__B (.DIODE(\mprj_logic1[294] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2538_A (.DIODE(\mprj_logic1[296] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2536_A (.DIODE(\mprj_logic1[297] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2530_A (.DIODE(\mprj_logic1[299] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__A (.DIODE(\mprj_logic1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2517_A (.DIODE(\mprj_logic1[302] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2514_A (.DIODE(\mprj_logic1[303] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2511_A (.DIODE(\mprj_logic1[304] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2505_A (.DIODE(\mprj_logic1[306] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2500_A (.DIODE(\mprj_logic1[308] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2497_A (.DIODE(\mprj_logic1[309] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__A (.DIODE(\mprj_logic1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2494_A (.DIODE(\mprj_logic1[310] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2491_A (.DIODE(\mprj_logic1[311] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2488_A (.DIODE(\mprj_logic1[312] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2481_A (.DIODE(\mprj_logic1[314] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2476_A (.DIODE(\mprj_logic1[316] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2468_A (.DIODE(\mprj_logic1[318] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2465_A (.DIODE(\mprj_logic1[319] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2461_A (.DIODE(\mprj_logic1[320] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2458_A (.DIODE(\mprj_logic1[321] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2454_A (.DIODE(\mprj_logic1[322] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2446_A (.DIODE(\mprj_logic1[324] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2442_A (.DIODE(\mprj_logic1[325] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2434_A (.DIODE(\mprj_logic1[327] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2430_A (.DIODE(\mprj_logic1[328] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__A (.DIODE(\mprj_logic1[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2421_A (.DIODE(\mprj_logic1[330] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2419_A (.DIODE(\mprj_logic1[331] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2416_A (.DIODE(\mprj_logic1[332] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2414_A (.DIODE(\mprj_logic1[333] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2407_A (.DIODE(\mprj_logic1[336] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2406_A (.DIODE(\mprj_logic1[337] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2404_A (.DIODE(\mprj_logic1[338] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2403_A (.DIODE(\mprj_logic1[339] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2391_A (.DIODE(\mprj_logic1[344] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2389_A (.DIODE(\mprj_logic1[345] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2385_A (.DIODE(\mprj_logic1[347] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2383_A (.DIODE(\mprj_logic1[348] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2381_A (.DIODE(\mprj_logic1[349] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__A (.DIODE(\mprj_logic1[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2379_A (.DIODE(\mprj_logic1[350] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2377_A (.DIODE(\mprj_logic1[351] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2376_A (.DIODE(\mprj_logic1[352] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2371_A (.DIODE(\mprj_logic1[354] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2367_A (.DIODE(\mprj_logic1[356] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2365_A (.DIODE(\mprj_logic1[357] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2364_A (.DIODE(\mprj_logic1[358] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__A (.DIODE(\mprj_logic1[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2358_A (.DIODE(\mprj_logic1[361] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2357_A (.DIODE(\mprj_logic1[362] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2354_A (.DIODE(\mprj_logic1[364] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2351_A (.DIODE(\mprj_logic1[366] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__A (.DIODE(\mprj_logic1[367] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2348_A (.DIODE(\mprj_logic1[369] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2347_A (.DIODE(\mprj_logic1[370] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2346_A (.DIODE(\mprj_logic1[371] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2345_A (.DIODE(\mprj_logic1[372] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2344_A (.DIODE(\mprj_logic1[373] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2343_A (.DIODE(\mprj_logic1[374] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2342_A (.DIODE(\mprj_logic1[375] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2341_A (.DIODE(\mprj_logic1[376] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2340_A (.DIODE(\mprj_logic1[377] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2339_A (.DIODE(\mprj_logic1[378] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A (.DIODE(\mprj_logic1[379] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A (.DIODE(\mprj_logic1[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2338_A (.DIODE(\mprj_logic1[380] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2337_A (.DIODE(\mprj_logic1[381] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2336_A (.DIODE(\mprj_logic1[382] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2335_A (.DIODE(\mprj_logic1[383] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2334_A (.DIODE(\mprj_logic1[384] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__A (.DIODE(\mprj_logic1[385] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2332_A (.DIODE(\mprj_logic1[387] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A (.DIODE(\mprj_logic1[388] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__A (.DIODE(\mprj_logic1[389] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__A (.DIODE(\mprj_logic1[392] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__A (.DIODE(\mprj_logic1[394] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__A (.DIODE(\mprj_logic1[399] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2329_A (.DIODE(\mprj_logic1[400] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2328_A (.DIODE(\mprj_logic1[401] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2327_A (.DIODE(\mprj_logic1[402] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2322_A (.DIODE(\mprj_logic1[405] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2320_A (.DIODE(\mprj_logic1[406] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2319_A (.DIODE(\mprj_logic1[407] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2318_A (.DIODE(\mprj_logic1[408] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2317_A (.DIODE(\mprj_logic1[409] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__A (.DIODE(\mprj_logic1[411] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A (.DIODE(\mprj_logic1[412] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2312_A (.DIODE(\mprj_logic1[414] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2311_A (.DIODE(\mprj_logic1[415] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2309_A (.DIODE(\mprj_logic1[417] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2305_A (.DIODE(\mprj_logic1[419] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__A (.DIODE(\mprj_logic1[420] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2301_A (.DIODE(\mprj_logic1[424] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2299_A (.DIODE(\mprj_logic1[426] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2297_A (.DIODE(\mprj_logic1[428] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2296_A (.DIODE(\mprj_logic1[429] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2295_A (.DIODE(\mprj_logic1[430] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A (.DIODE(\mprj_logic1[431] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__A (.DIODE(\mprj_logic1[433] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2292_A (.DIODE(\mprj_logic1[435] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2291_A (.DIODE(\mprj_logic1[436] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2289_A (.DIODE(\mprj_logic1[437] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2283_A (.DIODE(\mprj_logic1[439] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2280_A (.DIODE(\mprj_logic1[440] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2278_A (.DIODE(\mprj_logic1[441] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2275_A (.DIODE(\mprj_logic1[442] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2272_A (.DIODE(\mprj_logic1[443] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2269_A (.DIODE(\mprj_logic1[444] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2267_A (.DIODE(\mprj_logic1[445] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2263_A (.DIODE(\mprj_logic1[446] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2258_A (.DIODE(\mprj_logic1[448] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2255_A (.DIODE(\mprj_logic1[449] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2253_A (.DIODE(\mprj_logic1[44] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2252_A (.DIODE(\mprj_logic1[450] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2248_A (.DIODE(\mprj_logic1[451] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2245_A (.DIODE(\mprj_logic1[452] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2242_A (.DIODE(\mprj_logic1[453] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2239_A (.DIODE(\mprj_logic1[454] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2236_A (.DIODE(\mprj_logic1[455] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2233_A (.DIODE(\mprj_logic1[456] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2230_A (.DIODE(\mprj_logic1[457] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2220_A (.DIODE(\mprj_logic1[460] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__A (.DIODE(\mprj_logic1[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__A (.DIODE(\mprj_logic1[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2208_A (.DIODE(\mprj_logic1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A (.DIODE(\mprj_logic1[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2207_A (.DIODE(\mprj_logic1[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2206_A (.DIODE(\mprj_logic1[52] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2203_A (.DIODE(\mprj_logic1[54] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2201_A (.DIODE(\mprj_logic1[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__A (.DIODE(\mprj_logic1[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2198_A (.DIODE(\mprj_logic1[58] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2195_A (.DIODE(\mprj_logic1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2194_A (.DIODE(\mprj_logic1[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2193_A (.DIODE(\mprj_logic1[61] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2190_A (.DIODE(\mprj_logic1[63] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2189_A (.DIODE(\mprj_logic1[64] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2188_A (.DIODE(\mprj_logic1[65] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2181_A (.DIODE(\mprj_logic1[68] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2175_A (.DIODE(\mprj_logic1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2173_A (.DIODE(\mprj_logic1[70] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2169_A (.DIODE(\mprj_logic1[72] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2168_A (.DIODE(\mprj_logic1[73] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2167_A (.DIODE(\mprj_logic1[74] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2164_A (.DIODE(\mprj_logic1[75] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2161_A (.DIODE(\mprj_logic1[76] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2158_A (.DIODE(\mprj_logic1[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2155_A (.DIODE(\mprj_logic1[78] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2152_A (.DIODE(\mprj_logic1[79] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2149_A (.DIODE(\mprj_logic1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2143_A (.DIODE(\mprj_logic1[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2139_A (.DIODE(\mprj_logic1[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2121_A (.DIODE(\mprj_logic1[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2110_A (.DIODE(\mprj_logic1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2098_A (.DIODE(\mprj_logic1[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2091_A (.DIODE(\mprj_logic1[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2088_A (.DIODE(\mprj_logic1[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2085_A (.DIODE(\mprj_logic1[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2080_A (.DIODE(\mprj_logic1[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input454_A (.DIODE(mprj_sel_o_core[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input455_A (.DIODE(mprj_sel_o_core[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input456_A (.DIODE(mprj_sel_o_core[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input457_A (.DIODE(mprj_sel_o_core[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input458_A (.DIODE(mprj_stb_o_core));
 sky130_fd_sc_hd__diode_2 ANTENNA_input459_A (.DIODE(mprj_we_o_core));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_irq_gates[0]_A  (.DIODE(user_irq_core[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_irq_gates[1]_A  (.DIODE(user_irq_core[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_irq_gates[2]_A  (.DIODE(user_irq_core[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input460_A (.DIODE(user_irq_ena[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input461_A (.DIODE(user_irq_ena[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input462_A (.DIODE(user_irq_ena[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1327_A (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[31]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[30]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[29]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[26]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[25]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[24]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[23]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[22]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[21]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[14]_B  (.DIODE(wb_in_enable));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1936_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__C (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__C (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__C (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__C (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__C (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__C (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__C (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__C (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__C (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__C (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__C (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1919_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__C (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__C (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__C (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__C (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__C (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__C (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__C (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__C (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__C (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__C (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__C (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__C (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__C (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__C (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__C (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__C (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__C (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__C (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__C (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__C (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1644_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1642_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1639_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1635_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1634_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__C (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1633_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2063_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2062_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2061_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2059_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2058_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2053_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2047_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2039_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2037_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2032_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2029_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__C (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__0813__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2025_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2024_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2022_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2019_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2018_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2012_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2011_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2010_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__B (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__B (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__B (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__0717__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1993_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__0725__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__0731__B (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__B (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__0735__B (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__0741__B (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__0743__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1989_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1988_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1987_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1982_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1979_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__B (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__B (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1978_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__B (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1976_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__B (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__B (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__A_N (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1971_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__A_N (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1968_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__A_N (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1967_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__A_N (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1964_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__A_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1962_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__A_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1959_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1295__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1947_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__A_N (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1943_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__A_N (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1942_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__A_N (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1940_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__A_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A_N (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__A_N (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A_N (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A_N (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A_N (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__A_N (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__A_N (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__A_N (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__A_N (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__A_N (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__A_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1925_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1924_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA__1279__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__A_N (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A_N (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__A_N (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A_N (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1921_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A_N (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__A_N (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__A_N (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__A_N (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1915_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1913_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__A_N (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1912_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__A_N (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1910_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1909_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1906_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A_N (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A_N (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__A (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__A_N (.DIODE(net332));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1903_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A_N (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1900_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1898_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1897_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__A_N (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__A_N (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1883_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1882_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1881_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A_N (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1875_A (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A_N (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1873_A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1872_A (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1871_A (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1870_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1869_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1867_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1866_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1864_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A_N (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1858_A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1856_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1854_A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1852_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1850_A (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1848_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1846_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1844_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1842_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A_N (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__A_N (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__A (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__A_N (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__A_N (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1840_A (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__A_N (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1839_A (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__A_N (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1838_A (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__A_N (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1835_A (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__A_N (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1834_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__A_N (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A_N (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1830_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1817_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1806_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1801_A (.DIODE(net396));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1798_A (.DIODE(net397));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1793_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1789_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1785_A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1782_A (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1760_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1751_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1747_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1742_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1737_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1733_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1729_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1720_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1716_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1693_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__B (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1688_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1683_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1682_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1673_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__B (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__B (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__B (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__B (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1670_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1669_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1668_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1661_A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1659_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1657_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1653_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1651_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__B (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__B (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__B (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__B (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__B (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1148_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_output464_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1099_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_output470_A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_output472_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_output478_A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_output482_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_output483_A (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 ANTENNA_output484_A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_output486_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_output487_A (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_output488_A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_output489_A (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_output491_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_output492_A (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1138_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_output496_A (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_output505_A (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 ANTENNA_output506_A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_output508_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1131_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1128_A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1145_A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_output514_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1126_A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1121_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_output519_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_output520_A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_output521_A (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA_output522_A (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_output523_A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1144_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1120_A (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA_output529_A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_output530_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_output531_A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_output534_A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1143_A (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA_output536_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_output538_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_output544_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1142_A (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA_output550_A (.DIODE(net550));
 sky130_fd_sc_hd__diode_2 ANTENNA_output552_A (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA_output554_A (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA_output555_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_output556_A (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1141_A (.DIODE(net557));
 sky130_fd_sc_hd__diode_2 ANTENNA_output559_A (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA_output562_A (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA_output563_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_output564_A (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA_output565_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_output566_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_output567_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1118_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1117_A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1116_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1115_A (.DIODE(net572));
 sky130_fd_sc_hd__diode_2 ANTENNA_output574_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1113_A (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1112_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1111_A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_output579_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_output580_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1108_A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1107_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1106_A (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1105_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_output587_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1102_A (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire993_A (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA_output597_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire990_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire989_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire986_A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire985_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire981_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire971_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_output612_A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire970_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire969_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire968_A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire967_A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_output618_A (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA_output620_A (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_output621_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_output623_A (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA_output624_A (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA_output626_A (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA_output628_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1011_A (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_output633_A (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA_output635_A (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1009_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_output638_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1007_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_output644_A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1003_A (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1002_A (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_output648_A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_output651_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_output654_A (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire998_A (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA_output656_A (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_output657_A (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire997_A (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_output659_A (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA_output661_A (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_output664_A (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA_output667_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_output668_A (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA_output670_A (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_output671_A (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA_output689_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_output696_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_output703_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_output706_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_output707_A (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_output709_A (.DIODE(net709));
 sky130_fd_sc_hd__diode_2 ANTENNA_output718_A (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA_output721_A (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_output722_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output723_A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output724_A (.DIODE(net724));
 sky130_fd_sc_hd__diode_2 ANTENNA_output726_A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA_output727_A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA_output728_A (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA_output731_A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA_output732_A (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA_output733_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_output734_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_output735_A (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_output737_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_output739_A (.DIODE(net739));
 sky130_fd_sc_hd__diode_2 ANTENNA_output741_A (.DIODE(net741));
 sky130_fd_sc_hd__diode_2 ANTENNA_output743_A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_output744_A (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA_output756_A (.DIODE(net756));
 sky130_fd_sc_hd__diode_2 ANTENNA_output757_A (.DIODE(net757));
 sky130_fd_sc_hd__diode_2 ANTENNA_output758_A (.DIODE(net758));
 sky130_fd_sc_hd__diode_2 ANTENNA_output759_A (.DIODE(net759));
 sky130_fd_sc_hd__diode_2 ANTENNA_output769_A (.DIODE(net769));
 sky130_fd_sc_hd__diode_2 ANTENNA_output776_A (.DIODE(net776));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1092_A (.DIODE(net779));
 sky130_fd_sc_hd__diode_2 ANTENNA_output780_A (.DIODE(net780));
 sky130_fd_sc_hd__diode_2 ANTENNA_output782_A (.DIODE(net782));
 sky130_fd_sc_hd__diode_2 ANTENNA_output783_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_output785_A (.DIODE(net785));
 sky130_fd_sc_hd__diode_2 ANTENNA_output789_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_output790_A (.DIODE(net790));
 sky130_fd_sc_hd__diode_2 ANTENNA_output792_A (.DIODE(net792));
 sky130_fd_sc_hd__diode_2 ANTENNA_output793_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_output795_A (.DIODE(net795));
 sky130_fd_sc_hd__diode_2 ANTENNA_output798_A (.DIODE(net798));
 sky130_fd_sc_hd__diode_2 ANTENNA_output802_A (.DIODE(net802));
 sky130_fd_sc_hd__diode_2 ANTENNA_output803_A (.DIODE(net803));
 sky130_fd_sc_hd__diode_2 ANTENNA_output806_A (.DIODE(net806));
 sky130_fd_sc_hd__diode_2 ANTENNA_output807_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_output809_A (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output810_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_output818_A (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA_output820_A (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_output825_A (.DIODE(net825));
 sky130_fd_sc_hd__diode_2 ANTENNA_output827_A (.DIODE(net827));
 sky130_fd_sc_hd__diode_2 ANTENNA_output828_A (.DIODE(net828));
 sky130_fd_sc_hd__diode_2 ANTENNA_output829_A (.DIODE(net829));
 sky130_fd_sc_hd__diode_2 ANTENNA_output830_A (.DIODE(net830));
 sky130_fd_sc_hd__diode_2 ANTENNA_output831_A (.DIODE(net831));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1087_A (.DIODE(net833));
 sky130_fd_sc_hd__diode_2 ANTENNA_output839_A (.DIODE(net839));
 sky130_fd_sc_hd__diode_2 ANTENNA_output841_A (.DIODE(net841));
 sky130_fd_sc_hd__diode_2 ANTENNA_output844_A (.DIODE(net844));
 sky130_fd_sc_hd__diode_2 ANTENNA_output845_A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA_output847_A (.DIODE(net847));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1276_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1273_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1271_A (.DIODE(net852));
 sky130_fd_sc_hd__diode_2 ANTENNA_output855_A (.DIODE(net855));
 sky130_fd_sc_hd__diode_2 ANTENNA_output857_A (.DIODE(net857));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1262_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1290_A (.DIODE(net859));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1261_A (.DIODE(net860));
 sky130_fd_sc_hd__diode_2 ANTENNA_output861_A (.DIODE(net861));
 sky130_fd_sc_hd__diode_2 ANTENNA_output864_A (.DIODE(net864));
 sky130_fd_sc_hd__diode_2 ANTENNA_output865_A (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1254_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1253_A (.DIODE(net867));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1252_A (.DIODE(net868));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1251_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_output870_A (.DIODE(net870));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1289_A (.DIODE(net873));
 sky130_fd_sc_hd__diode_2 ANTENNA_output874_A (.DIODE(net874));
 sky130_fd_sc_hd__diode_2 ANTENNA_output877_A (.DIODE(net877));
 sky130_fd_sc_hd__diode_2 ANTENNA_output878_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1321_A (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA_output881_A (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_output882_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_output883_A (.DIODE(net883));
 sky130_fd_sc_hd__diode_2 ANTENNA_output884_A (.DIODE(net884));
 sky130_fd_sc_hd__diode_2 ANTENNA_output887_A (.DIODE(net887));
 sky130_fd_sc_hd__diode_2 ANTENNA_output889_A (.DIODE(net889));
 sky130_fd_sc_hd__diode_2 ANTENNA_output892_A (.DIODE(net892));
 sky130_fd_sc_hd__diode_2 ANTENNA_output901_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_output906_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_output908_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_output909_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire963_A (.DIODE(net910));
 sky130_fd_sc_hd__diode_2 ANTENNA_output911_A (.DIODE(net911));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1246_A (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1213_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1210_A (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1199_A (.DIODE(net918));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1196_A (.DIODE(net919));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1193_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1190_A (.DIODE(net921));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1187_A (.DIODE(net922));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1243_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1182_A (.DIODE(net925));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1173_A (.DIODE(net928));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1170_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1167_A (.DIODE(net930));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1164_A (.DIODE(net931));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1161_A (.DIODE(net932));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1158_A (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1240_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1152_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1150_A (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1237_A (.DIODE(net938));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1234_A (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1223_A (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1216_A (.DIODE(net944));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1295_A (.DIODE(net948));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1318_A (.DIODE(net949));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2217_A (.DIODE(net951));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2071_A (.DIODE(net952));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2855_A (.DIODE(net953));
 sky130_fd_sc_hd__diode_2 ANTENNA_output960_A (.DIODE(net960));
 sky130_fd_sc_hd__diode_2 ANTENNA_output625_A (.DIODE(net961));
 sky130_fd_sc_hd__diode_2 ANTENNA_output602_A (.DIODE(net962));
 sky130_fd_sc_hd__diode_2 ANTENNA_output910_A (.DIODE(net963));
 sky130_fd_sc_hd__diode_2 ANTENNA_output907_A (.DIODE(net964));
 sky130_fd_sc_hd__diode_2 ANTENNA_output903_A (.DIODE(net965));
 sky130_fd_sc_hd__diode_2 ANTENNA_output619_A (.DIODE(net966));
 sky130_fd_sc_hd__diode_2 ANTENNA_output617_A (.DIODE(net967));
 sky130_fd_sc_hd__diode_2 ANTENNA_output616_A (.DIODE(net968));
 sky130_fd_sc_hd__diode_2 ANTENNA_output615_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_output614_A (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_output611_A (.DIODE(net971));
 sky130_fd_sc_hd__diode_2 ANTENNA_output610_A (.DIODE(net972));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire972_A (.DIODE(net973));
 sky130_fd_sc_hd__diode_2 ANTENNA_output609_A (.DIODE(net974));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire974_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_output608_A (.DIODE(net976));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire976_A (.DIODE(net977));
 sky130_fd_sc_hd__diode_2 ANTENNA_output607_A (.DIODE(net978));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire978_A (.DIODE(net979));
 sky130_fd_sc_hd__diode_2 ANTENNA_output606_A (.DIODE(net980));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire980_A (.DIODE(net981));
 sky130_fd_sc_hd__diode_2 ANTENNA_output605_A (.DIODE(net982));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire982_A (.DIODE(net983));
 sky130_fd_sc_hd__diode_2 ANTENNA_output604_A (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire984_A (.DIODE(net985));
 sky130_fd_sc_hd__diode_2 ANTENNA_output603_A (.DIODE(net986));
 sky130_fd_sc_hd__diode_2 ANTENNA_output601_A (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire987_A (.DIODE(net988));
 sky130_fd_sc_hd__diode_2 ANTENNA_output600_A (.DIODE(net989));
 sky130_fd_sc_hd__diode_2 ANTENNA_output599_A (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_output598_A (.DIODE(net991));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire991_A (.DIODE(net992));
 sky130_fd_sc_hd__diode_2 ANTENNA_output596_A (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_output666_A (.DIODE(net994));
 sky130_fd_sc_hd__diode_2 ANTENNA_output665_A (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_output660_A (.DIODE(net996));
 sky130_fd_sc_hd__diode_2 ANTENNA_output658_A (.DIODE(net997));
 sky130_fd_sc_hd__diode_2 ANTENNA_output655_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_output650_A (.DIODE(net999));
 sky130_fd_sc_hd__diode_2 ANTENNA_output649_A (.DIODE(net1000));
 sky130_fd_sc_hd__diode_2 ANTENNA_output647_A (.DIODE(net1001));
 sky130_fd_sc_hd__diode_2 ANTENNA_output646_A (.DIODE(net1002));
 sky130_fd_sc_hd__diode_2 ANTENNA_output645_A (.DIODE(net1003));
 sky130_fd_sc_hd__diode_2 ANTENNA_output643_A (.DIODE(net1004));
 sky130_fd_sc_hd__diode_2 ANTENNA_output642_A (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA_output640_A (.DIODE(net1006));
 sky130_fd_sc_hd__diode_2 ANTENNA_output639_A (.DIODE(net1007));
 sky130_fd_sc_hd__diode_2 ANTENNA_output637_A (.DIODE(net1008));
 sky130_fd_sc_hd__diode_2 ANTENNA_output636_A (.DIODE(net1009));
 sky130_fd_sc_hd__diode_2 ANTENNA_output634_A (.DIODE(net1010));
 sky130_fd_sc_hd__diode_2 ANTENNA_output631_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_output629_A (.DIODE(net1012));
 sky130_fd_sc_hd__diode_2 ANTENNA__0544__A (.DIODE(net1013));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1013_A (.DIODE(net1014));
 sky130_fd_sc_hd__diode_2 ANTENNA__0543__A (.DIODE(net1015));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1015_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__0542__A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1017_A (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__0541__A (.DIODE(net1019));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1019_A (.DIODE(net1020));
 sky130_fd_sc_hd__diode_2 ANTENNA__0540__A (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1021_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1022_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__0539__A (.DIODE(net1024));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1024_A (.DIODE(net1025));
 sky130_fd_sc_hd__diode_2 ANTENNA__0538__A (.DIODE(net1026));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1026_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__0537__A (.DIODE(net1028));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1028_A (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1030_A (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA__0535__A (.DIODE(net1032));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1032_A (.DIODE(net1033));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1033_A (.DIODE(net1034));
 sky130_fd_sc_hd__diode_2 ANTENNA__0534__A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__0533__A (.DIODE(net1036));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1036_A (.DIODE(net1037));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1037_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__0532__A (.DIODE(net1039));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1039_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1040_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA__0531__A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1042_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA__0530__A (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1044_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__0529__A (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1046_A (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1047_A (.DIODE(net1048));
 sky130_fd_sc_hd__diode_2 ANTENNA__0528__A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1049_A (.DIODE(net1050));
 sky130_fd_sc_hd__diode_2 ANTENNA__0527__A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1051_A (.DIODE(net1052));
 sky130_fd_sc_hd__diode_2 ANTENNA__0526__A (.DIODE(net1053));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1053_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1054_A (.DIODE(net1055));
 sky130_fd_sc_hd__diode_2 ANTENNA__0525__A (.DIODE(net1056));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1056_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1057_A (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__0524__A (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1059_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__0523__A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1061_A (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__0522__A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1063_A (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1064_A (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1065_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__0521__A (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1067_A (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1068_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA__0520__A (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1070_A (.DIODE(net1071));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1071_A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__0519__A (.DIODE(net1073));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1073_A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__0518__A (.DIODE(net1075));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1075_A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__0517__A (.DIODE(net1077));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1077_A (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__0516__A (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__0515__A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__A (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1081_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__0547__A (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__0546__A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1084_A (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__0545__A (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA_output833_A (.DIODE(net1087));
 sky130_fd_sc_hd__diode_2 ANTENNA_output832_A (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA_output826_A (.DIODE(net1089));
 sky130_fd_sc_hd__diode_2 ANTENNA_output817_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_output786_A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA_output779_A (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA_output766_A (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA_output791_A (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA_output719_A (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA_output473_A (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA_output471_A (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA_output469_A (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA_output467_A (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_A (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output589_A (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output588_A (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1103_A (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output586_A (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output585_A (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output584_A (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA_output583_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output582_A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output581_A (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output578_A (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output576_A (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output575_A (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output573_A (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output572_A (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output571_A (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output570_A (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output569_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output533_A (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output525_A (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output518_A (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output517_A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1122_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output516_A (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1124_A (.DIODE(net1125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output515_A (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output512_A (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA_output511_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output510_A (.DIODE(net1129));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1129_A (.DIODE(net1130));
 sky130_fd_sc_hd__diode_2 ANTENNA_output509_A (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA_output503_A (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output501_A (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1133_A (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA_output498_A (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1135_A (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output495_A (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output494_A (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output590_A (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA_output568_A (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_output557_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_output546_A (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA_output535_A (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA_output524_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_output513_A (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_output502_A (.DIODE(net1146));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1146_A (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_output463_A (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA_output937_A (.DIODE(net1149));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1149_A (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA_output936_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1151_A (.DIODE(net1152));
 sky130_fd_sc_hd__diode_2 ANTENNA_output934_A (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1153_A (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1154_A (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output933_A (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1156_A (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1157_A (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA_output932_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1159_A (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1160_A (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output931_A (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1162_A (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1163_A (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA_output930_A (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1165_A (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1166_A (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA_output929_A (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1168_A (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1169_A (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_output928_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1171_A (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1172_A (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA_output927_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1174_A (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1175_A (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA_output926_A (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1177_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1178_A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output925_A (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1180_A (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1181_A (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output923_A (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1183_A (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1184_A (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output922_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1186_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output921_A (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1188_A (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1189_A (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output920_A (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1191_A (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1192_A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output919_A (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1194_A (.DIODE(net1195));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1195_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output918_A (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1197_A (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1198_A (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output917_A (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1200_A (.DIODE(net1201));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1201_A (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1202_A (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output916_A (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1204_A (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1205_A (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1206_A (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output915_A (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1208_A (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1209_A (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output914_A (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1211_A (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1212_A (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output944_A (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1214_A (.DIODE(net1215));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1215_A (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA_output943_A (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1217_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1218_A (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1219_A (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA_output942_A (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1221_A (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1222_A (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA_output941_A (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1224_A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1225_A (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1226_A (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output940_A (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1228_A (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1229_A (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1230_A (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA_output939_A (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1232_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1233_A (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA_output938_A (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1235_A (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1236_A (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA_output935_A (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1238_A (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1239_A (.DIODE(net1240));
 sky130_fd_sc_hd__diode_2 ANTENNA_output924_A (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1241_A (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1242_A (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA_output913_A (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1244_A (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1245_A (.DIODE(net1246));
 sky130_fd_sc_hd__diode_2 ANTENNA_output872_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1247_A (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA_output871_A (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1249_A (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA_output869_A (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA_output868_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_output867_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_output866_A (.DIODE(net1254));
 sky130_fd_sc_hd__diode_2 ANTENNA_output863_A (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1255_A (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output862_A (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1257_A (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1258_A (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA_output860_A (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1260_A (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA_output858_A (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA_output856_A (.DIODE(net1263));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1263_A (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1264_A (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA_output854_A (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA_output853_A (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1267_A (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1268_A (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA_output852_A (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1270_A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output851_A (.DIODE(net1272));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1272_A (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA_output850_A (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1274_A (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1275_A (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA_output849_A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1277_A (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1278_A (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1279_A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA_output879_A (.DIODE(net1281));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1281_A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1282_A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_output876_A (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1284_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1285_A (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA_output875_A (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1287_A (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output873_A (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output859_A (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output848_A (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output948_A (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1292_A (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1293_A (.DIODE(net1294));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1294_A (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output947_A (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1296_A (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1297_A (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1298_A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1299_A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA_output946_A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1301_A (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1302_A (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1303_A (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1304_A (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output945_A (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1306_A (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1307_A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1308_A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1309_A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA_output950_A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1311_A (.DIODE(net1312));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1312_A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1313_A (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA_output949_A (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1315_A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1316_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1317_A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA_output880_A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1319_A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1320_A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA_output955_A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1322_A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1323_A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1324_A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[4]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[7]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[2]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[8]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA_user_wb_ack_gate_B (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[1]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[0]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[6]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[5]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[19]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[10]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[17]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[12]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[15]_B  (.DIODE(net1326));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1326_A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[3]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[11]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[20]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[18]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[9]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[13]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[16]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[28]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_wb_dat_gates[27]_B  (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_user_to_mprj_in_gates[105]_B  (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__1460__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__1458__A (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__1456__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1331_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1337_A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__A (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1340_A (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1342_A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__A (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1344_A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1346_A (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__1388__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__A (.DIODE(net1349));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1349_A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__1382__A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1351_A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1353_A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__1376__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1355_A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__A (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1359_A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__A (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__1348__A (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__A (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__A (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__A (.DIODE(net1366));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__A (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__A (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__A (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1369_A (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__A (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1372_A (.DIODE(net1373));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__A (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__1322__A (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1375_A (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__A (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__A (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__1316__A (.DIODE(net1379));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1379_A (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__A (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__A (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1383_A (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__A (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__A (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__A (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__A (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1388_A (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__A (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__1298__A (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__A (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__1294__A (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1393_A (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__1292__A (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1395_A (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__A (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1397_A (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__A (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1399_A (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__A (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__1282__A (.DIODE(net1403));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__A (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__A (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__A (.DIODE(net1406));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__A (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__A (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__A (.DIODE(net1411));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__A (.DIODE(net1412));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__A (.DIODE(net1413));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__A (.DIODE(net1414));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__A (.DIODE(net1415));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1415_A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__A (.DIODE(net1417));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1417_A (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__A (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1419_A (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__A (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__A (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1422_A (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__1220__A (.DIODE(net1424));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1424_A (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__A (.DIODE(net1426));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1426_A (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1428_A (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__A (.DIODE(net1430));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1430_A (.DIODE(net1431));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__A (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1432_A (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1433_A (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__A (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1435_A (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1436_A (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__A (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1438_A (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1440_A (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__A (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1447_A (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A (.DIODE(net1449));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1449_A (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__A (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1451_A (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1453_A (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1454_A (.DIODE(net1455));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1456_A (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1458_A (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1460_A (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1462_A (.DIODE(net1463));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1464_A (.DIODE(net1465));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1466_A (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1467_A (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__A (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1469_A (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A (.DIODE(net1471));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1471_A (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A (.DIODE(net1473));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1473_A (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A (.DIODE(net1479));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1480_A (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__A (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1483_A (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__A (.DIODE(net1486));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__A (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__1062__A (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1493_A (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__1060__A (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__A (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1496_A (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__A (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__A (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1499_A (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__A (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__A (.DIODE(net1503));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1503_A (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__A (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__A (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__A (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__A (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__A (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__A (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1513_A (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1514_A (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1516_A (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__1006__A (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1518_A (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__A (.DIODE(net1520));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1520_A (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__A (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1526_A (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1528_A (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__A (.DIODE(net1531));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__A (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1533_A (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__A (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA__0960__A (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__A (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__0906__A (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__0890__A (.DIODE(net1543));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1543_A (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1544_A (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__0888__A (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1546_A (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__0884__A (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__0880__A (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__A (.DIODE(net1552));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__0820__A (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1556_A (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1558_A (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1559_A (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1561_A (.DIODE(net1562));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1562_A (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__0812__A (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1564_A (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1565_A (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A (.DIODE(net1567));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1567_A (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1568_A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__A (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1570_A (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__0806__A (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1572_A (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1573_A (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__A (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1575_A (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__A (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1577_A (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1578_A (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__A (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1580_A (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__A (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1582_A (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1583_A (.DIODE(net1584));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1585_A (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1586_A (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1588_A (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1589_A (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__A (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1591_A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1592_A (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1594_A (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1595_A (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__A (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1597_A (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1598_A (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__A (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1600_A (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1602_A (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1603_A (.DIODE(net1604));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__A (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1605_A (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1607_A (.DIODE(net1608));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__A (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1609_A (.DIODE(net1610));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1610_A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__A (.DIODE(net1612));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1612_A (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1613_A (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1615_A (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__A (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1617_A (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1618_A (.DIODE(net1619));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__A (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA__0766__A (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1621_A (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__A (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1623_A (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__A (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1625_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__A (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1627_A (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__A (.DIODE(net1629));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__C (.DIODE(net1633));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__C (.DIODE(net1634));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__C (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__C (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__C (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__C (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__C (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__C (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__C (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__C (.DIODE(net1642));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__C (.DIODE(net1643));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__C (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__C (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__C (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__C (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__C (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__B (.DIODE(net1649));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__B (.DIODE(net1650));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__B (.DIODE(net1651));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__B (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1652_A (.DIODE(net1653));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__B (.DIODE(net1654));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1654_A (.DIODE(net1655));
 sky130_fd_sc_hd__diode_2 ANTENNA__0967__B (.DIODE(net1656));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1656_A (.DIODE(net1657));
 sky130_fd_sc_hd__diode_2 ANTENNA__0965__B (.DIODE(net1658));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1658_A (.DIODE(net1659));
 sky130_fd_sc_hd__diode_2 ANTENNA__0963__B (.DIODE(net1660));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1660_A (.DIODE(net1661));
 sky130_fd_sc_hd__diode_2 ANTENNA__0961__B (.DIODE(net1662));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1662_A (.DIODE(net1663));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1663_A (.DIODE(net1664));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__B (.DIODE(net1665));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1665_A (.DIODE(net1666));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__B (.DIODE(net1667));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1667_A (.DIODE(net1668));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__B (.DIODE(net1669));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (.DIODE(net1670));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__B (.DIODE(net1671));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__C (.DIODE(net1672));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__B (.DIODE(net1673));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__B (.DIODE(net1674));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1674_A (.DIODE(net1675));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__B (.DIODE(net1676));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1676_A (.DIODE(net1677));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (.DIODE(net1678));
 sky130_fd_sc_hd__diode_2 ANTENNA__0957__B (.DIODE(net1679));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1679_A (.DIODE(net1680));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1680_A (.DIODE(net1681));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__B (.DIODE(net1682));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (.DIODE(net1683));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (.DIODE(net1684));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__B (.DIODE(net1685));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1685_A (.DIODE(net1686));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (.DIODE(net1687));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1687_A (.DIODE(net1688));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__B (.DIODE(net1689));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1689_A (.DIODE(net1690));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__B (.DIODE(net1691));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__B (.DIODE(net1692));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__B (.DIODE(net1693));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__B (.DIODE(net1694));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1694_A (.DIODE(net1695));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1695_A (.DIODE(net1696));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__B (.DIODE(net1697));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1697_A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1698_A (.DIODE(net1699));
 sky130_fd_sc_hd__diode_2 ANTENNA__0909__B (.DIODE(net1700));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1700_A (.DIODE(net1701));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1701_A (.DIODE(net1702));
 sky130_fd_sc_hd__diode_2 ANTENNA__0907__B (.DIODE(net1703));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1703_A (.DIODE(net1704));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1704_A (.DIODE(net1705));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1705_A (.DIODE(net1706));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1706_A (.DIODE(net1707));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__B (.DIODE(net1708));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1708_A (.DIODE(net1709));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1709_A (.DIODE(net1710));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1710_A (.DIODE(net1711));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1711_A (.DIODE(net1712));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1712_A (.DIODE(net1713));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__B (.DIODE(net1714));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1714_A (.DIODE(net1715));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1715_A (.DIODE(net1716));
 sky130_fd_sc_hd__diode_2 ANTENNA__0901__B (.DIODE(net1717));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1717_A (.DIODE(net1718));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1718_A (.DIODE(net1719));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1719_A (.DIODE(net1720));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__B (.DIODE(net1721));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1721_A (.DIODE(net1722));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1722_A (.DIODE(net1723));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1723_A (.DIODE(net1724));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1724_A (.DIODE(net1725));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__B (.DIODE(net1726));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1726_A (.DIODE(net1727));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1727_A (.DIODE(net1728));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1728_A (.DIODE(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__B (.DIODE(net1730));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1730_A (.DIODE(net1731));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1731_A (.DIODE(net1732));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1732_A (.DIODE(net1733));
 sky130_fd_sc_hd__diode_2 ANTENNA__0951__B (.DIODE(net1734));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1734_A (.DIODE(net1735));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1735_A (.DIODE(net1736));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1736_A (.DIODE(net1737));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__B (.DIODE(net1738));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1738_A (.DIODE(net1739));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1739_A (.DIODE(net1740));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1740_A (.DIODE(net1741));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1741_A (.DIODE(net1742));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__C (.DIODE(net1743));
 sky130_fd_sc_hd__diode_2 ANTENNA__0949__B (.DIODE(net1744));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1744_A (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1745_A (.DIODE(net1746));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1746_A (.DIODE(net1747));
 sky130_fd_sc_hd__diode_2 ANTENNA__0947__B (.DIODE(net1748));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1748_A (.DIODE(net1749));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1749_A (.DIODE(net1750));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1750_A (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__B (.DIODE(net1752));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1752_A (.DIODE(net1753));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1753_A (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1754_A (.DIODE(net1755));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1755_A (.DIODE(net1756));
 sky130_fd_sc_hd__diode_2 ANTENNA__0943__B (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1757_A (.DIODE(net1758));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1758_A (.DIODE(net1759));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1759_A (.DIODE(net1760));
 sky130_fd_sc_hd__diode_2 ANTENNA__0941__B (.DIODE(net1761));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1761_A (.DIODE(net1762));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1762_A (.DIODE(net1763));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1763_A (.DIODE(net1764));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1764_A (.DIODE(net1765));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__B (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1766_A (.DIODE(net1767));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1767_A (.DIODE(net1768));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1768_A (.DIODE(net1769));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1769_A (.DIODE(net1770));
 sky130_fd_sc_hd__diode_2 ANTENNA__0937__B (.DIODE(net1771));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1771_A (.DIODE(net1772));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1772_A (.DIODE(net1773));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1773_A (.DIODE(net1774));
 sky130_fd_sc_hd__diode_2 ANTENNA__0935__B (.DIODE(net1775));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1775_A (.DIODE(net1776));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1776_A (.DIODE(net1777));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__B (.DIODE(net1778));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1778_A (.DIODE(net1779));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1779_A (.DIODE(net1780));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1780_A (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1781_A (.DIODE(net1782));
 sky130_fd_sc_hd__diode_2 ANTENNA__0931__B (.DIODE(net1783));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1783_A (.DIODE(net1784));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1784_A (.DIODE(net1785));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__B (.DIODE(net1786));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1786_A (.DIODE(net1787));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1787_A (.DIODE(net1788));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1788_A (.DIODE(net1789));
 sky130_fd_sc_hd__diode_2 ANTENNA__0929__B (.DIODE(net1790));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1790_A (.DIODE(net1791));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1791_A (.DIODE(net1792));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1792_A (.DIODE(net1793));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__B (.DIODE(net1794));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1794_A (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1795_A (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1796_A (.DIODE(net1797));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1797_A (.DIODE(net1798));
 sky130_fd_sc_hd__diode_2 ANTENNA__0925__B (.DIODE(net1799));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1799_A (.DIODE(net1800));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1800_A (.DIODE(net1801));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__B (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1802_A (.DIODE(net1803));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1803_A (.DIODE(net1804));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1804_A (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1805_A (.DIODE(net1806));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__B (.DIODE(net1807));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1807_A (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1808_A (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1809_A (.DIODE(net1810));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1810_A (.DIODE(net1811));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__B (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1812_A (.DIODE(net1813));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1813_A (.DIODE(net1814));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__B (.DIODE(net1815));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1815_A (.DIODE(net1816));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1816_A (.DIODE(net1817));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__B (.DIODE(net1818));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1818_A (.DIODE(net1819));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1819_A (.DIODE(net1820));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1820_A (.DIODE(net1821));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__B (.DIODE(net1822));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1822_A (.DIODE(net1823));
 sky130_fd_sc_hd__diode_2 ANTENNA__0911__B (.DIODE(net1824));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1824_A (.DIODE(net1825));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__B (.DIODE(net1826));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1826_A (.DIODE(net1827));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1827_A (.DIODE(net1828));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1828_A (.DIODE(net1829));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1829_A (.DIODE(net1830));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A (.DIODE(net1831));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1831_A (.DIODE(net1832));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__A_N (.DIODE(net1832));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__A (.DIODE(net1833));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1833_A (.DIODE(net1834));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A (.DIODE(net1835));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__A (.DIODE(net1836));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1836_A (.DIODE(net1837));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__A_N (.DIODE(net1837));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__A (.DIODE(net1838));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A (.DIODE(net1839));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__A (.DIODE(net1840));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__A (.DIODE(net1841));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1841_A (.DIODE(net1842));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__A_N (.DIODE(net1842));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__A_N (.DIODE(net1843));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__A (.DIODE(net1843));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1843_A (.DIODE(net1844));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__A_N (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__A (.DIODE(net1845));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1845_A (.DIODE(net1846));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__A_N (.DIODE(net1847));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__A (.DIODE(net1847));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1847_A (.DIODE(net1848));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__A (.DIODE(net1849));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A_N (.DIODE(net1849));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1849_A (.DIODE(net1850));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__A_N (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__A (.DIODE(net1851));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1851_A (.DIODE(net1852));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__A_N (.DIODE(net1853));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__A (.DIODE(net1853));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1853_A (.DIODE(net1854));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__A_N (.DIODE(net1855));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A (.DIODE(net1855));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1855_A (.DIODE(net1856));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__A_N (.DIODE(net1857));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__A (.DIODE(net1857));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1857_A (.DIODE(net1858));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__A (.DIODE(net1859));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1859_A (.DIODE(net1860));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A_N (.DIODE(net1860));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__A_N (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__A (.DIODE(net1861));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1861_A (.DIODE(net1862));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__A_N (.DIODE(net1863));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__A (.DIODE(net1863));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1863_A (.DIODE(net1864));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (.DIODE(net1865));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__A_N (.DIODE(net1865));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1865_A (.DIODE(net1866));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__A (.DIODE(net1867));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A_N (.DIODE(net1867));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__A_N (.DIODE(net1868));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__A (.DIODE(net1868));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1868_A (.DIODE(net1869));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__A (.DIODE(net1870));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A_N (.DIODE(net1870));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A_N (.DIODE(net1871));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A_N (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__A (.DIODE(net1872));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__A (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A_N (.DIODE(net1873));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__A (.DIODE(net1874));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A_N (.DIODE(net1874));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__A_N (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A (.DIODE(net1875));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__A_N (.DIODE(net1876));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (.DIODE(net1876));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__A (.DIODE(net1877));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1877_A (.DIODE(net1878));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__A_N (.DIODE(net1878));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__A (.DIODE(net1879));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A (.DIODE(net1880));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1880_A (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__A_N (.DIODE(net1882));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__A (.DIODE(net1883));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__A (.DIODE(net1884));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__A_N (.DIODE(net1884));
 sky130_fd_sc_hd__diode_2 ANTENNA__1397__A (.DIODE(net1885));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A_N (.DIODE(net1885));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__A (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__A_N (.DIODE(net1886));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__A (.DIODE(net1887));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1887_A (.DIODE(net1888));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__A_N (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__A_N (.DIODE(net1890));
 sky130_fd_sc_hd__diode_2 ANTENNA__1391__A (.DIODE(net1890));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__A_N (.DIODE(net1891));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__A (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1892_A (.DIODE(net1893));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__C (.DIODE(net1894));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A_N (.DIODE(net1895));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__A (.DIODE(net1895));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__A_N (.DIODE(net1896));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__A (.DIODE(net1897));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1896_A (.DIODE(net1898));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__A (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__A_N (.DIODE(net1899));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__A (.DIODE(net1900));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A_N (.DIODE(net1900));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__A (.DIODE(net1901));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A_N (.DIODE(net1902));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A (.DIODE(net1903));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__A (.DIODE(net1904));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1904_A (.DIODE(net1905));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1905_A (.DIODE(net1906));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__C (.DIODE(net1907));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A (.DIODE(net1908));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1908_A (.DIODE(net1909));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A_N (.DIODE(net1910));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (.DIODE(net1911));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1911_A (.DIODE(net1912));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__A_N (.DIODE(net1913));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__A (.DIODE(net1914));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1914_A (.DIODE(net1915));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__A (.DIODE(net1916));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__A_N (.DIODE(net1916));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__A (.DIODE(net1917));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__A_N (.DIODE(net1918));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__C (.DIODE(net1919));
 sky130_fd_sc_hd__diode_2 ANTENNA__1349__A (.DIODE(net1920));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1920_A (.DIODE(net1921));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__A (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__A_N (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__C (.DIODE(net1923));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A_N (.DIODE(net1924));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__A (.DIODE(net1925));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__A (.DIODE(net1926));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A_N (.DIODE(net1926));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__A (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__A_N (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__A (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A_N (.DIODE(net1929));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A_N (.DIODE(net1930));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1930_A (.DIODE(net1931));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1931_A (.DIODE(net1932));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1932_A (.DIODE(net1933));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1933_A (.DIODE(net1934));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1934_A (.DIODE(net1935));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1935_A (.DIODE(net1936));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__A_N (.DIODE(net1937));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__A_N (.DIODE(net1938));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__A_N (.DIODE(net1939));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A_N (.DIODE(net1940));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A (.DIODE(net1940));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__A_N (.DIODE(net1941));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A (.DIODE(net1942));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A (.DIODE(net1943));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (.DIODE(net1944));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__A_N (.DIODE(net1944));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__A (.DIODE(net1945));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1945_A (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__A_N (.DIODE(net1946));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A (.DIODE(net1947));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A (.DIODE(net1948));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__A_N (.DIODE(net1948));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__C (.DIODE(net1949));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A (.DIODE(net1950));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__A_N (.DIODE(net1950));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A (.DIODE(net1951));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__A_N (.DIODE(net1951));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A (.DIODE(net1952));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__A_N (.DIODE(net1952));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A (.DIODE(net1953));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1953_A (.DIODE(net1954));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__A_N (.DIODE(net1954));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A (.DIODE(net1955));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__A_N (.DIODE(net1955));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__A (.DIODE(net1956));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__A_N (.DIODE(net1956));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A (.DIODE(net1957));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__A_N (.DIODE(net1957));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (.DIODE(net1958));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__A_N (.DIODE(net1958));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A (.DIODE(net1959));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__C (.DIODE(net1960));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A (.DIODE(net1961));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__A_N (.DIODE(net1961));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A (.DIODE(net1962));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A (.DIODE(net1963));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1963_A (.DIODE(net1964));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__A (.DIODE(net1965));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1965_A (.DIODE(net1966));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A (.DIODE(net1967));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A (.DIODE(net1968));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__A (.DIODE(net1969));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1969_A (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__A_N (.DIODE(net1970));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A (.DIODE(net1971));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__A (.DIODE(net1972));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1972_A (.DIODE(net1973));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__A_N (.DIODE(net1973));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__B (.DIODE(net1974));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__B (.DIODE(net1975));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1975_A (.DIODE(net1976));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__B (.DIODE(net1977));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1977_A (.DIODE(net1978));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__B (.DIODE(net1979));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__B (.DIODE(net1980));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__B (.DIODE(net1981));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1981_A (.DIODE(net1982));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__B (.DIODE(net1983));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1983_A (.DIODE(net1984));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__B (.DIODE(net1985));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1985_A (.DIODE(net1986));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B (.DIODE(net1987));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__B (.DIODE(net1988));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__B (.DIODE(net1989));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__B (.DIODE(net1990));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__B (.DIODE(net1991));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__B (.DIODE(net1992));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B (.DIODE(net1993));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__B (.DIODE(net1994));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (.DIODE(net1995));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__B (.DIODE(net1996));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__B (.DIODE(net1997));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__B (.DIODE(net1998));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__B (.DIODE(net1999));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__B (.DIODE(net2000));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__B (.DIODE(net2001));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__B (.DIODE(net2002));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B (.DIODE(net2003));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__B (.DIODE(net2004));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__B (.DIODE(net2005));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__B (.DIODE(net2006));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__C (.DIODE(net2007));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__B (.DIODE(net2008));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__B (.DIODE(net2009));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__B (.DIODE(net2010));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__B (.DIODE(net2011));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__B (.DIODE(net2012));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__B (.DIODE(net2013));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2013_A (.DIODE(net2014));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__B (.DIODE(net2015));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__B (.DIODE(net2016));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__B (.DIODE(net2017));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2017_A (.DIODE(net2018));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__B (.DIODE(net2019));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__B (.DIODE(net2020));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2020_A (.DIODE(net2021));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__B (.DIODE(net2022));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__B (.DIODE(net2023));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__B (.DIODE(net2024));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__B (.DIODE(net2025));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__B (.DIODE(net2026));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__B (.DIODE(net2027));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2027_A (.DIODE(net2028));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__C (.DIODE(net2029));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__C (.DIODE(net2030));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2030_A (.DIODE(net2031));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2031_A (.DIODE(net2032));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__C (.DIODE(net2033));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2033_A (.DIODE(net2034));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2034_A (.DIODE(net2035));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__C (.DIODE(net2036));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2036_A (.DIODE(net2037));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__C (.DIODE(net2038));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2038_A (.DIODE(net2039));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__C (.DIODE(net2040));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2040_A (.DIODE(net2041));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2041_A (.DIODE(net2042));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__C (.DIODE(net2043));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2043_A (.DIODE(net2044));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2044_A (.DIODE(net2045));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__C (.DIODE(net2046));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2046_A (.DIODE(net2047));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__C (.DIODE(net2048));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2048_A (.DIODE(net2049));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2049_A (.DIODE(net2050));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__C (.DIODE(net2051));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__C (.DIODE(net2052));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2052_A (.DIODE(net2053));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__C (.DIODE(net2054));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2054_A (.DIODE(net2055));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2055_A (.DIODE(net2056));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__C (.DIODE(net2057));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2057_A (.DIODE(net2058));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__C (.DIODE(net2059));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__C (.DIODE(net2060));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2060_A (.DIODE(net2061));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__C (.DIODE(net2062));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__C (.DIODE(net2063));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__C (.DIODE(net2064));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2064_A (.DIODE(net2065));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__B (.DIODE(net2066));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2066_A (.DIODE(net2067));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2067_A (.DIODE(net2068));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2068_A (.DIODE(net2069));
 sky130_fd_sc_hd__diode_2 ANTENNA_output952_A (.DIODE(net2070));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2070_A (.DIODE(net2071));
 sky130_fd_sc_hd__diode_2 ANTENNA_output954_A (.DIODE(net2072));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2072_A (.DIODE(net2073));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2073_A (.DIODE(net2074));
 sky130_fd_sc_hd__diode_2 ANTENNA__0889__A (.DIODE(net2075));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2075_A (.DIODE(net2076));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2076_A (.DIODE(net2077));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__B (.DIODE(net2078));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2078_A (.DIODE(net2079));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2079_A (.DIODE(net2080));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__B (.DIODE(net2081));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2081_A (.DIODE(net2082));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2082_A (.DIODE(net2083));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__B (.DIODE(net2084));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2084_A (.DIODE(net2085));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__B (.DIODE(net2086));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2086_A (.DIODE(net2087));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2087_A (.DIODE(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__B (.DIODE(net2089));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2089_A (.DIODE(net2090));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2090_A (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__B (.DIODE(net2092));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2092_A (.DIODE(net2093));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2093_A (.DIODE(net2094));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2094_A (.DIODE(net2095));
 sky130_fd_sc_hd__diode_2 ANTENNA__1057__B (.DIODE(net2096));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2096_A (.DIODE(net2097));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2097_A (.DIODE(net2098));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__B (.DIODE(net2099));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2099_A (.DIODE(net2100));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2100_A (.DIODE(net2101));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2101_A (.DIODE(net2102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__B (.DIODE(net2103));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2103_A (.DIODE(net2104));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2104_A (.DIODE(net2105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1051__B (.DIODE(net2106));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2106_A (.DIODE(net2107));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2107_A (.DIODE(net2108));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__A (.DIODE(net2109));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2109_A (.DIODE(net2110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(net2111));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2111_A (.DIODE(net2112));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2112_A (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2113_A (.DIODE(net2114));
 sky130_fd_sc_hd__diode_2 ANTENNA__1047__B (.DIODE(net2115));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2115_A (.DIODE(net2116));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2116_A (.DIODE(net2117));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2117_A (.DIODE(net2118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B (.DIODE(net2119));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2119_A (.DIODE(net2120));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2120_A (.DIODE(net2121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B (.DIODE(net2122));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2122_A (.DIODE(net2123));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2123_A (.DIODE(net2124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__B (.DIODE(net2125));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2125_A (.DIODE(net2126));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2126_A (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2127_A (.DIODE(net2128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B (.DIODE(net2129));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2129_A (.DIODE(net2130));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2130_A (.DIODE(net2131));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2131_A (.DIODE(net2132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B (.DIODE(net2133));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2133_A (.DIODE(net2134));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2134_A (.DIODE(net2135));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2135_A (.DIODE(net2136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B (.DIODE(net2137));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2137_A (.DIODE(net2138));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2138_A (.DIODE(net2139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__B (.DIODE(net2140));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2140_A (.DIODE(net2141));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2141_A (.DIODE(net2142));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2142_A (.DIODE(net2143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B (.DIODE(net2144));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2144_A (.DIODE(net2145));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2145_A (.DIODE(net2146));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2146_A (.DIODE(net2147));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A (.DIODE(net2148));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2148_A (.DIODE(net2149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__B (.DIODE(net2150));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2150_A (.DIODE(net2151));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2151_A (.DIODE(net2152));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__B (.DIODE(net2153));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2153_A (.DIODE(net2154));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2154_A (.DIODE(net2155));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__B (.DIODE(net2156));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2156_A (.DIODE(net2157));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2157_A (.DIODE(net2158));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B (.DIODE(net2159));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2159_A (.DIODE(net2160));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2160_A (.DIODE(net2161));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__B (.DIODE(net2162));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2162_A (.DIODE(net2163));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2163_A (.DIODE(net2164));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__B (.DIODE(net2165));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2165_A (.DIODE(net2166));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2166_A (.DIODE(net2167));
 sky130_fd_sc_hd__diode_2 ANTENNA__1017__A (.DIODE(net2168));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__A (.DIODE(net2169));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (.DIODE(net2170));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2170_A (.DIODE(net2171));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__A (.DIODE(net2172));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2172_A (.DIODE(net2173));
 sky130_fd_sc_hd__diode_2 ANTENNA__0883__A (.DIODE(net2174));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2174_A (.DIODE(net2175));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A (.DIODE(net2176));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2176_A (.DIODE(net2177));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2177_A (.DIODE(net2178));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2178_A (.DIODE(net2179));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__A (.DIODE(net2180));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2180_A (.DIODE(net2181));
 sky130_fd_sc_hd__diode_2 ANTENNA__1005__A (.DIODE(net2182));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2182_A (.DIODE(net2183));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2183_A (.DIODE(net2184));
 sky130_fd_sc_hd__diode_2 ANTENNA__1003__A (.DIODE(net2185));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2185_A (.DIODE(net2186));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2186_A (.DIODE(net2187));
 sky130_fd_sc_hd__diode_2 ANTENNA__1001__A (.DIODE(net2188));
 sky130_fd_sc_hd__diode_2 ANTENNA__0999__A (.DIODE(net2189));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__A (.DIODE(net2190));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__A (.DIODE(net2191));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2191_A (.DIODE(net2192));
 sky130_fd_sc_hd__diode_2 ANTENNA__0993__A (.DIODE(net2193));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__A (.DIODE(net2194));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__A (.DIODE(net2195));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__A (.DIODE(net2196));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2196_A (.DIODE(net2197));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (.DIODE(net2198));
 sky130_fd_sc_hd__diode_2 ANTENNA__0983__A (.DIODE(net2199));
 sky130_fd_sc_hd__diode_2 ANTENNA__0981__A (.DIODE(net2200));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2200_A (.DIODE(net2201));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(net2202));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2202_A (.DIODE(net2203));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__A (.DIODE(net2204));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2204_A (.DIODE(net2205));
 sky130_fd_sc_hd__diode_2 ANTENNA__0975__A (.DIODE(net2206));
 sky130_fd_sc_hd__diode_2 ANTENNA__0973__A (.DIODE(net2207));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (.DIODE(net2208));
 sky130_fd_sc_hd__diode_2 ANTENNA__0969__A (.DIODE(net2209));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(net2210));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2210_A (.DIODE(net2211));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2211_A (.DIODE(net2212));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2212_A (.DIODE(net2213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output951_A (.DIODE(net2214));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2214_A (.DIODE(net2215));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2215_A (.DIODE(net2216));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2216_A (.DIODE(net2217));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(net2218));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2218_A (.DIODE(net2219));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2219_A (.DIODE(net2220));
 sky130_fd_sc_hd__diode_2 ANTENNA__0865__A (.DIODE(net2221));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2221_A (.DIODE(net2222));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2222_A (.DIODE(net2223));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2223_A (.DIODE(net2224));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__A (.DIODE(net2225));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2225_A (.DIODE(net2226));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2226_A (.DIODE(net2227));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2227_A (.DIODE(net2228));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(net2229));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2229_A (.DIODE(net2230));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A (.DIODE(net2231));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2231_A (.DIODE(net2232));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2232_A (.DIODE(net2233));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (.DIODE(net2234));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2234_A (.DIODE(net2235));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2235_A (.DIODE(net2236));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A (.DIODE(net2237));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2237_A (.DIODE(net2238));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2238_A (.DIODE(net2239));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__A (.DIODE(net2240));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2240_A (.DIODE(net2241));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2241_A (.DIODE(net2242));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__A (.DIODE(net2243));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2243_A (.DIODE(net2244));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2244_A (.DIODE(net2245));
 sky130_fd_sc_hd__diode_2 ANTENNA__0849__A (.DIODE(net2246));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2246_A (.DIODE(net2247));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2247_A (.DIODE(net2248));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__A (.DIODE(net2249));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2249_A (.DIODE(net2250));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2250_A (.DIODE(net2251));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2251_A (.DIODE(net2252));
 sky130_fd_sc_hd__diode_2 ANTENNA__0959__A (.DIODE(net2253));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A (.DIODE(net2254));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2254_A (.DIODE(net2255));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A (.DIODE(net2256));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2256_A (.DIODE(net2257));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2257_A (.DIODE(net2258));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__A (.DIODE(net2259));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2259_A (.DIODE(net2260));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2260_A (.DIODE(net2261));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__A (.DIODE(net2262));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2262_A (.DIODE(net2263));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__A (.DIODE(net2264));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2264_A (.DIODE(net2265));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2265_A (.DIODE(net2266));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2266_A (.DIODE(net2267));
 sky130_fd_sc_hd__diode_2 ANTENNA__0835__A (.DIODE(net2268));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2268_A (.DIODE(net2269));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__A (.DIODE(net2270));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2270_A (.DIODE(net2271));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2271_A (.DIODE(net2272));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__A (.DIODE(net2273));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2273_A (.DIODE(net2274));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2274_A (.DIODE(net2275));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__A (.DIODE(net2276));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2276_A (.DIODE(net2277));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2277_A (.DIODE(net2278));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__A (.DIODE(net2279));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2279_A (.DIODE(net2280));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__A (.DIODE(net2281));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2281_A (.DIODE(net2282));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2282_A (.DIODE(net2283));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__A (.DIODE(net2284));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2284_A (.DIODE(net2285));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2285_A (.DIODE(net2286));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__A (.DIODE(net2287));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2287_A (.DIODE(net2288));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2288_A (.DIODE(net2289));
 sky130_fd_sc_hd__diode_2 ANTENNA__0819__A (.DIODE(net2290));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2290_A (.DIODE(net2291));
 sky130_fd_sc_hd__diode_2 ANTENNA__0817__A (.DIODE(net2292));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__A (.DIODE(net2293));
 sky130_fd_sc_hd__diode_2 ANTENNA__0811__A (.DIODE(net2294));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A (.DIODE(net2295));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__A (.DIODE(net2296));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (.DIODE(net2297));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A (.DIODE(net2298));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__A (.DIODE(net2299));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (.DIODE(net2300));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__A (.DIODE(net2301));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__A (.DIODE(net2302));
 sky130_fd_sc_hd__diode_2 ANTENNA__0791__A (.DIODE(net2303));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (.DIODE(net2304));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__A (.DIODE(net2305));
 sky130_fd_sc_hd__diode_2 ANTENNA__0783__A (.DIODE(net2306));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A (.DIODE(net2307));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2307_A (.DIODE(net2308));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2308_A (.DIODE(net2309));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A (.DIODE(net2310));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__A (.DIODE(net2311));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A (.DIODE(net2312));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A (.DIODE(net2313));
 sky130_fd_sc_hd__diode_2 ANTENNA__0767__A (.DIODE(net2314));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2314_A (.DIODE(net2315));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2315_A (.DIODE(net2316));
 sky130_fd_sc_hd__diode_2 ANTENNA__0765__A (.DIODE(net2317));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__A (.DIODE(net2318));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__A (.DIODE(net2319));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A (.DIODE(net2320));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A (.DIODE(net2321));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2321_A (.DIODE(net2322));
 sky130_fd_sc_hd__diode_2 ANTENNA__0755__A (.DIODE(net2323));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2323_A (.DIODE(net2324));
 sky130_fd_sc_hd__diode_2 ANTENNA__0753__A (.DIODE(net2325));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2325_A (.DIODE(net2326));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__A (.DIODE(net2327));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__A (.DIODE(net2328));
 sky130_fd_sc_hd__diode_2 ANTENNA__0747__A (.DIODE(net2329));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A (.DIODE(net2330));
 sky130_fd_sc_hd__diode_2 ANTENNA__0727__A (.DIODE(net2331));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (.DIODE(net2332));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__A (.DIODE(net2333));
 sky130_fd_sc_hd__diode_2 ANTENNA__0715__A (.DIODE(net2334));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A (.DIODE(net2335));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A (.DIODE(net2336));
 sky130_fd_sc_hd__diode_2 ANTENNA__0709__A (.DIODE(net2337));
 sky130_fd_sc_hd__diode_2 ANTENNA__0707__A (.DIODE(net2338));
 sky130_fd_sc_hd__diode_2 ANTENNA__0703__A (.DIODE(net2339));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__A (.DIODE(net2340));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A (.DIODE(net2341));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__A (.DIODE(net2342));
 sky130_fd_sc_hd__diode_2 ANTENNA__0695__A (.DIODE(net2343));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A (.DIODE(net2344));
 sky130_fd_sc_hd__diode_2 ANTENNA__0691__A (.DIODE(net2345));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A (.DIODE(net2346));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A (.DIODE(net2347));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A (.DIODE(net2348));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (.DIODE(net2349));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2349_A (.DIODE(net2350));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (.DIODE(net2351));
 sky130_fd_sc_hd__diode_2 ANTENNA__0677__A (.DIODE(net2352));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2352_A (.DIODE(net2353));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A (.DIODE(net2354));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A (.DIODE(net2355));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2355_A (.DIODE(net2356));
 sky130_fd_sc_hd__diode_2 ANTENNA__0671__A (.DIODE(net2357));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A (.DIODE(net2358));
 sky130_fd_sc_hd__diode_2 ANTENNA__0667__A (.DIODE(net2359));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2359_A (.DIODE(net2360));
 sky130_fd_sc_hd__diode_2 ANTENNA__0665__A (.DIODE(net2361));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2361_A (.DIODE(net2362));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A (.DIODE(net2363));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2363_A (.DIODE(net2364));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__A (.DIODE(net2365));
 sky130_fd_sc_hd__diode_2 ANTENNA__0659__A (.DIODE(net2366));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2366_A (.DIODE(net2367));
 sky130_fd_sc_hd__diode_2 ANTENNA__0657__A (.DIODE(net2368));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2368_A (.DIODE(net2369));
 sky130_fd_sc_hd__diode_2 ANTENNA__0655__A (.DIODE(net2370));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2370_A (.DIODE(net2371));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A (.DIODE(net2372));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2372_A (.DIODE(net2373));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2373_A (.DIODE(net2374));
 sky130_fd_sc_hd__diode_2 ANTENNA__0651__A (.DIODE(net2375));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2375_A (.DIODE(net2376));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A (.DIODE(net2377));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__A (.DIODE(net2378));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2378_A (.DIODE(net2379));
 sky130_fd_sc_hd__diode_2 ANTENNA__0645__A (.DIODE(net2380));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2380_A (.DIODE(net2381));
 sky130_fd_sc_hd__diode_2 ANTENNA__0643__A (.DIODE(net2382));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2382_A (.DIODE(net2383));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__A (.DIODE(net2384));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2384_A (.DIODE(net2385));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__A (.DIODE(net2386));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2386_A (.DIODE(net2387));
 sky130_fd_sc_hd__diode_2 ANTENNA__0637__A (.DIODE(net2388));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2388_A (.DIODE(net2389));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__A (.DIODE(net2390));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2390_A (.DIODE(net2391));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__A (.DIODE(net2392));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2392_A (.DIODE(net2393));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2393_A (.DIODE(net2394));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2394_A (.DIODE(net2395));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__A (.DIODE(net2396));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2396_A (.DIODE(net2397));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2397_A (.DIODE(net2398));
 sky130_fd_sc_hd__diode_2 ANTENNA__0629__A (.DIODE(net2399));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2399_A (.DIODE(net2400));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2400_A (.DIODE(net2401));
 sky130_fd_sc_hd__diode_2 ANTENNA__0627__A (.DIODE(net2402));
 sky130_fd_sc_hd__diode_2 ANTENNA__0625__A (.DIODE(net2403));
 sky130_fd_sc_hd__diode_2 ANTENNA__0623__A (.DIODE(net2404));
 sky130_fd_sc_hd__diode_2 ANTENNA__0621__A (.DIODE(net2405));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2405_A (.DIODE(net2406));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__A (.DIODE(net2407));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__A (.DIODE(net2408));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2408_A (.DIODE(net2409));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__A (.DIODE(net2410));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2410_A (.DIODE(net2411));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2411_A (.DIODE(net2412));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__A (.DIODE(net2413));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2413_A (.DIODE(net2414));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__A (.DIODE(net2415));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2415_A (.DIODE(net2416));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__A (.DIODE(net2417));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2417_A (.DIODE(net2418));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2418_A (.DIODE(net2419));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A (.DIODE(net2420));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2420_A (.DIODE(net2421));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__B (.DIODE(net2422));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2422_A (.DIODE(net2423));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2423_A (.DIODE(net2424));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2424_A (.DIODE(net2425));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2425_A (.DIODE(net2426));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B (.DIODE(net2427));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2427_A (.DIODE(net2428));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2428_A (.DIODE(net2429));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2429_A (.DIODE(net2430));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__B (.DIODE(net2431));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2431_A (.DIODE(net2432));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2432_A (.DIODE(net2433));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2433_A (.DIODE(net2434));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__B (.DIODE(net2435));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2435_A (.DIODE(net2436));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2436_A (.DIODE(net2437));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2437_A (.DIODE(net2438));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__B (.DIODE(net2439));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2439_A (.DIODE(net2440));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2440_A (.DIODE(net2441));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2441_A (.DIODE(net2442));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__B (.DIODE(net2443));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2443_A (.DIODE(net2444));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2444_A (.DIODE(net2445));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2445_A (.DIODE(net2446));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__B (.DIODE(net2447));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2447_A (.DIODE(net2448));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2448_A (.DIODE(net2449));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2449_A (.DIODE(net2450));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__B (.DIODE(net2451));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2451_A (.DIODE(net2452));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2452_A (.DIODE(net2453));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2453_A (.DIODE(net2454));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__B (.DIODE(net2455));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2455_A (.DIODE(net2456));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2456_A (.DIODE(net2457));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2457_A (.DIODE(net2458));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__B (.DIODE(net2459));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2459_A (.DIODE(net2460));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2460_A (.DIODE(net2461));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A (.DIODE(net2462));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__B (.DIODE(net2463));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2463_A (.DIODE(net2464));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2464_A (.DIODE(net2465));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__B (.DIODE(net2466));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2466_A (.DIODE(net2467));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2467_A (.DIODE(net2468));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__B (.DIODE(net2469));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2469_A (.DIODE(net2470));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2470_A (.DIODE(net2471));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2471_A (.DIODE(net2472));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__B (.DIODE(net2473));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2473_A (.DIODE(net2474));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2474_A (.DIODE(net2475));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2475_A (.DIODE(net2476));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__B (.DIODE(net2477));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2477_A (.DIODE(net2478));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2478_A (.DIODE(net2479));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__B (.DIODE(net2480));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2480_A (.DIODE(net2481));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__B (.DIODE(net2482));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2482_A (.DIODE(net2483));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2483_A (.DIODE(net2484));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__B (.DIODE(net2485));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2485_A (.DIODE(net2486));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2486_A (.DIODE(net2487));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2487_A (.DIODE(net2488));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__B (.DIODE(net2489));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2489_A (.DIODE(net2490));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2490_A (.DIODE(net2491));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__B (.DIODE(net2492));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2492_A (.DIODE(net2493));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2493_A (.DIODE(net2494));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__B (.DIODE(net2495));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2495_A (.DIODE(net2496));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2496_A (.DIODE(net2497));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__B (.DIODE(net2498));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2498_A (.DIODE(net2499));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2499_A (.DIODE(net2500));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__B (.DIODE(net2501));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2501_A (.DIODE(net2502));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2502_A (.DIODE(net2503));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__B (.DIODE(net2504));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2504_A (.DIODE(net2505));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__B (.DIODE(net2506));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2506_A (.DIODE(net2507));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2507_A (.DIODE(net2508));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__B (.DIODE(net2509));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2509_A (.DIODE(net2510));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2510_A (.DIODE(net2511));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__B (.DIODE(net2512));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2512_A (.DIODE(net2513));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2513_A (.DIODE(net2514));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__B (.DIODE(net2515));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2515_A (.DIODE(net2516));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2516_A (.DIODE(net2517));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__B (.DIODE(net2518));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2518_A (.DIODE(net2519));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2519_A (.DIODE(net2520));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__B (.DIODE(net2521));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2521_A (.DIODE(net2522));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2522_A (.DIODE(net2523));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(net2524));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2524_A (.DIODE(net2525));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2525_A (.DIODE(net2526));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2526_A (.DIODE(net2527));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2527_A (.DIODE(net2528));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__B (.DIODE(net2529));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2529_A (.DIODE(net2530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__B (.DIODE(net2531));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2531_A (.DIODE(net2532));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2532_A (.DIODE(net2533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__B (.DIODE(net2534));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2534_A (.DIODE(net2535));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2535_A (.DIODE(net2536));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__B (.DIODE(net2537));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2537_A (.DIODE(net2538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1461__B (.DIODE(net2539));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2539_A (.DIODE(net2540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__B (.DIODE(net2541));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__B (.DIODE(net2542));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__B (.DIODE(net2543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__B (.DIODE(net2544));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2544_A (.DIODE(net2545));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2545_A (.DIODE(net2546));
 sky130_fd_sc_hd__diode_2 ANTENNA__0927__A (.DIODE(net2547));
 sky130_fd_sc_hd__diode_2 ANTENNA__1449__B (.DIODE(net2548));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2548_A (.DIODE(net2549));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2549_A (.DIODE(net2550));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__B (.DIODE(net2551));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2551_A (.DIODE(net2552));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2552_A (.DIODE(net2553));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2553_A (.DIODE(net2554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1445__B (.DIODE(net2555));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2555_A (.DIODE(net2556));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2556_A (.DIODE(net2557));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__B (.DIODE(net2558));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2558_A (.DIODE(net2559));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2559_A (.DIODE(net2560));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__B (.DIODE(net2561));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2561_A (.DIODE(net2562));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2562_A (.DIODE(net2563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1439__B (.DIODE(net2564));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2564_A (.DIODE(net2565));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2565_A (.DIODE(net2566));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2566_A (.DIODE(net2567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__B (.DIODE(net2568));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2568_A (.DIODE(net2569));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__B (.DIODE(net2570));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2570_A (.DIODE(net2571));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2571_A (.DIODE(net2572));
 sky130_fd_sc_hd__diode_2 ANTENNA__1433__B (.DIODE(net2573));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2573_A (.DIODE(net2574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__B (.DIODE(net2575));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2575_A (.DIODE(net2576));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2576_A (.DIODE(net2577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__B (.DIODE(net2578));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2578_A (.DIODE(net2579));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2579_A (.DIODE(net2580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__B (.DIODE(net2581));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2581_A (.DIODE(net2582));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2582_A (.DIODE(net2583));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__B (.DIODE(net2584));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2584_A (.DIODE(net2585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__B (.DIODE(net2586));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2586_A (.DIODE(net2587));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__B (.DIODE(net2588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__B (.DIODE(net2589));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2589_A (.DIODE(net2590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__B (.DIODE(net2591));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2591_A (.DIODE(net2592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__B (.DIODE(net2593));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__B (.DIODE(net2594));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__B (.DIODE(net2595));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2595_A (.DIODE(net2596));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__A (.DIODE(net2597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__B (.DIODE(net2598));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__B (.DIODE(net2599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__B (.DIODE(net2600));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__B (.DIODE(net2601));
 sky130_fd_sc_hd__diode_2 ANTENNA__1385__B (.DIODE(net2602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__B (.DIODE(net2603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1379__B (.DIODE(net2604));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__B (.DIODE(net2605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__B (.DIODE(net2606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__B (.DIODE(net2607));
 sky130_fd_sc_hd__diode_2 ANTENNA__1357__B (.DIODE(net2608));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__B (.DIODE(net2609));
 sky130_fd_sc_hd__diode_2 ANTENNA__1343__B (.DIODE(net2610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__B (.DIODE(net2611));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__B (.DIODE(net2612));
 sky130_fd_sc_hd__diode_2 ANTENNA__1337__B (.DIODE(net2613));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2613_A (.DIODE(net2614));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__B (.DIODE(net2615));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__B (.DIODE(net2616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__B (.DIODE(net2617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__B (.DIODE(net2618));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2618_A (.DIODE(net2619));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__B (.DIODE(net2620));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2620_A (.DIODE(net2621));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B (.DIODE(net2622));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__B (.DIODE(net2623));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2623_A (.DIODE(net2624));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2624_A (.DIODE(net2625));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__B (.DIODE(net2626));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__B (.DIODE(net2627));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__B (.DIODE(net2628));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2628_A (.DIODE(net2629));
 sky130_fd_sc_hd__diode_2 ANTENNA__1313__B (.DIODE(net2630));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2630_A (.DIODE(net2631));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__B (.DIODE(net2632));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2632_A (.DIODE(net2633));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2633_A (.DIODE(net2634));
 sky130_fd_sc_hd__diode_2 ANTENNA__0913__A (.DIODE(net2635));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__B (.DIODE(net2636));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2636_A (.DIODE(net2637));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__B (.DIODE(net2638));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2638_A (.DIODE(net2639));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__B (.DIODE(net2640));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2640_A (.DIODE(net2641));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__B (.DIODE(net2642));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2642_A (.DIODE(net2643));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2643_A (.DIODE(net2644));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__B (.DIODE(net2645));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2645_A (.DIODE(net2646));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2646_A (.DIODE(net2647));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__B (.DIODE(net2648));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__B (.DIODE(net2649));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2649_A (.DIODE(net2650));
 sky130_fd_sc_hd__diode_2 ANTENNA__1295__B (.DIODE(net2651));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2651_A (.DIODE(net2652));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2652_A (.DIODE(net2653));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__B (.DIODE(net2654));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2654_A (.DIODE(net2655));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2655_A (.DIODE(net2656));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__B (.DIODE(net2657));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2657_A (.DIODE(net2658));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__B (.DIODE(net2659));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2659_A (.DIODE(net2660));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__B (.DIODE(net2661));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2661_A (.DIODE(net2662));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2662_A (.DIODE(net2663));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__B (.DIODE(net2664));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2664_A (.DIODE(net2665));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2665_A (.DIODE(net2666));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__B (.DIODE(net2667));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2667_A (.DIODE(net2668));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__B (.DIODE(net2669));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2669_A (.DIODE(net2670));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2670_A (.DIODE(net2671));
 sky130_fd_sc_hd__diode_2 ANTENNA__1279__B (.DIODE(net2672));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2672_A (.DIODE(net2673));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2673_A (.DIODE(net2674));
 sky130_fd_sc_hd__diode_2 ANTENNA__1277__B (.DIODE(net2675));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2675_A (.DIODE(net2676));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2676_A (.DIODE(net2677));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__B (.DIODE(net2678));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2678_A (.DIODE(net2679));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__B (.DIODE(net2680));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2680_A (.DIODE(net2681));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2681_A (.DIODE(net2682));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__B (.DIODE(net2683));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2683_A (.DIODE(net2684));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2684_A (.DIODE(net2685));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2685_A (.DIODE(net2686));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__B (.DIODE(net2687));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2687_A (.DIODE(net2688));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2688_A (.DIODE(net2689));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2689_A (.DIODE(net2690));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__B (.DIODE(net2691));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2691_A (.DIODE(net2692));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2692_A (.DIODE(net2693));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2693_A (.DIODE(net2694));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__B (.DIODE(net2695));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2695_A (.DIODE(net2696));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2696_A (.DIODE(net2697));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__B (.DIODE(net2698));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2698_A (.DIODE(net2699));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2699_A (.DIODE(net2700));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__B (.DIODE(net2701));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2701_A (.DIODE(net2702));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2702_A (.DIODE(net2703));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2703_A (.DIODE(net2704));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__B (.DIODE(net2705));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2705_A (.DIODE(net2706));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2706_A (.DIODE(net2707));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__B (.DIODE(net2708));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2708_A (.DIODE(net2709));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2709_A (.DIODE(net2710));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__B (.DIODE(net2711));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2711_A (.DIODE(net2712));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2712_A (.DIODE(net2713));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__B (.DIODE(net2714));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2714_A (.DIODE(net2715));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__B (.DIODE(net2716));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2716_A (.DIODE(net2717));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2717_A (.DIODE(net2718));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__B (.DIODE(net2719));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2719_A (.DIODE(net2720));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2720_A (.DIODE(net2721));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__B (.DIODE(net2722));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2722_A (.DIODE(net2723));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2723_A (.DIODE(net2724));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__B (.DIODE(net2725));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2725_A (.DIODE(net2726));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__B (.DIODE(net2727));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2727_A (.DIODE(net2728));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__B (.DIODE(net2729));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2729_A (.DIODE(net2730));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2730_A (.DIODE(net2731));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__B (.DIODE(net2732));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2732_A (.DIODE(net2733));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__B (.DIODE(net2734));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2734_A (.DIODE(net2735));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__B (.DIODE(net2736));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2736_A (.DIODE(net2737));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2737_A (.DIODE(net2738));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__B (.DIODE(net2739));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2739_A (.DIODE(net2740));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__B (.DIODE(net2741));
 sky130_fd_sc_hd__diode_2 ANTENNA__0905__A (.DIODE(net2742));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__B (.DIODE(net2743));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2743_A (.DIODE(net2744));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__B (.DIODE(net2745));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__B (.DIODE(net2746));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2746_A (.DIODE(net2747));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__B (.DIODE(net2748));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2748_A (.DIODE(net2749));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__B (.DIODE(net2750));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__B (.DIODE(net2751));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2751_A (.DIODE(net2752));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__B (.DIODE(net2753));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__B (.DIODE(net2754));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__B (.DIODE(net2755));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__B (.DIODE(net2756));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__B (.DIODE(net2757));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2757_A (.DIODE(net2758));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__B (.DIODE(net2759));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__B (.DIODE(net2760));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__B (.DIODE(net2761));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__B (.DIODE(net2762));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__B (.DIODE(net2763));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__B (.DIODE(net2764));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2764_A (.DIODE(net2765));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2765_A (.DIODE(net2766));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__B (.DIODE(net2767));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2767_A (.DIODE(net2768));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2768_A (.DIODE(net2769));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2769_A (.DIODE(net2770));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2770_A (.DIODE(net2771));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__B (.DIODE(net2772));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2772_A (.DIODE(net2773));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2773_A (.DIODE(net2774));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2774_A (.DIODE(net2775));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__B (.DIODE(net2776));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2776_A (.DIODE(net2777));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2777_A (.DIODE(net2778));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2778_A (.DIODE(net2779));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B (.DIODE(net2780));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2780_A (.DIODE(net2781));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2781_A (.DIODE(net2782));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__B (.DIODE(net2783));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2783_A (.DIODE(net2784));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2784_A (.DIODE(net2785));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2785_A (.DIODE(net2786));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__B (.DIODE(net2787));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2787_A (.DIODE(net2788));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2788_A (.DIODE(net2789));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2789_A (.DIODE(net2790));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__B (.DIODE(net2791));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2791_A (.DIODE(net2792));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2792_A (.DIODE(net2793));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2793_A (.DIODE(net2794));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__B (.DIODE(net2795));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2795_A (.DIODE(net2796));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2796_A (.DIODE(net2797));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2797_A (.DIODE(net2798));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__B (.DIODE(net2799));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2799_A (.DIODE(net2800));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__B (.DIODE(net2801));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2801_A (.DIODE(net2802));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2802_A (.DIODE(net2803));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__B (.DIODE(net2804));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2804_A (.DIODE(net2805));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2805_A (.DIODE(net2806));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__B (.DIODE(net2807));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2807_A (.DIODE(net2808));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2808_A (.DIODE(net2809));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__A (.DIODE(net2810));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__B (.DIODE(net2811));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2811_A (.DIODE(net2812));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__B (.DIODE(net2813));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2813_A (.DIODE(net2814));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2814_A (.DIODE(net2815));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__B (.DIODE(net2816));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2816_A (.DIODE(net2817));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__B (.DIODE(net2818));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2818_A (.DIODE(net2819));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__B (.DIODE(net2820));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2820_A (.DIODE(net2821));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__B (.DIODE(net2822));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2822_A (.DIODE(net2823));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__B (.DIODE(net2824));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__B (.DIODE(net2825));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2825_A (.DIODE(net2826));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__B (.DIODE(net2827));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__B (.DIODE(net2828));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A (.DIODE(net2829));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__B (.DIODE(net2830));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__B (.DIODE(net2831));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__B (.DIODE(net2832));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__B (.DIODE(net2833));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__B (.DIODE(net2834));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__B (.DIODE(net2835));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__B (.DIODE(net2836));
 sky130_fd_sc_hd__diode_2 ANTENNA__0891__A (.DIODE(net2837));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__B (.DIODE(net2838));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__B (.DIODE(net2839));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__B (.DIODE(net2840));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__B (.DIODE(net2841));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__B (.DIODE(net2842));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2842_A (.DIODE(net2843));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__B (.DIODE(net2844));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__B (.DIODE(net2845));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2845_A (.DIODE(net2846));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__B (.DIODE(net2847));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B (.DIODE(net2848));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2848_A (.DIODE(net2849));
 sky130_fd_sc_hd__diode_2 ANTENNA_output953_A (.DIODE(net2850));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2850_A (.DIODE(net2851));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2851_A (.DIODE(net2852));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2852_A (.DIODE(net2853));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2853_A (.DIODE(net2854));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2854_A (.DIODE(net2855));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3081 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3666 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1191 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1419 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1501 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1510 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1528 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1536 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1547 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1598 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1613 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1620 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1637 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1669 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1686 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1692 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1715 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1723 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1743 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1749 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1763 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1791 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1812 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1836 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1846 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1849 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1859 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1871 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1879 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1885 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1893 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1901 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1911 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1923 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1931 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1939 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1947 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1959 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1970 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1977 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1997 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2003 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2013 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2017 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2023 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2031 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2039 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2051 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2079 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2085 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2099 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2106 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2112 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2123 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2127 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2135 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2143 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2173 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2182 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2185 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2197 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2206 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2214 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2219 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2247 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2267 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2274 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2291 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2308 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2316 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2333 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2347 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2368 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2382 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2389 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2395 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2416 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2424 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2431 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2438 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2451 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2465 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2470 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2476 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2481 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2501 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2515 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2527 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2535 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2542 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2550 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2562 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2596 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2602 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2607 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2614 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2622 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2627 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2649 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2669 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2683 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2689 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2703 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2709 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2723 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2731 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2738 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2751 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2765 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2781 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2789 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2801 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2817 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2837 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2845 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2852 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2873 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2895 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2927 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2935 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2943 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_2957 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2965 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_2969 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2981 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3005 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3019 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3023 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3025 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3037 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3061 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3069 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3076 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3087 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3094 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3101 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3111 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3117 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3132 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3144 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3153 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3173 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3181 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3198 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3213 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3227 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3235 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3243 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3247 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3255 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3263 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3269 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3274 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3280 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3290 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3302 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3305 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3316 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3324 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3334 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3342 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3348 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3359 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3395 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3408 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3414 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3428 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3432 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3442 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3450 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3458 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3466 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3491 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3511 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3519 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3534 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3538 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3543 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3563 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3590 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3597 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3617 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3625 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3638 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3651 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3671 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3684 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3692 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3705 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3725 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3732 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3738 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3748 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3759 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3779 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3793 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3806 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3813 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3833 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3846 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3859 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3863 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3887 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3900 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3907 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3914 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3945 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_3957 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_3968 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4031 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_4033 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4047 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4071 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_4083 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1059 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1184 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1280 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1302 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1331 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1397 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1447 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1455 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1508 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1520 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1528 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1546 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1565 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1586 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1590 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1594 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1617 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1631 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1643 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1649 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1664 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1672 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1675 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1683 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1695 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1714 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1725 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1732 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1743 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1750 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1758 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1762 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1774 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1780 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1783 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1792 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1804 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1810 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1845 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1848 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1852 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1855 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1863 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1867 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1882 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1894 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1901 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1907 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1911 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1915 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1922 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1928 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1939 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1951 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1960 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1968 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1972 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1978 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1995 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2002 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2010 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2015 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2021 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2027 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2045 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2050 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2056 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2059 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2065 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2077 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2087 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2101 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2105 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2113 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2117 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2121 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2147 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2153 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2171 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2183 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2188 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2194 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2200 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2206 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2213 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2218 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2225 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2237 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2250 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2256 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2260 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2273 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2287 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2293 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2301 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2306 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2310 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2320 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2331 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2337 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2345 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2349 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2356 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2362 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2368 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2374 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2386 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2394 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2398 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2405 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2423 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2430 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2437 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2441 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2452 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2458 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2464 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2470 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2476 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2501 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2508 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2514 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2520 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2524 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2531 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2539 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2546 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2554 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2560 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2568 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2572 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2578 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2596 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2602 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2605 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2610 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2616 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2620 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2626 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2635 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2640 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2651 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2657 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2665 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2671 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2679 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2685 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2693 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2708 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2714 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2721 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2727 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2733 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2740 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2747 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2753 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2762 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2768 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2773 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2788 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2794 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2800 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2806 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2819 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2834 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2838 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2843 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2850 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2854 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2858 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2865 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2872 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2879 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2890 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_2896 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2904 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2908 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2915 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2925 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2941 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2963 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2973 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_2981 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_2997 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3003 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3013 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3021 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3028 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3032 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3043 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3050 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3065 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3079 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3084 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3088 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3100 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3106 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3115 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3122 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3130 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3144 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3154 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3177 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3201 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3209 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3221 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3229 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3238 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3245 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3252 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3260 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3268 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3274 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3284 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3294 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3301 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3308 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3314 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3318 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3322 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3326 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3330 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3338 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3342 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3346 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3354 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3362 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3382 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3399 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3405 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3415 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3425 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3433 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3440 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3450 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3454 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3458 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3465 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3478 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3485 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3492 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3498 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3501 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3527 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3532 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3546 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3557 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3568 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3582 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3589 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3600 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3610 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3613 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3621 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3627 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3632 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3638 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3643 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3674 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3681 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3694 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3702 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3709 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3716 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3722 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3725 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3730 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3737 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3744 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3750 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3756 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3766 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3777 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3781 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3797 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3815 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_3833 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3843 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3850 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3856 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3861 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3874 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3887 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3891 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3899 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3906 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3912 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3918 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3930 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_3938 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3961 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3973 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_3984 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3990 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1327 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1354 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1372 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1382 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1407 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1474 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1484 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1506 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1523 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1529 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1532 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1543 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1557 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1579 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1586 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1592 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1598 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1610 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1614 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1652 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1656 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1711 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1722 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1728 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1734 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1741 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1744 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1752 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1758 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1762 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1768 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1771 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1805 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1815 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1853 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1865 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1876 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1888 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1892 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1895 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1905 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1909 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1927 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1957 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1969 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1972 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1976 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1979 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1988 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1996 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2005 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2049 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2054 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2060 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2079 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2123 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2143 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2151 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2159 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2164 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2170 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2191 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2203 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2211 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2215 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2227 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2247 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2253 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2259 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2291 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2301 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2309 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2315 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2323 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2357 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2364 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2370 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2376 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2388 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2392 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2395 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2413 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2419 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2425 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2431 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2443 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2446 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_2454 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2477 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2483 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2495 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2507 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2515 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2521 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2525 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2538 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2544 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2550 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2556 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2560 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2581 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2607 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2617 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2626 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2637 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2641 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2679 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2686 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2697 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2703 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2710 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2716 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2726 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2736 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2742 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2749 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2753 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2756 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2762 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2768 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_2774 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2782 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2786 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2792 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2805 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2811 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2817 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2823 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2847 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_2853 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2861 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2867 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2873 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2879 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2891 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2903 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2925 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2931 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2937 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2943 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2952 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2960 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2966 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2975 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2979 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2984 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_2992 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3000 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3006 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3014 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3018 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3034 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3040 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3046 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3052 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3058 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3062 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3067 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3074 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3085 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3100 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3117 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3123 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3135 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3137 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3141 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3149 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3153 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3161 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3167 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3179 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3187 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3191 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3208 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3216 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3224 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3232 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3238 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3246 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3255 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3262 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3271 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3279 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3287 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3295 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3316 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3322 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3328 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3334 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3338 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3342 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3347 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3367 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3375 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3383 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3387 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3395 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3401 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3405 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3411 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3415 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3423 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3428 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3436 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3441 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3447 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3453 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3457 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3464 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3470 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3477 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3483 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3495 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3507 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3513 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3519 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3525 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3547 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3555 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3562 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3568 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3580 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3591 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3597 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3612 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3616 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3624 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3631 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3638 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3650 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3658 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3664 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3672 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3679 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3687 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3693 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3702 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3708 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3714 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3720 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3724 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3727 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3736 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3742 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3748 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3757 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3763 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3771 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3784 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3792 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3798 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3803 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3807 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3820 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3827 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3834 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3838 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3843 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3854 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3861 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3865 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3871 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3877 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3884 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3891 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3901 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3906 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3918 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3975 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3977 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_3982 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3988 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4012 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_4024 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1519 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1531 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1547 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1554 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1564 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1576 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1580 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1583 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1609 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1731 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1743 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1753 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1759 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1939 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1951 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1963 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1998 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2004 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2016 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2028 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2040 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2123 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2135 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2164 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2176 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2184 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2225 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2235 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2243 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2255 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2279 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2299 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2365 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2393 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2399 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2402 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2408 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2411 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2461 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2464 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2472 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2478 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2566 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2578 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2582 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2586 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2592 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2596 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2601 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2609 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2613 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2616 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2620 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2623 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2646 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2658 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2721 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2727 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2733 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2744 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2750 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2756 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2760 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2778 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2787 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2795 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2803 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2809 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2815 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2841 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2853 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2859 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2865 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2871 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2889 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2895 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2908 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2914 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2920 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2926 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2932 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_2937 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2947 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2951 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2955 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2959 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_2964 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2972 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2976 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2984 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2992 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3005 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3013 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3019 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3031 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3037 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3043 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3063 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3069 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3076 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3090 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3094 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3099 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3105 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3113 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3119 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3127 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3132 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3138 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3144 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3150 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3156 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3169 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3175 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3181 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3187 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3206 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3214 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3221 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3226 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3234 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3241 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3249 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3255 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3267 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3274 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3282 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3288 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3294 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3307 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3317 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3323 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3329 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3333 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3341 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3350 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3356 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3360 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3371 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3387 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3395 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3401 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3407 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3413 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3419 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3425 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3429 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3432 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3440 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3449 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3455 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3461 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3467 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3470 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3476 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3482 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3488 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3494 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3511 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3519 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3529 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3535 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3540 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3555 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3557 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3562 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3571 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3578 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3590 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3596 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3602 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3608 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3617 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3623 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3632 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3638 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3642 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3646 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3652 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3667 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3675 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3682 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3688 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3694 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3700 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3706 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3718 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3725 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3729 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3739 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3758 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3770 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3778 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3787 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3793 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3801 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3807 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3819 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3824 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3830 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3837 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3841 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3850 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3856 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3862 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3868 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3874 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3880 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3886 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3897 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3909 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3913 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3922 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3934 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3961 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3973 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3980 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3986 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3998 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1302 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1567 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1575 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1587 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1594 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1604 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1612 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1630 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1636 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1660 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1820 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1832 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1844 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1873 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1881 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1884 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2097 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2107 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2119 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2141 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2144 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2190 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2194 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2229 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2312 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2320 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2328 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2334 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2346 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2421 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2424 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2432 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2444 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2456 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2499 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2561 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2597 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2602 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2610 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2618 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2626 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2644 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2652 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2670 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2676 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2731 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2742 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2754 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2762 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2770 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2778 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2792 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2809 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2816 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2822 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2828 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2834 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2840 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2846 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2861 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2870 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2880 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_2888 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2896 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2901 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2905 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2910 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2921 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2929 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2935 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2953 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2959 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_2965 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2973 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2981 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2993 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3003 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3007 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3012 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3018 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3029 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3033 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3038 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3048 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3054 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3060 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3072 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3078 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3085 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3091 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3097 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3103 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3115 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3127 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3143 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3149 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3155 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3161 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3179 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3191 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3197 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3203 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3209 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3215 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3227 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3233 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3239 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3245 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3253 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3259 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3265 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3271 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3283 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3295 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3305 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3311 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3317 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3324 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3330 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3336 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3344 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3349 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3359 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3365 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3372 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3380 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3386 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3400 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3406 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3412 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3421 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3427 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3439 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3451 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3468 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3478 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3484 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3492 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3498 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3508 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3514 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3520 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3533 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3545 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3551 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3563 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3569 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3575 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3591 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3599 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3605 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3611 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3623 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3629 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3635 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3639 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3645 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3651 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3655 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3658 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3664 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3670 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3674 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3677 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3683 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3765 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3777 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3785 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3789 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3797 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3809 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3821 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3829 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3835 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3841 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3847 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3856 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3862 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3881 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3893 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3901 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3906 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_3912 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4087 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_4094 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1512 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1797 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1883 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1888 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1900 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1912 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1924 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2027 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2033 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2036 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2093 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2097 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2110 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2122 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2134 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2140 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2148 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2154 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2162 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2174 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2192 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2198 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2295 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2303 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2312 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2320 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2348 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2360 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2372 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2388 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2394 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2406 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2420 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2428 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2461 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2479 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2611 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2614 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2618 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2621 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2627 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2632 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2638 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2648 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2675 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2687 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2691 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2699 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2711 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2717 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2731 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2743 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2753 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2763 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2769 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2787 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2795 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2810 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2820 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2839 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2851 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2861 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2871 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2879 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2883 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2907 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2915 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2925 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2937 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2953 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2959 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2965 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2977 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2985 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2994 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3005 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3011 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3015 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3031 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3035 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3042 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3050 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3053 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3062 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3068 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3074 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3080 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3086 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3092 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3096 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3103 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3107 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3119 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3125 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3131 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3143 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3155 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3171 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3177 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3187 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3195 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3200 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3208 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3214 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3227 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3233 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3239 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3245 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3251 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3257 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3263 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3275 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3281 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3293 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3296 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3304 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3310 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3316 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3322 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3328 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3339 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3347 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3353 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3359 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3367 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3373 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3379 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3385 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3399 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3405 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3417 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3423 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3426 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3439 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3443 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3455 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3469 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3475 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3479 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3484 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3490 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3496 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3501 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3507 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3515 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3519 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3523 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3529 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3533 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3536 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3542 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3552 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3561 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3567 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3575 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3583 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3587 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3593 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3599 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3627 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3639 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3643 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3651 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3656 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3660 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3663 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3681 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3693 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3700 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3706 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3718 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3835 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3842 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3848 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3858 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3876 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1789 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1799 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1804 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1816 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1957 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1965 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1977 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1983 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2013 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2021 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2024 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2032 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2040 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2053 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2057 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2060 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2066 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2085 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2091 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2097 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2101 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2107 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2116 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2122 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2155 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2167 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2173 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2195 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2201 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2207 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2224 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2236 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2245 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2277 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2280 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2288 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2337 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2369 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2423 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2431 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2477 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2486 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2497 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2509 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2533 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2561 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2589 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2597 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2602 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2611 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2619 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2625 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2641 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2647 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2655 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2658 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2671 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2683 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2695 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2701 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2707 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2713 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2725 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2731 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2735 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2742 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2760 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2789 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2796 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2801 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2817 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2835 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2849 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2854 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2868 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2882 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2894 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2900 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2910 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2921 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2931 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2937 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2949 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2957 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2965 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2973 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2986 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2994 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3001 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3014 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3022 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3037 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3050 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3061 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3067 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3079 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3085 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3091 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3097 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3107 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3119 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3134 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3141 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3147 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3153 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3158 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3177 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3191 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3197 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3203 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3209 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3215 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3219 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3231 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3237 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3243 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3247 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3253 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3266 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3293 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3299 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3309 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3315 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3323 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3329 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3341 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3349 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3365 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3371 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3377 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3383 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3387 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3395 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3398 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3414 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3441 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3445 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3452 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3460 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3473 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3485 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3491 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3497 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3501 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3508 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3516 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3533 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3545 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3550 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3565 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3573 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3579 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3597 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3613 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3625 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3629 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3635 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3681 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3697 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3709 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3717 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3722 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3732 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_3744 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3765 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3777 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3786 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3792 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3849 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3877 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3908 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3914 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3921 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3935 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4005 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4010 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4016 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1459 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1479 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1491 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1516 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1528 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1535 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1559 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1571 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1582 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1591 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1629 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1641 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1647 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1671 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1683 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1703 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1727 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1744 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1756 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1759 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1763 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1769 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1772 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1778 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1800 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1808 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1815 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1841 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1853 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1859 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1867 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1871 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1881 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1904 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1916 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1920 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1936 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1944 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1947 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1953 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1965 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1971 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1983 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2005 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2013 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2023 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2031 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2037 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2039 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2047 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2053 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2060 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2067 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2079 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2088 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2095 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2105 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2110 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2118 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2126 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2132 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2138 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2155 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2161 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2175 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2189 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2194 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2202 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2207 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2211 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2223 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2229 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2235 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2239 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2244 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2250 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2256 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2263 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2271 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2317 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2319 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2335 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2365 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2399 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2411 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2419 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2431 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2447 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2459 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2471 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2483 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2487 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2495 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2513 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2525 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2539 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2543 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2559 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2583 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2599 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2611 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2617 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2625 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2641 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2652 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2655 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2659 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2665 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2675 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_2683 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2691 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2694 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2700 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2704 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3086 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3092 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3096 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3103 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3117 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3123 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3133 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3150 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3156 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3162 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3164 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3173 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3179 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3185 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3191 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3209 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3215 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3226 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3232 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3238 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3250 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3262 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3300 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3318 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3324 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3327 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3332 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3337 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3343 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3349 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3352 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3358 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3364 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3370 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3376 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3456 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3468 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3472 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3478 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3486 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3512 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3536 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3556 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_3568 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3576 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3594 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3606 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3624 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3704 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3716 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3760 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3778 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3785 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3797 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3821 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3928 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3940 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3996 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4002 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_4004 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_4010 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4019 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4043 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4057 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4066 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4078 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_4090 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4098 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1431 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1463 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1475 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1478 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1488 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1494 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1543 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1552 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1560 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1563 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1568 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1576 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1584 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1596 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1602 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1610 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1616 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1619 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1631 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1655 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1667 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1675 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1699 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1711 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1719 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1724 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1731 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1735 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1741 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1744 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1750 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1758 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1770 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1778 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1784 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1787 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1791 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1799 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1820 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1828 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1836 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1843 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1853 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1861 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1874 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1882 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1890 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1895 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1899 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1903 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1909 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1912 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1920 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1930 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1938 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1944 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1952 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1955 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1965 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1973 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1985 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1990 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1996 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2008 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2011 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2021 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2031 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2039 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2043 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2048 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2056 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2064 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2067 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2081 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2089 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2097 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2105 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2123 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2129 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2135 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2149 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2166 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2179 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2193 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2201 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2209 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2221 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2226 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2232 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2235 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2243 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2251 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2263 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2276 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2282 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2291 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2327 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2345 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2347 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2362 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2368 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2380 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2392 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2403 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2427 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2445 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2459 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2471 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2491 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2503 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2509 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2515 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2527 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2539 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2547 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2552 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2560 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2568 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2571 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2595 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2607 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2615 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_2623 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2627 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2631 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2637 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2643 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2649 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2662 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2674 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2680 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2683 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2691 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2694 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2700 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2704 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3090 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3096 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3102 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3114 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3120 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3126 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3132 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3142 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3148 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3154 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3160 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3166 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3172 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3178 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3190 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3192 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3196 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3208 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3214 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3222 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3228 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3234 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3246 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3260 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3284 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3296 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3302 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3316 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3328 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3340 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3355 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3360 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3364 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3372 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3380 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3386 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3398 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3410 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3414 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3416 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3428 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3436 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3440 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3453 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3461 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3540 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3552 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3562 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3575 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3596 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3603 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3633 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3644 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3656 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3692 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3696 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3702 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3711 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3735 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3747 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3752 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3764 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3772 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3778 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3784 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3790 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3796 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3844 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3856 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3862 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3876 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3900 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3912 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3920 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_3925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3931 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3943 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3952 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3964 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3988 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4012 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_4024 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4029 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4068 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4080 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4086 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_4088 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1179 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1291 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1447 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1459 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1467 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1479 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1483 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1502 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1506 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1511 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1520 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1535 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1547 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1572 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1580 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1591 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1603 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1608 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1615 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1619 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1624 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1628 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1647 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1651 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1659 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1663 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1674 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1682 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1696 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1714 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1722 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1730 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1738 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1748 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1756 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1759 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1769 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1779 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1787 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1795 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1799 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1804 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1812 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1815 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1827 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1831 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1836 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1844 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1852 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1860 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1868 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1871 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1890 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1894 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1908 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1916 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1924 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1927 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1932 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1940 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1944 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1949 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1958 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1964 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1972 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1980 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1983 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1995 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2003 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2011 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2019 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2032 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2039 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2049 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2065 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2086 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2092 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2095 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2117 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2125 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2133 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2147 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2159 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2171 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2181 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2189 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2195 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2204 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2207 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2220 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2228 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2234 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2240 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2252 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2260 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2263 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2267 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2280 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2286 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2298 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2302 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2311 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2319 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2355 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2367 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2387 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2407 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2419 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2427 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2431 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2450 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2462 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2474 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2487 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2491 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2494 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2502 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2514 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2526 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2538 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2543 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2555 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2567 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2572 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2578 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2590 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2599 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2603 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2611 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2619 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2625 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2631 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2643 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2655 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2675 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2683 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2691 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_2694 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3090 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3098 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3104 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3112 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3118 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3124 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3130 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3142 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3154 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3160 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3174 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3180 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3186 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3192 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3198 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3204 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3210 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3218 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3220 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3226 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3232 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3239 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3245 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3253 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3257 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3263 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3312 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3330 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3344 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3356 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3368 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3376 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3381 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3424 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3436 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3456 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3480 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3492 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3498 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3506 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3518 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3530 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3542 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3554 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3556 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3562 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3570 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3575 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3605 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3624 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3636 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3642 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3692 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3698 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3706 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3712 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3748 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3760 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3770 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3780 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3792 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3795 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3802 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3817 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3823 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3892 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3904 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3908 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3913 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3925 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3937 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3945 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3959 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3971 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3983 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3995 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4016 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4040 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4052 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4072 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4084 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4096 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4102 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1211 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1295 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1323 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1395 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1407 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1419 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1476 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1488 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1507 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1518 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1524 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1532 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1535 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1542 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1551 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1563 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1574 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1578 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1588 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1591 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1608 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1616 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1630 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1643 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1647 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1651 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1667 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1672 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1675 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1682 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1690 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1698 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1703 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1711 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1724 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1731 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1742 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1756 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1759 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1770 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1780 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1787 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1791 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1799 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1815 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1819 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1823 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1839 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1843 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1847 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1855 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1868 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1871 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1881 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1896 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1899 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1910 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1916 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1924 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1927 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1931 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1936 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1944 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1952 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1955 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1960 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1973 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1977 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1980 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1983 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1990 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1998 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2008 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2011 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2022 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2028 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2036 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2039 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2050 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2056 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2064 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2067 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2079 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2092 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2095 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2106 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2114 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2120 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2123 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2137 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2145 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2149 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2174 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2179 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2190 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2198 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2204 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2207 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2218 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2228 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2235 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2241 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2247 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2259 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2263 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2267 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2284 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2291 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2296 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2308 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2316 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2319 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2323 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2329 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2344 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2347 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2363 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2371 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2387 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2399 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2403 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2411 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2423 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2429 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2431 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2442 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2448 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2456 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2459 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2467 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2478 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2484 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2499 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2515 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2534 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2540 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2543 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2553 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2565 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2583 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_2595 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2599 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2603 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2615 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2619 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2622 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2627 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2635 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2638 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2655 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2659 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2662 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2668 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2674 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2680 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2683 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2687 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3090 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3098 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3104 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3120 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3126 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3136 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3152 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3158 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3174 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3180 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3188 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3192 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3205 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3217 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3230 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3240 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3246 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3248 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3252 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3255 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3266 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3290 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3302 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3304 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3316 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3324 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3330 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3336 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3348 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3356 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3372 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3384 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3400 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3428 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3456 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3468 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3472 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3484 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3496 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3500 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3506 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3518 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3528 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3540 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3552 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3556 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3568 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3576 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3592 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3604 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3610 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3624 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3652 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3664 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3674 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3690 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3694 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3696 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3704 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3708 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3714 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3736 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3792 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3820 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3832 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3841 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3853 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3861 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3864 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3872 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3879 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3904 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3916 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3920 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3931 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3943 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3960 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3972 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3976 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3982 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3985 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3994 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4016 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4032 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_4044 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4052 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4057 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4072 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1335 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1403 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1423 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1437 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2256 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2262 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2268 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2285 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2291 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2318 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2322 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2327 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2335 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2371 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2374 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2383 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2399 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2423 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2435 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2499 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2511 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2523 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2529 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2539 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2545 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2551 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2559 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2565 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2578 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2590 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2593 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2608 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2611 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2615 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2628 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2640 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2652 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2658 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2664 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2671 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2674 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2693 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3090 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3100 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3106 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3116 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3122 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3128 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3134 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3152 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3158 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3174 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3180 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3186 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3198 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3210 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3218 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3230 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3262 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3274 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3276 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3284 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3288 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3299 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3311 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3315 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3318 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3328 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3332 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3339 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3349 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3364 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3372 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3384 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3388 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3400 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3408 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3413 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3429 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3435 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3456 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3468 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3480 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3490 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3497 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3500 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3508 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3514 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3520 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3538 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3550 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3554 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3556 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3564 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3571 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3577 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3601 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3624 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3680 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3696 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3708 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3711 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3717 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3724 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3732 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3738 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3750 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3762 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3834 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3836 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3847 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3859 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3879 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3928 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3940 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3946 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3948 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3953 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3962 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3974 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3982 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3990 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4016 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4028 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4036 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4048 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_4056 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4069 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4081 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_4093 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1299 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1323 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1351 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1375 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1393 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1421 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2255 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2261 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2278 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2284 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2290 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2300 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2312 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2318 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2324 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2330 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2336 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2342 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2354 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2363 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2399 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2411 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2419 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2449 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2461 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2469 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2501 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2513 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2516 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2522 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2541 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2547 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2553 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2559 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2565 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2571 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2577 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2581 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2591 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2597 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2618 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2643 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2649 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2655 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2661 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2665 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2670 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2676 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2692 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3090 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3100 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3108 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3116 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3122 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3127 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3158 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3170 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3176 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3180 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3188 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3196 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3208 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3220 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3223 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3229 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3232 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3238 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3242 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3245 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3248 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3260 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3278 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3292 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3298 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3301 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3304 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3310 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3318 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3329 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3366 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3378 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3390 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3402 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3410 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3414 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3416 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3424 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3431 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3437 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3449 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3461 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3472 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3476 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3480 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3483 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3496 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3504 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3510 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3516 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3520 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3525 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3532 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3538 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3550 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3560 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3573 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3596 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3608 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3618 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3626 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3638 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3644 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3656 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3668 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3688 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3693 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3696 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3705 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3718 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3730 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3742 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3752 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3764 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3768 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3801 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3808 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3816 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3820 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3826 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3838 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3843 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3855 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3864 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3870 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3883 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3907 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3932 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3944 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3952 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3969 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3976 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3984 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3988 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4000 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4006 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4018 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4030 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4032 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4039 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4050 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4056 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4068 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4080 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4086 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1391 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1420 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2258 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2266 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2272 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2285 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2291 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2297 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2308 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2314 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2320 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2326 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2347 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2366 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2372 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2384 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2387 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2399 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2407 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2428 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2440 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2448 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2459 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_2465 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2473 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2497 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2499 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2504 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2519 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2525 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2535 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2545 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_2551 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2569 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2576 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2582 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2600 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2606 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2617 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2624 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2630 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2636 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2642 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2648 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2654 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_2660 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2673 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2682 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_2690 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3093 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3101 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3114 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3120 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3126 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3132 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3143 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3149 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3155 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3160 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3164 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3170 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3184 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3202 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3214 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3218 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3232 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3244 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3254 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3267 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3288 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3304 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3316 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3320 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3328 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3344 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3356 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3364 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3375 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3388 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3393 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3399 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3411 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3429 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3441 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3444 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3449 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3453 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3458 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3464 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3472 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3487 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3493 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3500 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3506 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3510 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3515 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3527 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3551 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3556 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3572 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3578 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3590 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3602 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3610 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3616 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3630 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3636 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3647 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3653 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3659 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3668 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3684 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3698 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3709 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3715 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3736 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3760 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3772 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3778 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3816 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3828 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3848 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3860 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3866 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3878 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3904 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3916 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3924 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3928 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3940 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3960 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_3972 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3980 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3984 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_3993 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4011 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4023 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4035 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_4040 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4046 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_4060 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_4072 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_4078 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_4081 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1240 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1283 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1337 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1339 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1374 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1386 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1415 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2267 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2286 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2292 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2298 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2303 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2313 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2319 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2325 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2329 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2334 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2342 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2348 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2356 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2367 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2373 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2403 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2412 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2420 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2431 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2445 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2451 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2457 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2469 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2490 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2498 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2508 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2514 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2518 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2523 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2527 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_2531 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2545 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2552 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2558 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2564 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2570 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2580 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2589 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2597 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2609 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2622 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2628 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2634 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2648 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_2656 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_2664 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_2683 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3103 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3111 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3119 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3131 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3142 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3154 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3162 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3168 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3174 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3186 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3190 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3196 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3210 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3218 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3226 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3234 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3244 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3248 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3260 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3266 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3272 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3284 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3296 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3304 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3313 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3319 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3327 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3332 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3340 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3348 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3356 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3368 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3382 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3395 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3399 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3404 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3410 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3414 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3422 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3434 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3442 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3454 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3466 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3472 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3476 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3489 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3495 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3512 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3525 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3545 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3568 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3581 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3594 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3600 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3608 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3619 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3625 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3631 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3637 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3640 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3651 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3660 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3672 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3680 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3689 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3696 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3708 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3712 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3718 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3727 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3733 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3739 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3788 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3800 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3806 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3820 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3832 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3843 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3855 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3871 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3883 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3895 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3899 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_3908 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3916 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3920 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3926 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3937 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3963 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3976 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3982 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_3985 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3994 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4006 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4018 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_4030 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_4032 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_4042 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4052 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4064 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_4076 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1311 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1350 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1362 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2249 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2271 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2287 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2315 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2329 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2335 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2347 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2364 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2372 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2378 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2383 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2387 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2392 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2400 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2412 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2440 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2475 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2483 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2497 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2499 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2505 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2520 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2531 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2541 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_2551 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2555 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2559 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2571 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2581 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2590 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2598 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2606 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2611 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2615 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2621 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2635 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2641 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2646 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_2659 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_2665 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2667 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_2675 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_2690 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3093 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3119 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3127 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3142 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3153 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3161 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3179 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3187 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3199 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3205 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3213 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3231 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3235 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3241 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3252 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3266 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3272 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3280 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3292 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3306 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3312 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3322 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3326 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3329 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3332 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3338 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3350 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3362 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3370 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3378 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3384 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3388 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3394 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3400 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3410 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3422 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3427 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3435 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3444 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3450 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3458 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3468 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3485 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3491 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3497 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3500 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3505 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3513 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3517 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3527 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3539 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3551 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3556 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3560 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3566 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3576 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3592 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3601 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3607 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3612 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3618 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3624 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3630 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3638 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3651 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3657 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3704 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3716 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3722 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3724 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3730 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3741 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3765 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3777 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3780 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3788 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3791 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3799 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3807 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3812 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3818 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3830 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3848 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3860 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3872 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3878 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3884 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3890 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3930 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3942 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3945 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3948 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3956 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_3964 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_3969 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_3978 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_3986 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3989 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_4004 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_4009 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4015 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4027 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_4039 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4043 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4046 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4072 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_4084 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_4096 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4102 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1227 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1239 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1327 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1339 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1364 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1388 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2260 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2268 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2276 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2285 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2300 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2317 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2333 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2347 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2357 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2366 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2372 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2378 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2384 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2396 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2407 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2413 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2415 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2419 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2426 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2459 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2469 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_2471 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2489 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2509 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2514 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2524 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2540 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2544 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2550 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2558 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2568 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2580 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2591 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2601 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2607 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_2617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2623 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2633 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2637 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2643 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2649 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2660 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2670 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_2678 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_2682 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2692 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3101 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3109 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3121 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3128 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3134 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3147 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3160 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3168 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3174 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3184 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3190 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3192 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3196 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3202 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3214 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3231 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3241 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3248 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3255 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3274 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3286 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3291 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3297 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3304 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3309 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3318 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3326 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3329 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3349 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3355 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3360 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3364 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3370 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3376 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3379 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3390 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3398 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3413 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3420 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3432 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3444 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3452 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3456 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3459 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3463 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3466 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3470 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3472 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3478 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3488 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3501 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3512 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3523 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3536 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3542 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3548 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3554 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3560 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3568 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3573 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3579 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3588 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3592 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3597 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3606 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3615 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3624 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3630 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3652 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3676 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3688 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3708 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3720 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3724 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3730 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3739 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3788 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3800 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3803 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3808 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3814 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3817 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3824 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3836 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3850 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3858 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3862 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3864 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3868 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3874 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3880 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3886 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3898 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3910 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3918 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3956 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3968 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3974 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3976 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3988 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_3994 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4000 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_4006 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_4014 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4019 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_4028 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_4032 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_4038 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_4042 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4048 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4072 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1255 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1311 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1339 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1367 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1392 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1404 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1420 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2263 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2271 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2275 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2286 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2292 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2298 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2315 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2329 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2337 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2351 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2367 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2375 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2385 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2387 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2391 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2397 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2400 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2410 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2417 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2425 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2433 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_2439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2452 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2456 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2463 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2480 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2488 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2494 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2505 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_2509 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2521 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2527 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2541 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2549 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2553 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2568 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2576 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2584 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2592 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2598 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_2604 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2615 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2618 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2628 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2638 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2642 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2649 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2655 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2661 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_2665 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2677 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_2690 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3093 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3101 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3108 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3119 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3127 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3132 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3142 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3155 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3175 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3188 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3203 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3209 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3217 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3220 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3226 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3237 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3246 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3252 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3258 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3264 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3270 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3274 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3276 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3284 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3301 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3306 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3310 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3325 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3332 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3338 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3343 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3354 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3358 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3364 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3373 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3381 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3388 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3392 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3402 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3410 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3422 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3432 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3440 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3444 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3452 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3458 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3470 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3479 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3485 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3491 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3497 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3500 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3504 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3507 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3515 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3525 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3542 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3550 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3554 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3556 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3565 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3569 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3575 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3583 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3599 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3605 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3612 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3620 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3626 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3632 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3651 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3663 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3680 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3704 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3716 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3722 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3724 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3730 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3733 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3744 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3756 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3768 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3776 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3780 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3788 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3793 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3799 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3820 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3829 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3836 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3844 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3849 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3857 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3860 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3875 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3887 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3892 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3897 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3903 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3914 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3932 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3984 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3996 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4011 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4023 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4036 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_4048 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_4056 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_4066 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_4078 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_4081 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1352 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1386 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1408 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1414 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2262 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2266 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2271 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2282 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2288 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2300 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2307 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2311 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2323 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2329 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2338 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2344 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2356 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2363 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2369 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2382 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2395 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2407 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2433 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2436 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2447 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2451 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2454 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2460 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2468 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_2471 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2483 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2487 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2496 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2509 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2515 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2521 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2525 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2531 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2544 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2550 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2567 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2573 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2579 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2589 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2595 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_2601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2609 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2611 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2615 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2620 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2626 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2630 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2635 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2644 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2650 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2664 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_2667 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2671 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_2678 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_2691 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3089 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3093 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3103 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3127 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3152 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3158 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3174 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3185 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3192 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3196 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3202 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3213 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3232 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3244 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3252 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3258 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3264 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3270 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3273 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3276 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3287 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3296 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3304 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3310 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3322 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3330 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3332 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3337 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3341 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3347 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3353 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3360 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3364 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3370 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3382 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3386 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3388 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3399 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3403 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3406 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3410 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3413 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3416 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3422 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3428 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3437 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3444 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3452 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3464 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3470 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3472 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3476 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3482 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3494 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3498 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3500 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3504 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3512 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3522 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3526 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3532 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3538 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3544 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3552 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3556 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3560 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3575 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3590 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3596 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3604 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3609 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3612 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3616 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3622 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3630 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3633 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3640 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3652 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3696 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3708 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3720 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3724 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_3732 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3735 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3741 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3764 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3792 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3804 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3808 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3814 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3820 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3832 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3836 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3840 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3847 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3853 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3868 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3880 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3888 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3892 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3899 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3905 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3920 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3932 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3960 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3988 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4000 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4008 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_4020 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_4026 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_4029 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_4032 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_4053 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4060 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4072 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4084 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1225 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1347 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1359 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2263 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2273 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2275 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2283 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2295 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2315 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2321 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2327 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2331 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2335 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2343 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2348 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2352 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2355 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2366 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2372 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2378 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2384 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2393 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2413 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2417 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2424 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2440 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2443 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2455 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2459 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2462 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2470 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2485 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2496 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2503 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2509 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2515 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2523 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2529 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2540 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2546 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2552 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2559 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2565 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2571 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2574 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_2586 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2598 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2608 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2611 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_2615 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2623 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2628 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2634 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2640 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2652 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2658 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2664 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2672 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_2678 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_2690 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_2703 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3087 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3100 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3106 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3116 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3122 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3128 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3134 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3140 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3152 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3158 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3178 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3184 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3190 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3196 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3208 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3232 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3256 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3268 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3273 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3276 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3287 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3293 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3305 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3311 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3314 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3320 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3328 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3332 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3336 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3341 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3347 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3359 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3371 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3377 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3382 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3386 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3392 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3404 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3416 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3419 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3429 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3437 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3444 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3450 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3457 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3463 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3467 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3470 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3481 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3487 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3497 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3500 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3507 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3513 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3523 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3533 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3541 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3553 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3556 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3560 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3571 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3584 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3588 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3595 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3601 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3612 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3624 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3636 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3645 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3657 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3674 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3686 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3698 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3710 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3724 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3736 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3748 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3754 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3760 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3763 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3775 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3784 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3798 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3810 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3814 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3822 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3826 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3833 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3844 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3856 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3868 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3880 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3892 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3904 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3916 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3924 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3928 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3937 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3943 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3972 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3984 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_3990 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3994 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_4000 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4004 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4009 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4016 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4022 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_4034 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4042 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4047 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_4053 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4060 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_4065 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4071 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_4083 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1273 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1316 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1335 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1358 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1368 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1422 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2256 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2264 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2270 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2276 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2282 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2288 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2300 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2310 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2316 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2322 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2328 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2344 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2356 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2359 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2365 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2370 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2378 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2384 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2392 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2397 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2411 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2422 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2430 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2436 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2445 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2451 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2455 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2458 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2468 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2483 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2489 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2508 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2520 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2527 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2532 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2540 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2548 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2554 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_2560 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2572 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2580 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2583 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_2587 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2595 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2602 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2608 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2636 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2639 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2643 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2648 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2654 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_2660 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2668 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2674 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2680 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2692 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3082 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3089 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3097 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3104 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3110 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3122 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3128 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3134 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3136 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3160 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3178 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3192 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3204 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3241 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3248 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3260 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3272 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3275 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3291 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3304 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3312 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3323 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3335 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3347 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3351 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3360 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3364 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3367 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3376 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3384 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3396 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3408 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3414 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3416 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3428 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3433 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3441 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3465 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3472 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3477 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3483 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3495 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3499 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3511 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3515 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3525 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3538 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3549 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3559 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3565 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3571 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3584 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3588 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3594 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3604 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3616 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3628 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3636 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3640 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3652 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3664 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3676 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3688 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3694 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3696 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3708 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3711 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3723 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3735 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3740 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3746 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3749 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3752 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3759 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3766 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3772 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3777 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3786 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3794 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3802 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3806 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3808 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3818 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3830 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3843 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_3855 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3864 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3868 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3871 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3879 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3885 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3896 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3908 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3913 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3920 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_3924 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3944 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3956 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3968 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3974 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3988 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4000 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4006 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_4013 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_4019 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4023 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4032 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_4047 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4053 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4065 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_4077 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1294 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1348 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1390 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1400 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1403 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1424 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2265 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2271 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2275 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2284 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2292 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2304 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2310 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2316 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2324 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2328 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2340 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2348 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2354 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2367 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2373 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2385 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2387 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2399 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2403 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2406 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2412 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2418 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2424 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2432 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2455 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2477 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2489 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2497 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2504 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2513 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2530 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2534 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2541 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2547 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2553 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_2559 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2571 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2579 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2588 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2594 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_2607 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2611 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2615 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2621 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2627 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2654 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_2660 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2671 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_2675 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2678 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2684 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_2692 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_2703 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3082 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3093 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3101 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3108 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3112 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3118 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3124 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3130 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3142 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3146 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3149 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3155 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3164 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3169 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3175 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3179 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3182 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3194 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3206 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3218 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3220 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3232 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3256 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3268 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3274 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3291 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3318 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3330 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3332 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3340 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3348 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3352 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3367 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3379 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3388 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3396 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3409 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3421 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3433 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3456 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3460 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3468 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3474 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3480 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3488 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3494 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3500 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3512 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3524 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3527 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3545 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3551 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3556 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3560 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3566 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3572 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3585 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3591 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3597 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3600 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3612 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3624 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3632 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3635 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3648 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3660 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3668 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3680 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3692 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3704 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3710 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3721 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3724 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3732 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3738 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3744 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3756 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3768 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3776 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3780 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3784 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3796 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3808 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3820 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3828 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3832 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3836 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3840 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3852 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3864 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3876 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3892 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3904 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3907 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3915 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3926 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3938 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_3946 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3948 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3960 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3972 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3984 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_3996 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4004 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4010 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4014 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4017 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4031 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4043 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4055 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_4060 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_4072 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4078 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_4081 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_982 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1263 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1336 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1360 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1368 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1374 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2287 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2295 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2301 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2307 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2313 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2322 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2330 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2342 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2350 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2356 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2370 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2374 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2387 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2397 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2410 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2420 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2434 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2446 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2451 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2460 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2466 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_2481 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2495 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2513 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2516 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2524 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2527 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2533 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2537 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2544 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2552 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2558 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_2566 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2574 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2580 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2583 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2587 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_2611 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2618 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2629 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_2635 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2651 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2662 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2672 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_2678 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2692 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2695 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_2703 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3082 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3086 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3096 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3102 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3112 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3118 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3124 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3130 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3133 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3136 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3147 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3156 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3168 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3176 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3179 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3192 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3196 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3208 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3220 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3226 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3232 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3244 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3248 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3255 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3261 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3267 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3273 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3285 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3297 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3301 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3304 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3310 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3316 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3322 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3330 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3334 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3342 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3350 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3353 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3360 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3372 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3384 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3396 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3408 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3411 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3416 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3428 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3440 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3458 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3468 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3472 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3478 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3484 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3490 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3496 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3508 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3520 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3526 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3528 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3534 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3543 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3547 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3570 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3577 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3584 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3596 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3608 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3616 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3621 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3630 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3636 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3640 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3648 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3666 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3680 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3692 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3696 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3701 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3707 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3716 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3722 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3728 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3740 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3748 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3752 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3764 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3776 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3788 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3800 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3805 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3808 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3813 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3819 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3830 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3838 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3843 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3851 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3864 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3876 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_3888 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3899 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3911 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3915 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3920 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_3928 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3933 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3941 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3955 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_3967 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3976 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3985 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3997 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_4009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4017 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_4021 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4029 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_4032 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_4040 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4050 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4062 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4074 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4086 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_4088 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_4100 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1168 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1299 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1398 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2263 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2271 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2281 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2293 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2298 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2310 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2314 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2319 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2327 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2331 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2339 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2353 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2357 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2373 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2379 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2385 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2387 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2393 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2412 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2422 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2430 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2434 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2439 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2443 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2451 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2455 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2463 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2469 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2488 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2494 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2499 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2507 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2510 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2524 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2539 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2548 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2555 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2559 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2565 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_2570 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2583 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2591 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2599 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2607 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2611 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2619 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2625 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2636 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2639 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2652 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2658 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2664 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2673 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2692 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2695 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2711 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2719 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2723 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2731 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2740 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2748 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2751 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2758 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2768 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2776 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2790 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2794 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2804 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2818 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2831 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2843 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2857 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2861 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2869 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2873 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_2883 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2889 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2891 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2902 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2906 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2916 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2930 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_2943 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2958 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2966 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2972 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_2975 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_2986 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2990 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3000 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3003 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3007 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3011 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3021 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3027 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3031 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3042 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3052 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3059 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3071 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3081 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3085 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3087 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3091 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3095 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3102 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3108 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3115 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3122 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3130 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3140 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3143 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3161 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3165 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3168 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3171 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3177 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3189 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3193 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3211 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3223 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3227 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3233 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3246 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3252 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3255 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3266 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3281 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3283 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3297 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3311 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3315 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3327 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3335 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3339 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3351 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3363 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3373 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3385 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3393 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3395 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3409 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3420 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3429 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3441 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3449 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3451 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3459 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3462 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3474 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3479 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3490 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3502 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3507 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3519 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3535 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3541 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3548 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3554 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3563 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3567 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3580 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3588 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3591 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3603 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3615 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3619 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3626 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3632 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3638 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3642 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3647 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3659 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3671 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3675 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3679 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3684 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3696 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3703 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3715 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3728 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3731 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_3757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3771 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3783 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3787 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3799 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3804 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3815 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3827 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3833 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3839 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3843 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3855 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3871 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3883 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3895 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3899 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3912 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3924 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3927 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3932 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3938 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_3950 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3955 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3967 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_3979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3998 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4011 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4023 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_4026 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4030 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_4033 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_4039 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4045 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4057 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4065 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4067 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_4079 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_4091 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_982 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2263 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2287 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2293 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2299 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2303 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2315 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2321 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2324 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2332 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2338 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2344 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2349 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2355 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2363 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2369 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2377 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2389 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2409 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2412 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2415 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2421 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2447 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2455 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2461 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2465 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2468 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2495 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2504 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2510 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2522 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2527 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2532 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2538 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2549 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2555 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2566 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2572 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2580 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2583 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2587 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2595 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2609 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2615 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2625 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2637 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_2643 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2655 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2663 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2674 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2680 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2692 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2695 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2702 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2708 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2716 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2725 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2733 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2739 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2743 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2748 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2751 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2755 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2759 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2780 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2791 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2804 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2818 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2822 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2830 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2842 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2848 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2858 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2871 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2903 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_2911 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_2917 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2930 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2938 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2951 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_2959 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_2971 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_2975 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2983 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_2991 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3002 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3015 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3028 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3031 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3039 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3043 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3050 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3062 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3070 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3078 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3084 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3087 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3098 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3104 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3112 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3123 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3126 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3132 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3139 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3143 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3150 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3156 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3168 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3182 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3211 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3252 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3255 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3261 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3269 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3282 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3294 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3298 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3308 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3311 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3323 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3327 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3339 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3353 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3362 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3367 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3378 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3390 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3402 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3410 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3413 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3421 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3435 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3458 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3464 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3476 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3479 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3490 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3502 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3514 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3520 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3523 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3532 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3535 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3542 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3548 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3564 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3576 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3588 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3591 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3603 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3627 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3635 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3639 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3647 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3659 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3675 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3687 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3699 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3703 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3708 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3718 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3724 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3733 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3741 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3750 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3771 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3791 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3803 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3811 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3815 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3827 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3851 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3863 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3871 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3883 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3907 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3919 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3925 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3934 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3946 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3954 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3963 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3975 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3981 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3995 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4007 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4019 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_4022 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_4031 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_4037 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4039 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_4044 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4050 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4062 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_4074 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_4086 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1210 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1228 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2255 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2261 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2273 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2275 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2282 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2288 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2300 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2305 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2329 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2331 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2345 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2357 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2369 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2381 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2387 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2395 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2419 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2431 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2443 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2455 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2467 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2479 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2491 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2497 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2499 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2511 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2525 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2537 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2549 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2553 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2555 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2563 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2569 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2581 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2599 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2609 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2611 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2621 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2627 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2632 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_2644 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_2656 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2664 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_2667 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2672 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2693 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2696 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2710 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2716 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2723 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2727 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2733 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2747 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2753 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2761 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2770 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2776 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2787 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2796 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2806 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2816 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2822 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2826 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2832 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2842 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2848 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2852 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2859 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2867 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2875 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2879 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2884 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2891 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2905 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2911 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2917 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2928 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2936 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2942 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2953 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_2967 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2972 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2980 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_2990 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3000 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3003 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3015 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3034 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3038 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3043 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3049 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3055 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3059 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3065 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3071 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3079 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3083 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3089 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3095 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3113 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3115 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3127 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3151 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3163 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3169 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3171 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3183 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3207 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3225 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3227 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3239 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3247 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3252 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3256 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3259 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3268 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3275 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3281 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3283 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3289 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3294 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3300 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3316 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3322 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3326 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3336 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3339 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3351 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3375 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3393 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3395 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3413 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3425 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3432 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3444 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3451 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3456 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3468 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3480 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3486 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3498 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3507 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3519 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3537 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3549 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3555 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3561 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3563 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3575 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3599 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3611 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3617 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3619 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3631 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3643 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3655 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3663 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3669 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3673 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3675 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3687 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3697 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3706 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3714 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3719 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3723 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_3727 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3731 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3743 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3755 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3767 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3772 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3778 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3787 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3795 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3807 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3819 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3824 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3830 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3843 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3855 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3879 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3891 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3897 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3899 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3911 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3923 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3930 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3942 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3955 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3967 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3979 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3991 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3995 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_4004 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4011 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4023 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4035 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_4050 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_4056 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4064 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_4067 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_4081 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1381 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1423 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2253 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2265 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2278 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2284 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2296 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2303 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2315 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2327 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2343 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2346 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2355 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2359 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2363 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2375 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2387 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2399 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2411 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2427 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2445 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2448 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2456 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2468 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2471 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2483 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2495 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2507 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2517 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2523 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2563 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2575 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2583 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2595 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2607 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2619 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2631 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2637 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2651 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2663 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2675 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2692 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2695 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2699 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2705 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_2715 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2727 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2733 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2739 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2745 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2749 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2751 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2755 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2758 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2767 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2777 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2787 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2797 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2803 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2807 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2814 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2822 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2829 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2837 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2849 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2857 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2861 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2863 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_2867 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2880 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2884 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2909 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2915 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_2919 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2923 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2929 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2934 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2940 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2946 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2952 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_2958 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2964 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2969 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2973 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_2975 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2982 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2986 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_2991 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_2995 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3001 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3011 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3023 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3029 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3031 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3037 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3045 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3051 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3055 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3061 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3067 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3079 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3084 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3087 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3117 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3141 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3155 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3179 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3191 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3197 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3199 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3211 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3235 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3247 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3253 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3255 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3267 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3270 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3288 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3300 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3308 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3311 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3323 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3347 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3359 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3365 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3379 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3403 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3415 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3421 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3435 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3459 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3471 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3477 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3479 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3484 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3490 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3502 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3514 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3526 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3535 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3547 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3571 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3583 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3589 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3591 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3603 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3627 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3639 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3647 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3659 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3671 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3679 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3685 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3691 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3699 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3703 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3715 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3739 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3751 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3757 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3759 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3771 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3783 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3789 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3792 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3813 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3815 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3827 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3835 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3848 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3860 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3868 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3871 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3883 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3887 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3899 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3903 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3907 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3911 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3917 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3925 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3927 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3939 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3963 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3975 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_3981 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3983 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3995 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4019 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4031 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4037 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_4039 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4045 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_4048 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4069 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4093 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_4095 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1442 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1450 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1467 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1507 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1510 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1519 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1533 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1547 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1557 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1561 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1597 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1604 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1629 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1638 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1646 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1669 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1673 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1687 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1709 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1718 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1735 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1737 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1741 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1772 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1780 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1788 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1797 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1801 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1821 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1841 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1846 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1860 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1866 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1874 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1886 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1892 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1911 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1925 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1939 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1947 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1956 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1968 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1978 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1993 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2006 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2028 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2034 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2056 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2062 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2079 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2085 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2098 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2107 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2127 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2137 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2143 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2147 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2154 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2169 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2196 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2211 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2220 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2232 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2238 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2241 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2247 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2263 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2281 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2364 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2370 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2378 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2393 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2414 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2432 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2437 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2457 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2465 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2483 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2488 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2493 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2505 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2516 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2533 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2561 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2565 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2570 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2577 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2586 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2598 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2605 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2613 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2623 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2737 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2742 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2745 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2751 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2756 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2762 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2768 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2787 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2795 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2799 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2808 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_2814 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2820 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2843 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2853 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2875 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_2881 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2889 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2895 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2901 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2911 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2919 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2925 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2929 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2932 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2938 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2945 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2951 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2957 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2963 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2967 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2973 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2979 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_2985 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_2989 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2994 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3003 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3009 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3019 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3023 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3029 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3035 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3041 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3047 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3051 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3063 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3069 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3075 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3079 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3085 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3091 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3121 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3205 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3317 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3345 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3373 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3401 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3457 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3485 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3501 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3517 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3541 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3569 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3597 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3625 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3637 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3646 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3658 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3666 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3681 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3688 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3709 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3737 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3765 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3781 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3796 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3833 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3837 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_3841 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3844 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3853 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3877 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3905 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3933 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3961 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4017 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1374 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1438 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1499 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1508 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1531 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1539 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1550 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1558 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1577 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1601 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1609 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1641 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1657 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1687 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1695 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1715 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1722 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1735 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1747 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1753 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1759 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1767 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1773 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1778 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1784 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1790 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1803 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1814 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1820 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1826 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1835 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1847 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1856 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1864 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1872 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1878 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1886 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1905 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1911 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1923 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1931 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1935 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1941 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1950 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1958 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1967 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1975 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1985 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1991 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1996 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2015 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2023 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2028 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2036 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2044 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2052 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2071 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2079 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2087 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2095 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2103 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2119 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2125 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2144 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2148 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2153 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2169 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2183 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2191 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2195 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2201 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2215 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2365 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2377 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2391 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2397 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2405 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2409 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2414 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2420 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2426 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2438 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2450 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2462 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2465 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2477 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2485 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2503 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2515 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2518 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2527 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2539 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2551 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2563 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2709 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_2721 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2733 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2741 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2745 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2751 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2754 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2760 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2763 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2784 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2792 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2798 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2819 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2825 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2831 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2837 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2845 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2851 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2861 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2867 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2875 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2879 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2882 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2888 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2894 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2900 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2904 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2913 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_2930 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_2936 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2947 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2953 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2959 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2965 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2974 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_2980 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2990 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_2996 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3002 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3008 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3014 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3020 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3025 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3029 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3039 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3048 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3054 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3060 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3072 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3117 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3123 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3303 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3311 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3318 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3324 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3336 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3348 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3585 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3597 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3607 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3627 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3863 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1278 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1353 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1459 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1522 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1526 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1559 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1567 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1593 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1603 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1608 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1616 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1626 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1632 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1649 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1653 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1657 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1671 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1677 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1683 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1695 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1707 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1713 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1717 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1720 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1724 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1729 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1735 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1739 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1744 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1750 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1762 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1770 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1776 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1800 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1833 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1845 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1855 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1862 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1868 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1874 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1883 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1896 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1902 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1910 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1920 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1928 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1939 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1948 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1956 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1964 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1969 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1977 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1983 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1987 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1989 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1995 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2008 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2020 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2028 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2036 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2041 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2045 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2051 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2061 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2069 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2077 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2101 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2107 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2119 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2127 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2135 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2143 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2151 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2155 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2163 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2171 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2181 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2189 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2195 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2201 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2267 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2275 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2281 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2289 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2300 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2306 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2318 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2603 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2605 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2613 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2620 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2626 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_2638 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2646 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2650 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2658 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2753 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2760 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2764 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2767 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2773 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2777 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2783 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2786 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2790 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2795 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2807 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2819 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2829 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2833 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2841 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2853 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2859 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2865 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2871 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2957 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_2963 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2975 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_2984 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_2990 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3001 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3007 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3019 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3031 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3043 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3357 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3369 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3376 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3457 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3477 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3489 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3525 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_3536 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3542 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3554 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1268 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1450 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1467 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1479 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1517 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1531 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1538 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1546 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1560 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1566 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1575 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1587 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1593 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1600 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1608 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1619 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1631 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1639 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1642 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1648 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1654 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1662 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1670 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1674 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1681 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1689 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1699 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1711 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1723 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1749 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1761 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1769 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1772 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1784 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1847 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1849 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1855 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1858 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1864 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1872 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1876 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1884 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1892 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1915 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1927 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1932 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1938 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1942 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1945 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1967 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1973 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1979 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1982 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1992 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2002 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2008 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2014 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2022 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2030 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2040 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2048 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2052 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2058 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2062 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2067 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2071 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2079 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2091 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2103 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2119 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2123 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2126 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2135 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2140 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2148 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2153 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2167 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2183 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2185 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2189 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2195 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2198 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2204 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2216 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2228 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2593 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2605 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2613 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2618 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2626 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2669 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2693 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2705 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2765 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2770 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2778 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2784 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2788 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2791 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2805 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2811 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2817 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2823 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2835 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2847 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2893 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2900 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_2910 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2981 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2987 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_2999 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3011 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3037 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3049 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3057 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3063 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3069 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3247 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_3255 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1482 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1535 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1538 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1551 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1561 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1569 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1577 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1594 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1603 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1606 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1616 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1627 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1633 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1640 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1661 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1666 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1690 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1702 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1706 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1821 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1833 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1841 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1863 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1875 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1877 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1881 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1890 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1906 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1951 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1963 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1989 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1997 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2000 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2008 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2018 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2024 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2032 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2035 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2042 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2051 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2065 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2071 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2077 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2083 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2089 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2101 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2113 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2124 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2128 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2131 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2135 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2138 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2146 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2155 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2167 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2173 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2197 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2209 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2217 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2224 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2230 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2242 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2254 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2266 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2339 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2351 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2359 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2366 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2372 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2393 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2397 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2402 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2408 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2420 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2432 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2461 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2473 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2479 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2483 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2517 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_2529 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2536 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2542 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2555 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2771 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2773 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2777 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2780 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2786 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2792 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2798 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2806 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2811 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2817 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2823 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2827 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2833 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_2845 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2853 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2864 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2870 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2882 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2953 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_2957 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_2960 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2970 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2982 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_2994 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3555 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3563 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3569 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3581 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3586 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3592 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3604 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3667 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3674 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3680 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3692 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3704 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3716 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_4073 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1501 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1591 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1805 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1843 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1846 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1856 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1870 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1882 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1890 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1965 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1973 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1977 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1991 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2004 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2010 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2023 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2035 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2047 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2063 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2095 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2107 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2123 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2126 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2147 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2159 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2171 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2321 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2329 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2335 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2343 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2415 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2427 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2439 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2451 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2471 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2481 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2487 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2499 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2631 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_2639 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_2967 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2978 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_2990 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3002 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3014 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3022 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3415 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_3423 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1443 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1565 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1585 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1591 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1628 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1640 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1677 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1685 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1692 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1799 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1811 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1845 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1853 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1866 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1883 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1899 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1911 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1923 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1981 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1986 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1993 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2019 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2031 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2051 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2057 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2065 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2125 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2137 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2143 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2155 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_2157 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_2165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2170 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2182 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2194 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2225 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_2242 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2255 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2262 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2285 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_2321 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2339 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2363 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2375 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2953 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_2965 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2972 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2984 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3333 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3345 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3351 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3354 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3367 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_3379 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1623 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1631 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1636 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1660 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1829 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1849 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1857 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1862 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1874 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1886 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1892 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1997 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2141 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2153 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2168 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2225 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2309 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2329 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2341 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2377 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_2389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2406 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2413 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2425 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2449 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2461 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2472 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2478 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2490 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2494 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2498 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2504 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_2516 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2669 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_2681 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2686 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2695 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2707 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2719 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2731 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3273 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3285 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3289 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3294 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3300 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3999 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4011 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_4023 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1633 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1645 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1745 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1757 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1819 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1821 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1829 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1841 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1855 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1867 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1933 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1963 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1987 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1989 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1997 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2009 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2021 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_2033 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2121 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2133 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_2145 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_2153 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2785 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_2797 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_2808 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2814 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_2826 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3245 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3252 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3258 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3270 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3389 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_3401 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3411 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3424 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_3436 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3555 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3563 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_4073 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1471 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1681 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1693 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1699 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1710 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1722 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1743 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1755 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1767 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1779 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1793 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1813 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1825 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1829 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1861 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1873 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1881 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1884 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1959 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1967 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1997 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2029 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2041 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2049 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2052 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2064 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2073 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2081 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2086 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2100 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2112 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2124 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2136 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_2142 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_2150 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2161 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2167 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3005 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3021 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3029 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3041 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3385 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3403 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3415 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3430 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3442 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3454 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3466 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3527 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3529 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3537 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_3544 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3550 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3562 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3574 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_3582 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1476 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1573 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1707 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1709 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1717 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1777 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1791 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1799 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1803 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1806 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1875 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1883 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1888 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1900 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1904 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1907 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1919 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2043 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2045 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2051 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2056 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2068 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2080 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_2092 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_2106 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2112 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2124 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2136 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_2148 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_2164 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2170 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2182 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2194 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2206 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_2337 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2341 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2357 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_2369 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3221 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3233 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3239 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3244 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3250 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3262 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3421 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_3433 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3793 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3807 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3816 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3822 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3834 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3893 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_3905 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_3911 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4038 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_4050 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_4058 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1328 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1555 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1623 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1625 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1632 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1715 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1723 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1737 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1758 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1770 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1788 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1797 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1815 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1827 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1839 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1873 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1885 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1891 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2309 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2324 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2336 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2348 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2360 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2366 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2372 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2382 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2388 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2400 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2757 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2837 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2845 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_2851 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2861 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2873 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2897 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2913 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2935 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2947 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_2959 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3217 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3243 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3247 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3253 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3265 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3277 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3297 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3367 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3845 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3857 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3862 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_3872 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3878 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3884 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3888 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3900 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3912 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_4031 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4040 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4052 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4064 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4076 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1416 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1464 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1621 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1630 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1653 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1672 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1678 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1690 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1702 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1727 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1739 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1800 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1812 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1818 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1827 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1839 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1851 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1863 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2013 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2025 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2030 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2042 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2069 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2081 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2092 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2211 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2213 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2219 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2229 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2235 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2247 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_2259 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2267 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2273 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2276 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2288 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2294 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_2311 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2322 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2337 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2349 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2364 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_2370 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_2378 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2885 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_2907 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2917 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3009 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3021 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3026 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3034 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3046 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3053 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3073 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3078 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3090 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3102 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3163 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3183 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3277 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3289 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3295 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3708 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3720 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3849 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3869 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3881 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3889 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3898 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3916 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3928 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_3940 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_4073 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1267 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1527 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1535 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1540 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1552 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1564 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1577 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1583 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1599 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1612 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1618 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1658 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1664 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1676 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1705 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1717 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1725 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1732 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1753 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1773 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1883 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1895 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2015 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2023 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2127 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2134 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2140 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2152 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2164 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2176 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2197 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_2205 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2211 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2217 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2229 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2241 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2254 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2268 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2286 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_2294 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2309 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2327 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2339 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2477 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2489 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2497 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2503 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2515 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2655 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2869 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_2879 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2889 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_2901 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3845 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3857 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_3861 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3874 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3880 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3892 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3904 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3908 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1393 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1502 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1514 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1526 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1554 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1566 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1578 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1612 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1620 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1632 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1789 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1796 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1802 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1814 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1889 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1893 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1898 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1904 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1916 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1928 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1945 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1964 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1970 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1978 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2013 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2025 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_2033 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_2057 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2065 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_2082 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_2088 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2094 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2629 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_2641 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2649 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2673 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_2685 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2692 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2704 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3163 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3170 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3176 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3188 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3200 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3212 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4029 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_4041 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4045 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_4049 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1252 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1500 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1510 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1637 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1645 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1648 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1662 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1674 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1695 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1701 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1713 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1721 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1727 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1791 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1801 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1917 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1935 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1947 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2127 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_2129 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_2137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2143 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2167 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2183 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2196 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2208 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2220 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_2232 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2505 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2633 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2645 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_2656 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2662 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2674 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_2686 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2696 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2708 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2720 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2732 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3037 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3041 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3044 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3058 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3070 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_3078 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3093 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3118 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3130 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3485 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3497 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_3505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3518 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3524 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1468 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1536 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1564 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1572 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1582 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1588 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1597 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1605 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1608 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1616 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1628 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1632 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1651 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1763 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1765 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1771 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1776 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1782 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1794 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1806 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1833 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1845 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1851 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1854 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2001 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2010 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2022 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_2034 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_2042 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2056 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2068 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2080 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2113 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2125 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_2132 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_2146 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_2154 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_2995 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_2997 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3003 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3006 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3018 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3030 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3042 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_3050 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3345 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3364 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3376 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3400 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3406 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3410 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3427 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3439 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3569 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3588 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3600 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3949 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3961 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3964 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3978 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3990 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4002 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1249 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1267 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1318 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1437 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1445 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1545 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1548 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1555 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1559 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1573 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1585 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1589 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1599 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1611 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1625 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1633 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1773 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1781 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1787 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1793 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1808 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1812 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1815 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1823 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1835 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1847 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1849 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1857 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1862 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1868 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1880 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1892 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1985 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1991 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1994 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2014 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2017 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_2029 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2037 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2044 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2050 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_2062 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2070 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2141 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2145 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2148 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2162 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_2174 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2182 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2389 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_2392 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_2406 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_2981 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_2993 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_2999 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3004 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3018 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3043 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3055 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3067 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3134 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3141 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3153 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3247 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3256 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3262 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3274 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3286 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3298 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3359 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3367 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3371 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3376 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3388 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3400 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3412 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3453 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3465 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3470 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3479 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3491 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3515 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3583 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3592 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3604 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3616 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3628 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3665 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_3677 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3683 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3777 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3793 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3799 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_4087 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_4094 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1362 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1441 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1456 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1459 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1556 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1570 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1582 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1594 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1609 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1647 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1665 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1677 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1683 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1704 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1789 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1806 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1812 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1816 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1825 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1931 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1943 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1951 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1963 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1975 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2213 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2225 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_2233 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2247 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_2259 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2853 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2865 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2871 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_2882 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_2995 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_2997 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3008 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3020 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3032 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3044 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3301 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3313 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3321 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3326 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3849 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3872 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_3884 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1314 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1559 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1567 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1584 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1590 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1602 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1614 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1622 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1632 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1644 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1656 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1668 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1681 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1699 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1711 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1723 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1793 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1805 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1812 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1818 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1830 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1842 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1929 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1941 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1946 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3751 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_3766 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3772 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3784 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3796 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3863 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3865 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3871 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3882 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3894 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3906 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3918 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1225 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1338 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1344 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1651 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1653 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1659 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1667 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1691 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1703 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1906 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1930 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1945 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1969 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2281 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_2293 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_2301 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2307 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_2319 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2529 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2549 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2567 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2579 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2591 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_2610 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2616 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2628 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2640 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_2652 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3065 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3089 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3201 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_3213 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3218 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3443 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3451 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3723 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3725 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3733 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3743 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3767 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1340 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2029 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_2085 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2093 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2098 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2104 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2116 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2141 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_2153 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_2161 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2173 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2221 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3229 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_4087 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_4097 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1169 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1281 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1406 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1440 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1482 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1502 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1520 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1613 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1631 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1665 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1677 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1685 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1690 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1704 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1765 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1783 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1786 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1790 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1875 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1888 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1894 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1906 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1918 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1930 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1939 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1945 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1957 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1968 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1974 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1986 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2043 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_2045 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2050 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2056 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2068 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2080 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2092 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_2181 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2194 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2200 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2349 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2361 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2375 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2435 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2437 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2445 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2448 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2456 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2459 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2471 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2505 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2517 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2529 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_2543 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2697 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2773 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2793 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2805 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_2817 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3051 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3069 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3093 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3625 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3779 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3785 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3797 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3885 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_3947 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3953 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3965 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_4073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_4085 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1360 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1417 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1421 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1461 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1569 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1589 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1629 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1635 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1645 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1673 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1678 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1687 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1690 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1702 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1714 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1749 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1785 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1790 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1799 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1813 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1861 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1873 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1878 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1884 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1890 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1902 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1905 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1911 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1917 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1957 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1961 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1971 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1981 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2001 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2013 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2025 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2037 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2085 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2093 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2099 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2105 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2111 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2125 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2145 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2168 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2174 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2180 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2185 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2217 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2229 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2237 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2265 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2277 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2287 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2321 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2341 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2351 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2385 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2397 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2433 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2441 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2446 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2453 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2489 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2511 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_2517 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2525 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2545 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2553 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2559 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2571 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2575 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2581 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2687 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2719 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2731 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2739 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2743 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2749 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2775 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2779 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2782 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2796 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2825 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2837 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2845 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2855 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2887 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2899 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2911 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2943 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_2955 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_2963 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_2967 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_2993 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3005 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3013 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3023 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3049 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3055 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3064 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3070 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3076 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3085 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3117 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3131 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3137 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3149 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3159 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3163 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3174 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3180 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3186 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3193 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3237 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3245 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3291 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3329 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3341 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3359 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3361 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3365 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3385 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3394 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3400 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3408 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3411 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3415 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3421 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3441 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3455 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3467 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3497 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3509 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3517 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3527 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3533 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3583 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3609 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3621 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3635 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3639 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3645 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3657 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3669 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3681 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3695 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3697 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3741 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3749 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3792 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3798 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3804 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3833 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3845 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3853 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3863 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3869 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3919 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3921 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3945 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3952 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3958 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3966 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_3971 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1393 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1425 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1449 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1517 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1561 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1585 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1589 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1594 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1617 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1649 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1653 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1661 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1665 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1685 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1709 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1729 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1765 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1785 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1809 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1817 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1821 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1829 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1833 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1853 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1873 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1877 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1897 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1929 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1933 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1953 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1977 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1985 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1989 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1997 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2001 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2021 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2041 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2045 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2065 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2077 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2097 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2121 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2141 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2153 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2175 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2195 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2211 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2233 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2265 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2289 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2309 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2325 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2343 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2363 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2375 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2378 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2401 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_2425 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2431 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2434 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2457 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2477 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2487 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2490 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2511 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2531 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2543 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2546 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2549 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2569 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2593 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2625 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2645 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2657 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2679 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2699 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2706 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2712 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2737 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2769 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2793 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2867 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2873 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_2881 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2885 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2905 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2929 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2935 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2939 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2961 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_2981 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_2987 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_2995 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3015 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3035 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3041 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3045 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3050 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3053 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3073 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3097 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3105 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3129 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3149 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3163 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3183 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3203 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3209 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3217 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3221 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3241 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3271 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3274 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3297 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3317 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3323 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3331 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3351 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3371 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3377 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3385 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3389 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3409 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3433 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3439 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3443 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3465 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3485 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3497 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3519 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3539 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3545 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3553 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3557 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3577 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3607 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3611 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3633 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3687 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3707 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3713 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3719 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3722 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3725 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3745 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3769 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_3775 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3778 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3801 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3821 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3833 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3855 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3875 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3881 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3889 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3893 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3913 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_3937 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_3945 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3949 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_3969 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3989 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_4001 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4023 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4047 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_4085 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4097 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1286 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1405 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1454 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1482 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1510 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1518 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1538 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1546 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1573 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1593 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1597 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1601 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1605 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1622 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1630 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1650 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1653 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1661 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1678 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1686 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1706 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1714 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1734 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1741 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1761 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1765 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1769 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1773 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1790 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1798 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1818 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1821 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1829 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1846 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1854 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1874 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1881 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1885 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1902 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1905 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1938 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1958 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1961 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1969 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1986 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1989 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1994 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2014 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2022 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2042 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2045 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2053 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2070 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2073 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2091 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2099 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2119 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2125 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2147 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2151 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2154 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2157 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2175 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2179 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2182 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2185 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2203 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2211 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2213 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2239 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2241 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2259 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2267 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2287 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2294 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2297 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2315 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2323 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2325 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2343 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2351 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2353 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2371 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2379 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2381 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2399 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2407 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2409 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2427 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2435 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2437 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2455 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2462 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2483 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2487 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2490 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2493 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2511 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2519 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2539 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2543 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2546 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2567 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2571 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2574 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2577 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2595 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2603 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2623 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2627 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2630 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2633 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2651 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2659 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2661 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2679 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2687 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2707 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2735 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2741 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2745 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2763 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2771 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2791 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2801 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2819 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2825 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2829 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2847 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2855 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_2875 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2883 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2903 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2909 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2931 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2937 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2959 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2965 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2969 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_2987 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_2993 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_2997 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3015 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3021 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3043 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3049 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3053 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3071 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3075 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3078 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3081 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3099 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3107 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3109 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3127 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3135 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3155 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3162 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3165 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3183 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3191 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3211 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3217 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3239 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3245 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3267 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3273 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3295 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3299 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3302 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3305 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3323 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3331 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3351 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3357 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3361 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3379 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3387 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3389 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3407 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3415 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3435 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3441 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3445 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3463 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3471 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3491 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3519 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3525 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3529 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3547 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3553 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3575 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3581 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3603 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3609 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3631 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3637 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3659 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3663 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3666 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3669 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3687 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3695 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3715 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3721 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3725 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3743 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3751 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3771 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3777 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3781 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3799 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3807 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3827 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3833 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3855 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3861 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3865 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3883 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3891 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3911 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3917 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3921 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_3939 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_3945 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3949 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3967 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_3975 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_3977 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3995 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4003 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4005 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_4023 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4045 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_4073 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_4085 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4089 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4101 ();
endmodule
