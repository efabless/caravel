* NGSPICE file created from caravan.ext - technology: sky130A

.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VPWR Y VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_93# a_229_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_229_47# a_27_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_229_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfbbn_2 CLK_N D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_790_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_790_47# a_944_21# a_650_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 Q_N a_1431_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_894_329# a_476_47# a_650_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_476_47# a_27_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_650_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_2236_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_650_21# a_560_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1547_47# a_944_21# a_1431_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 Q a_2236_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1115_329# a_650_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_476_47# a_193_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_584_47# a_27_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 VPWR a_944_21# a_894_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_1162_47# a_650_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 VGND a_1431_21# Q_N VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Q a_2236_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND a_1431_21# a_2236_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR RESET_B a_944_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 Q_N a_1431_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR a_1431_21# a_1343_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR a_944_21# a_1665_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 VGND a_1431_21# a_1366_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND a_2236_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_1431_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VPWR a_1431_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1366_47# a_193_47# a_1257_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X30 a_1665_329# a_1257_47# a_1431_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 a_1257_47# a_27_47# a_1162_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X33 a_1343_413# a_27_47# a_1257_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1547_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_650_21# a_476_47# a_790_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1257_47# a_193_47# a_1115_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_1431_21# a_1257_47# a_1547_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 a_650_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X40 VPWR a_1431_21# a_2236_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 VGND RESET_B a_944_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 a_560_413# a_193_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X43 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VPWR X VNB VPB
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VPWR X VNB VPB
X0 a_204_297# A1 a_396_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR S a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_396_47# A0 a_314_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_206_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_396_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_396_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_490_47# A1 a_396_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND S a_490_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_396_47# A0 a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_396_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR S a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_396_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND S a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_0 A B VGND VPWR X VNB VPB
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VPWR X VNB VPB
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=5.36e+06u area=4.347e+11p
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_0 A B VGND VPWR X VNB VPB
X0 VGND A a_68_355# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_150_355# B a_68_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_68_355# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_68_355# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_150_355# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_68_355# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_2 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_2 A B VGND VPWR Y VNB VPB
X0 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__macro_sparecell VNB LO VPB VGND VPWR
Xsky130_fd_sc_hd__nand2_2_1 LO LO VGND VPWR sky130_fd_sc_hd__nor2_2_1/B VNB VPB sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__nand2_2_0 LO LO VGND VPWR sky130_fd_sc_hd__nor2_2_0/B VNB VPB sky130_fd_sc_hd__nand2_2
Xsky130_fd_sc_hd__inv_2_0 sky130_fd_sc_hd__inv_2_0/A VGND VPWR sky130_fd_sc_hd__inv_2_0/Y
+ VNB VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__inv_2_1 sky130_fd_sc_hd__inv_2_1/A VGND VPWR sky130_fd_sc_hd__inv_2_1/Y
+ VNB VPB sky130_fd_sc_hd__inv_2
Xsky130_fd_sc_hd__nor2_2_0 sky130_fd_sc_hd__nor2_2_0/B sky130_fd_sc_hd__nor2_2_0/B
+ VGND VPWR sky130_fd_sc_hd__inv_2_0/A VNB VPB sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__nor2_2_1 sky130_fd_sc_hd__nor2_2_1/B sky130_fd_sc_hd__nor2_2_1/B
+ VGND VPWR sky130_fd_sc_hd__inv_2_1/A VNB VPB sky130_fd_sc_hd__nor2_2
Xsky130_fd_sc_hd__conb_1_0 VGND VNB VPB VPWR sky130_fd_sc_hd__conb_1_0/HI LO sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_logic1 gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_4_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VPWR X VNB VPB
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_115_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A1 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A2 a_115_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_115_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VPWR X VNB VPB
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VPWR X VNB VPB
X0 a_109_53# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_215_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_53# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_373_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_215_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_215_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_215_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_301_53# a_109_53# a_215_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_215_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_373_53# B a_301_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_109_53# a_215_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 zero vssd1 vssd
X_062_ _106_/Q user_gpio_out vssd vccd _062_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_131_ _131_/CLK hold4/X _086_/A vssd vccd hold3/A vssd vccd sky130_fd_sc_hd__dfrtp_4
X_114_ _101__9/Y hold4/X _084_/X _085_/Y vssd vccd _114_/Q _114_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xoutput7 _116_/Q vssd vccd pad_gpio_ana_en vssd vccd sky130_fd_sc_hd__buf_16
Xoutput20 _134_/X vssd vccd resetn_out vssd vccd sky130_fd_sc_hd__buf_16
X_104__12 _100__8/A vssd vccd _104__12/Y vssd vccd sky130_fd_sc_hd__inv_2
X_130_ _130_/CLK hold9/X _086_/A vssd vccd hold4/A vssd vccd sky130_fd_sc_hd__dfrtp_4
X_094__2 _101__9/A vssd vccd _094__2/Y vssd vccd sky130_fd_sc_hd__inv_2
X_061_ user_gpio_oeb _060_/X _106_/Q vssd vccd _061_/X vssd vccd sky130_fd_sc_hd__mux2_4
X_113_ _100__8/Y hold9/X _082_/X _083_/Y vssd vccd _113_/Q _113_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xclkbuf_1_0__f_serial_load clkbuf_0_serial_load/X vssd vccd _100__8/A vssd vccd sky130_fd_sc_hd__clkbuf_16
X_059__14 _130_/CLK vssd vccd _132_/CLK vssd vccd sky130_fd_sc_hd__inv_2
Xoutput8 _118_/Q vssd vccd pad_gpio_ana_pol vssd vccd sky130_fd_sc_hd__buf_16
Xoutput10 _113_/Q vssd vccd pad_gpio_dm[0] vssd vccd sky130_fd_sc_hd__buf_16
Xoutput21 _132_/Q vssd vccd serial_data_out vssd vccd sky130_fd_sc_hd__buf_16
X_060_ _112_/Q _063_/C vssd vccd _060_/X vssd vccd sky130_fd_sc_hd__and2_0
X_112_ _099__7/Y hold6/X _080_/X _081_/Y vssd vccd _112_/Q _112_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xhold10 _127_/Q vssd vccd _128_/D vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xoutput9 _117_/Q vssd vccd pad_gpio_ana_sel vssd vccd sky130_fd_sc_hd__buf_16
Xoutput11 _114_/Q vssd vccd pad_gpio_dm[1] vssd vccd sky130_fd_sc_hd__buf_16
Xoutput22 _067_/X vssd vccd user_gpio_in vssd vccd sky130_fd_sc_hd__buf_16
X_111_ _098__6/Y hold8/X _078_/X _079_/Y vssd vccd _111_/Q _111_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xhold11 _126_/Q vssd vccd _127_/D vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xoutput12 _115_/Q vssd vccd pad_gpio_dm[2] vssd vccd sky130_fd_sc_hd__buf_16
XANTENNA__072__B gpio_defaults[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_fanout29_A _082_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_110_ _097__5/Y hold7/X _076_/X _077_/Y vssd vccd _110_/Q _110_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xhold12 _125_/Q vssd vccd _126_/D vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xoutput13 _107_/Q vssd vccd pad_gpio_holdover vssd vccd sky130_fd_sc_hd__buf_16
X_097__5 _101__9/A vssd vccd _097__5/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__080__B gpio_defaults[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__075__B gpio_defaults[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__083__B gpio_defaults[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xhold13 _124_/Q vssd vccd _125_/D vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__078__B gpio_defaults[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput14 _111_/Q vssd vccd pad_gpio_ib_mode_sel vssd vccd sky130_fd_sc_hd__buf_16
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__091__B gpio_defaults[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__086__B gpio_defaults[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput15 _110_/Q vssd vccd pad_gpio_inenb vssd vccd sky130_fd_sc_hd__buf_16
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__089__B gpio_defaults[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xconst_source vssd vssd vccd vccd one_buffer/A zero_buffer/A sky130_fd_sc_hd__conb_1
XANTENNA_fanout27_A _082_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput16 _066_/Y vssd vccd pad_gpio_out vssd vccd sky130_fd_sc_hd__buf_16
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput17 _061_/X vssd vccd pad_gpio_outenb vssd vccd sky130_fd_sc_hd__buf_16
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xfanout30 fanout31/X vssd vccd _082_/A vssd vccd sky130_fd_sc_hd__buf_2
X_079_ _088_/A gpio_defaults[4] vssd vccd _079_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
Xoutput18 _108_/Q vssd vccd pad_gpio_slow_sel vssd vccd sky130_fd_sc_hd__buf_16
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input4_A resetn vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xfanout31 input4/X vssd vccd fanout31/X vssd vccd sky130_fd_sc_hd__buf_2
X_100__8 _100__8/A vssd vccd _100__8/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__061__A0 user_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_078_ _088_/A gpio_defaults[4] vssd vccd _078_/X vssd vccd sky130_fd_sc_hd__or2_0
Xoutput19 _109_/Q vssd vccd pad_gpio_vtrip_sel vssd vccd sky130_fd_sc_hd__buf_16
X_103__11 _100__8/A vssd vccd _103__11/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_077_ _076_/A gpio_defaults[3] vssd vccd _077_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_129_ _131_/CLK hold2/X _074_/A vssd vccd hold9/A vssd vccd sky130_fd_sc_hd__dfrtp_4
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_093_ _092_/A gpio_defaults[7] vssd vccd _093_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_076_ _076_/A gpio_defaults[3] vssd vccd _076_/X vssd vccd sky130_fd_sc_hd__or2_0
Xinput1 mgmt_gpio_oeb vssd vccd _063_/C vssd vccd sky130_fd_sc_hd__buf_2
X_128_ _131_/CLK _128_/D _074_/A vssd vccd hold2/A vssd vccd sky130_fd_sc_hd__dfrtp_4
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xfanout23 _092_/A vssd vccd _088_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_input2_A mgmt_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_092_ _092_/A gpio_defaults[7] vssd vccd _092_/X vssd vccd sky130_fd_sc_hd__or2_0
Xinput2 mgmt_gpio_out vssd vccd input2/X vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_0_serial_load_A serial_load vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_075_ _074_/A gpio_defaults[9] vssd vccd _075_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_127_ _130_/CLK _127_/D _092_/A vssd vccd _127_/Q vssd vccd sky130_fd_sc_hd__dfrtp_4
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xfanout24 fanout31/X vssd vccd _092_/A vssd vccd sky130_fd_sc_hd__buf_2
X_095__3 _100__8/A vssd vccd _095__3/Y vssd vccd sky130_fd_sc_hd__inv_2
X_074_ _074_/A gpio_defaults[9] vssd vccd _074_/X vssd vccd sky130_fd_sc_hd__or2_0
X_091_ _088_/A gpio_defaults[6] vssd vccd _091_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
Xinput3 pad_gpio_in vssd vccd _133_/A vssd vccd sky130_fd_sc_hd__buf_2
X_126_ _130_/CLK _126_/D _088_/A vssd vccd _126_/Q vssd vccd sky130_fd_sc_hd__dfrtp_4
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_109_ _096__4/Y hold2/X _074_/X _075_/Y vssd vccd _109_/Q _109_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xfanout25 _080_/A vssd vccd _076_/A vssd vccd sky130_fd_sc_hd__buf_2
X_090_ _092_/A gpio_defaults[6] vssd vccd _090_/X vssd vccd sky130_fd_sc_hd__or2_0
Xinput4 resetn vssd vccd input4/X vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__062__B user_gpio_out vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_073_ _074_/A gpio_defaults[8] vssd vccd _073_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_125_ _130_/CLK _125_/D _088_/A vssd vccd _125_/Q vssd vccd sky130_fd_sc_hd__dfrtp_4
XANTENNA__070__B gpio_defaults[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_108_ _095__3/Y _128_/D _072_/X _073_/Y vssd vccd _108_/Q _108_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xfanout26 fanout31/X vssd vccd _080_/A vssd vccd sky130_fd_sc_hd__buf_2
X_072_ _074_/A gpio_defaults[8] vssd vccd _072_/X vssd vccd sky130_fd_sc_hd__or2_0
Xinput5 serial_data_in vssd vccd _119_/D vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__068__B gpio_defaults[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__073__B gpio_defaults[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_124_ _130_/CLK hold8/X _092_/A vssd vccd _124_/Q vssd vccd sky130_fd_sc_hd__dfrtp_4
X_107_ _094__2/Y hold5/X _070_/X _071_/Y vssd vccd _107_/Q _107_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xfanout27 _082_/A vssd vccd _074_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__076__B gpio_defaults[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__081__B gpio_defaults[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_071_ _076_/A gpio_defaults[2] vssd vccd _071_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
XANTENNA__084__B gpio_defaults[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_106_ _058__1/Y hold1/X _068_/X _069_/Y vssd vccd _106_/Q _106_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
X_123_ _131_/CLK hold7/X _092_/A vssd vccd hold8/A vssd vccd sky130_fd_sc_hd__dfrtp_4
X_098__6 _100__8/A vssd vccd _098__6/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__079__B gpio_defaults[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xfanout28 _082_/A vssd vccd _086_/A vssd vccd sky130_fd_sc_hd__buf_2
XANTENNA__087__B gpio_defaults[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__092__B gpio_defaults[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_070_ _076_/A gpio_defaults[2] vssd vccd _070_/X vssd vccd sky130_fd_sc_hd__or2_0
X_122_ _130_/CLK hold5/X _076_/A vssd vccd hold7/A vssd vccd sky130_fd_sc_hd__dfrtp_4
Xspare_cell vssd spare_cell/LO vccd vssd vccd sky130_fd_sc_hd__macro_sparecell
Xserial_clock_out_buffer _131_/CLK vssd vccd serial_clock_out vssd vccd sky130_fd_sc_hd__clkbuf_16
Xfanout29 _082_/A vssd vccd _134_/A vssd vccd sky130_fd_sc_hd__buf_2
X_121_ _130_/CLK hold6/X _076_/A vssd vccd hold5/A vssd vccd sky130_fd_sc_hd__dfrtp_4
X_120_ _130_/CLK hold1/X _076_/A vssd vccd hold6/A vssd vccd sky130_fd_sc_hd__dfrtp_4
X_102__10 _101__9/A vssd vccd _102__10/Y vssd vccd sky130_fd_sc_hd__inv_2
X_058__1 _101__9/A vssd vccd _058__1/Y vssd vccd sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd vccd hold1/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_serial_load serial_load vssd vccd clkbuf_0_serial_load/X vssd vccd sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f_serial_clock clkbuf_0_serial_clock/X vssd vccd _130_/CLK vssd vccd
+ sky130_fd_sc_hd__clkbuf_16
Xhold2 hold2/A vssd vccd hold2/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xgpio_logic_high _067_/A vccd1 vssd1 gpio_logic_high
Xone_buffer one_buffer/A vssd vccd one vssd vccd sky130_fd_sc_hd__buf_16
XPHY_40 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xhold3 hold3/A vssd vccd hold3/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
X_101__9 _101__9/A vssd vccd _101__9/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_30 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_fanout28_A _082_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd vccd hold4/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xhold5 hold5/A vssd vccd hold5/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_32 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_089_ _088_/A gpio_defaults[5] vssd vccd _089_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
Xhold6 hold6/A vssd vccd hold6/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
Xzero_buffer zero_buffer/A vssd vccd zero vssd vccd sky130_fd_sc_hd__buf_16
XANTENNA_input5_A serial_data_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xclkbuf_0_serial_clock serial_clock vssd vccd clkbuf_0_serial_clock/X vssd vccd sky130_fd_sc_hd__clkbuf_16
X_105__13 _100__8/A vssd vccd _105__13/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_088_ _088_/A gpio_defaults[5] vssd vccd _088_/X vssd vccd sky130_fd_sc_hd__or2_0
Xhold7 hold7/A vssd vccd hold7/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
X_096__4 _101__9/A vssd vccd _096__4/Y vssd vccd sky130_fd_sc_hd__inv_2
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_087_ _134_/A gpio_defaults[12] vssd vccd _087_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
Xclkbuf_1_1__f_serial_load clkbuf_0_serial_load/X vssd vccd _101__9/A vssd vccd sky130_fd_sc_hd__clkbuf_16
Xhold8 hold8/A vssd vccd hold8/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__071__B gpio_defaults[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__082__A _082_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__074__B gpio_defaults[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_086_ _086_/A gpio_defaults[12] vssd vccd _086_/X vssd vccd sky130_fd_sc_hd__or2_0
Xclkbuf_1_1__f_serial_clock clkbuf_0_serial_clock/X vssd vccd _131_/CLK vssd vccd
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__069__B gpio_defaults[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_069_ _086_/A gpio_defaults[0] vssd vccd _069_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
Xhold9 hold9/A vssd vccd hold9/X vssd vccd sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__082__B gpio_defaults[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__077__B gpio_defaults[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input3_A pad_gpio_in vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__085__B gpio_defaults[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__090__B gpio_defaults[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_085_ _086_/A gpio_defaults[11] vssd vccd _085_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_068_ _086_/A gpio_defaults[0] vssd vccd _068_/X vssd vccd sky130_fd_sc_hd__or2_0
XANTENNA__093__B gpio_defaults[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__088__B gpio_defaults[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_067_ _067_/A _133_/A vssd vccd _067_/X vssd vccd sky130_fd_sc_hd__and2_2
X_084_ _086_/A gpio_defaults[11] vssd vccd _084_/X vssd vccd sky130_fd_sc_hd__or2_0
X_099__7 _101__9/A vssd vccd _099__7/Y vssd vccd sky130_fd_sc_hd__inv_2
X_119_ _131_/CLK _119_/D _080_/A vssd vccd hold1/A vssd vccd sky130_fd_sc_hd__dfrtp_4
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_083_ _074_/A gpio_defaults[10] vssd vccd _083_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_066_ _064_/X _065_/Y _062_/Y vssd vccd _066_/Y vssd vccd sky130_fd_sc_hd__o21ai_4
X_118_ _105__13/Y _127_/D _092_/X _093_/Y vssd vccd _118_/Q _118_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input1_A mgmt_gpio_oeb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_065_ input2/X _064_/B _106_/Q vssd vccd _065_/Y vssd vccd sky130_fd_sc_hd__o21ai_2
X_082_ _082_/A gpio_defaults[10] vssd vccd _082_/X vssd vccd sky130_fd_sc_hd__or2_0
X_134_ _134_/A vssd vccd _134_/X vssd vccd sky130_fd_sc_hd__buf_2
Xserial_load_out_buffer _101__9/A vssd vccd serial_load_out vssd vccd sky130_fd_sc_hd__clkbuf_16
X_117_ _104__12/Y _126_/D _090_/X _091_/Y vssd vccd _117_/Q _117_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_081_ _080_/A gpio_defaults[1] vssd vccd _081_/Y vssd vccd sky130_fd_sc_hd__nand2b_2
X_064_ _113_/Q_N _064_/B vssd vccd _064_/X vssd vccd sky130_fd_sc_hd__and2b_2
X_133_ _133_/A vssd vccd _133_/X vssd vccd sky130_fd_sc_hd__buf_2
X_116_ _103__11/Y _125_/D _088_/X _089_/Y vssd vccd _116_/Q _116_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_0_serial_clock_A serial_clock vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_063_ _115_/Q _114_/Q _063_/C vssd vccd _064_/B vssd vccd sky130_fd_sc_hd__and3b_2
X_080_ _080_/A gpio_defaults[1] vssd vccd _080_/X vssd vccd sky130_fd_sc_hd__or2_0
X_132_ _132_/CLK hold3/A _134_/A vssd vccd _132_/Q vssd vccd sky130_fd_sc_hd__dfrtp_2
X_115_ _102__10/Y hold3/X _086_/X _087_/Y vssd vccd _115_/Q _115_/Q_N vssd vccd sky130_fd_sc_hd__dfbbn_2
Xoutput6 _133_/X vssd vccd mgmt_gpio_in vssd vccd sky130_fd_sc_hd__buf_16
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt gpio_defaults_block VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
+ VGND
Xgpio_default_value\[8\] VGND VGND VPWR VPWR gpio_default_value\[8\]/HI gpio_defaults[8]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[6\] VGND VGND VPWR VPWR gpio_default_value\[6\]/HI gpio_defaults[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[4\] VGND VGND VPWR VPWR gpio_default_value\[4\]/HI gpio_defaults[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[2\] VGND VGND VPWR VPWR gpio_default_value\[2\]/HI gpio_defaults[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xgpio_default_value\[12\] VGND VGND VPWR VPWR gpio_default_value\[12\]/HI gpio_defaults[12]
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[0\] VGND VGND VPWR VPWR gpio_default_value\[0\]/HI gpio_defaults[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[10\] VGND VGND VPWR VPWR gpio_defaults[10] gpio_default_value\[10\]/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[9\] VGND VGND VPWR VPWR gpio_default_value\[9\]/HI gpio_defaults[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xgpio_default_value\[7\] VGND VGND VPWR VPWR gpio_default_value\[7\]/HI gpio_defaults[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[5\] VGND VGND VPWR VPWR gpio_default_value\[5\]/HI gpio_defaults[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[3\] VGND VGND VPWR VPWR gpio_default_value\[3\]/HI gpio_defaults[3]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xgpio_default_value\[1\] VGND VGND VPWR VPWR gpio_defaults[1] gpio_default_value\[1\]/LO
+ sky130_fd_sc_hd__conb_1
Xgpio_default_value\[11\] VGND VGND VPWR VPWR gpio_default_value\[11\]/HI gpio_defaults[11]
+ sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VPWR Y VNB VPB
X0 a_27_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_560_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_297# a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_474_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A a_560_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_27_47# B a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_474_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_560_47# a_27_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_27_297# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_560_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 a_79_21# A1 a_348_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# C1 a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_299_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_585_297# B1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_348_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_1 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_470_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_384_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_384_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VPWR Z VNB VPB
X0 VPWR a_27_47# a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X1 a_204_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_215_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Z A a_215_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND TE a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_215_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X9 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_8 A TE_B VGND VPWR Z VNB VPB
X0 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X7 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X12 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X17 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X19 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X23 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X24 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X30 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_80_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_674_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_386_47# D1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_674_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_566_47# B1 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_566_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_566_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_458_47# C1 a_386_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR S a_591_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_591_369# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_306_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND S a_578_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_306_369# a_257_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_79_21# A0 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_288_47# a_257_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_257_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_578_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_257_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_80_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_80_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_386_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_80_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_80_199# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_386_297# B1 a_80_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_458_47# A1 a_80_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A1 a_386_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_458_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvn_4 A TE_B VGND VPWR Z VNB VPB
X0 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X4 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X6 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Z A a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR TE_B a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X10 a_204_309# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=940000u l=150000u
X11 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47# A Z VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_204_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR TE_B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Z A a_204_309# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND TE_B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_108_21# B1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_346_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_108_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_108_21# A3 a_430_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_430_297# A2 a_346_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_108_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_346_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_108_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR B1 a_108_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_108_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_346_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 a_27_47# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_373_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_182_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_182_47# B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_373_297# A2 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_110_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A1 a_182_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_301_47# B2 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_383_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_301_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_81_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_81_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_579_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_81_21# B1 a_301_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_579_297# A2 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_81_21# B2 a_383_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VPWR Y VNB VPB
X0 a_408_47# B a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_408_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y a_27_47# a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_218_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_218_47# B a_408_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VPWR X VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VPWR Y VNB VPB
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VPWR Y VNB VPB
X0 VGND C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_277_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_277_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_381_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_2 A B VGND VPWR X VNB VPB
X0 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_470_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_470_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_112_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_470_47# B X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_470_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_112_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR B a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_112_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_297# B a_112_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_112_47# a_470_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_470_297# a_112_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X B a_470_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_112_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VPWR Y VNB VPB
X0 Y a_61_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_217_297# a_61_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_479_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_217_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y a_61_47# a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_61_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2 a_637_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_61_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_479_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B1_N a_61_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_637_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A3 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_352_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_549_47# A1 a_21_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_21_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_21_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_665_47# A2 a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_299_297# B1 a_21_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_21_199# B2 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND A3 a_665_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_21_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_21_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_21_199# B1 a_352_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_294_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A2_N a_295_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR B1 a_665_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_581_47# a_295_369# a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_665_369# B2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND B2 a_581_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_295_369# A2_N a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_84_21# a_295_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_295_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_581_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__einvp_1 A TE VGND VPWR Z VNB VPB
X0 a_276_297# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Z A a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR TE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Z A a_276_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_204_47# TE VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND TE a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VPWR Y VNB VPB
X0 VGND A2 a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A1 a_114_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_114_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VPWR X VNB VPB
X0 VPWR a_193_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# a_27_413# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_193_413# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_193_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_141_47# B2 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_497_297# A2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_225_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR C1 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_237_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_38_47# B2 a_237_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_225_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_141_47# C1 a_38_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_225_47# B1 a_141_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_2 A B C VGND VPWR X VNB VPB
X0 VPWR a_29_311# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_29_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_29_311# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_184_53# B a_112_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR C a_29_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_29_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_53# A a_29_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_29_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_184_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VPWR X VNB VPB
X0 VGND B1_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND A2 a_478_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_478_47# a_27_93# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_478_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A1 a_574_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B1_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_574_297# A2 a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_174_21# a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_429_297# A2 a_345_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_345_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_345_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_629_297# B2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B1 a_629_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_79_21# B2 a_345_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_345_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_79_21# A3 a_429_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_345_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR A2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_277_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_79_21# B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_277_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_361_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_277_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# A1 a_361_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 A VGND VPWR Y VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_2 A B VGND VPWR X VNB VPB
X0 a_121_297# B a_39_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_39_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_39_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_39_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_39_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A a_121_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND A a_39_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_39_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VPWR Y VNB VPB
X0 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_471_47# B a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# C a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_277_47# B a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A a_471_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_471_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND D a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt digital_pll VPWR clockp[1] dco div[0] div[1] div[2] div[3] div[4] enable ext_trim[0]
+ ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14] ext_trim[15] ext_trim[16]
+ ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20] ext_trim[21] ext_trim[22]
+ ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3] ext_trim[4] ext_trim[5]
+ ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb clockp[0] VGND
X_294_ _397_/A _325_/A VGND VPWR _313_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
X_363_ _348_/X ext_trim[2] _398_/B _362_/Y VGND VPWR _363_/X VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_13_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_432_ _437_/A _433_/B VGND VPWR _432_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[1\].id.delayint0 ringosc.dstage\[1\].id.delayen1/Z VGND VPWR ringosc.dstage\[1\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_346_ _346_/A VGND VPWR _456_/D VGND VPWR sky130_fd_sc_hd__buf_2
X_415_ _376_/A _370_/A _468_/Q VGND VPWR _416_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_10_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_277_ _420_/B _302_/A VGND VPWR _278_/D VGND VPWR sky130_fd_sc_hd__nor2_2
X_329_ _463_/Q _291_/X _328_/Y VGND VPWR _463_/D VGND VPWR sky130_fd_sc_hd__o21a_2
Xringosc.dstage\[11\].id.delayen1 ringosc.dstage\[11\].id.delayen1/A _423_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_2_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__392__A2 ext_trim[13] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__383__A2 ext_trim[9] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[10\].id.delayenb0 ringosc.dstage\[10\].id.delayenb1/A _385_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delayenb0 ringosc.dstage\[9\].id.delayenb1/A _383_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_13_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_293_ _293_/A VGND VPWR _328_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_431_ _437_/A _433_/B VGND VPWR _431_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_362_ _397_/A _438_/A VGND VPWR _362_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XANTENNA__410__A1 _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_414_ _406_/B _359_/A _371_/Y _403_/B _413_/X VGND VPWR _414_/X VGND VPWR sky130_fd_sc_hd__o2111a_2
X_276_ _465_/Q VGND VPWR _302_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_345_ _455_/Q _456_/Q _345_/S VGND VPWR _346_/A VGND VPWR sky130_fd_sc_hd__mux2_2
X_259_ _288_/B _288_/C _258_/X VGND VPWR _259_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_328_ _463_/Q _328_/B VGND VPWR _328_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[9\].id.delayenb1 ringosc.dstage\[9\].id.delayenb1/A _421_/X VGND
+ VPWR ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[10\].id.delayenb1 ringosc.dstage\[10\].id.delayenb1/A _422_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_15_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_292_ _397_/A _325_/A _278_/Y _291_/X VGND VPWR _293_/A VGND VPWR sky130_fd_sc_hd__o31a_2
XFILLER_13_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_430_ _437_/A _433_/B VGND VPWR _430_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_361_ _367_/A dco VGND VPWR _398_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_3_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_344_ _344_/A VGND VPWR _457_/D VGND VPWR sky130_fd_sc_hd__buf_2
X_413_ _301_/Y _367_/Y _386_/Y _412_/X VGND VPWR _413_/X VGND VPWR sky130_fd_sc_hd__o211a_2
X_275_ _466_/Q VGND VPWR _420_/B VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA__410__A2 ext_trim[18] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[4\].id.delayen0 ringosc.dstage\[4\].id.delayen0/A _369_/X VGND VPWR
+ ringosc.dstage\[4\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_2_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_258_ div[1] _258_/B VGND VPWR _258_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_327_ _327_/A VGND VPWR _464_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_16_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[5\].id.delayenb0 ringosc.dstage\[5\].id.delayenb1/A _373_/X VGND
+ VPWR ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[9\].id.delaybuf0 ringosc.dstage\[8\].id.delayen0/Z VGND VPWR ringosc.dstage\[9\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[10\].id.delaybuf0 ringosc.dstage\[9\].id.delayen0/Z VGND VPWR ringosc.dstage\[10\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_291_ _285_/X _291_/B _291_/C VGND VPWR _291_/X VGND VPWR sky130_fd_sc_hd__and3b_2
X_360_ _352_/X ext_trim[1] _403_/A VGND VPWR _360_/X VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_9_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__244__A div[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_274_ _464_/Q _463_/Q VGND VPWR _324_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_412_ _420_/B _283_/B _381_/A _376_/Y VGND VPWR _412_/X VGND VPWR sky130_fd_sc_hd__o22a_2
X_343_ _456_/Q _457_/Q _345_/S VGND VPWR _344_/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[4\].id.delayen1 ringosc.dstage\[4\].id.delayen1/A _409_/X VGND VPWR
+ ringosc.dstage\[4\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_257_ div[0] _257_/B _257_/C VGND VPWR _288_/C VGND VPWR sky130_fd_sc_hd__nand3b_2
X_326_ _464_/Q _325_/X _328_/B VGND VPWR _327_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XANTENNA__252__A div[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__427__A _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_309_ _309_/A _309_/B VGND VPWR _309_/X VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_15_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[5\].id.delayenb1 ringosc.dstage\[5\].id.delayenb1/A _410_/X VGND
+ VPWR ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[9\].id.delaybuf1 ringosc.dstage\[9\].id.delayenb1/A VGND VPWR ringosc.dstage\[9\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xringosc.dstage\[10\].id.delaybuf1 ringosc.dstage\[10\].id.delayenb1/A VGND VPWR ringosc.dstage\[10\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__350__A ext_trim[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__422__A1 _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_290_ _266_/X _290_/B _290_/C _290_/D VGND VPWR _291_/C VGND VPWR sky130_fd_sc_hd__nand4b_2
XANTENNA__404__A1 _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_273_ _467_/Q VGND VPWR _376_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_342_ _342_/A _347_/B _342_/C VGND VPWR _458_/D VGND VPWR sky130_fd_sc_hd__nand3_2
X_411_ _379_/X ext_trim[19] _403_/A _403_/B VGND VPWR _411_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_325_ _325_/A _325_/B VGND VPWR _325_/X VGND VPWR sky130_fd_sc_hd__xor2_2
X_256_ _256_/A VGND VPWR _257_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_0_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_239_ _262_/A _239_/B VGND VPWR _240_/C VGND VPWR sky130_fd_sc_hd__nand2b_2
X_308_ _420_/A _325_/A VGND VPWR _309_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_20_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__348__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__258__A div[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__422__A2 ext_trim[23] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[5\].id.delaybuf0 ringosc.dstage\[4\].id.delayen0/Z VGND VPWR ringosc.dstage\[5\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA__404__A2 ext_trim[16] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_272_ _302_/B VGND VPWR _325_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_341_ _342_/C _340_/Y _347_/B VGND VPWR _459_/D VGND VPWR sky130_fd_sc_hd__a21boi_2
X_410_ _428_/A ext_trim[18] _398_/X VGND VPWR _410_/X VGND VPWR sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[1\].id.delayenb0 ringosc.dstage\[1\].id.delayenb1/A _360_/X VGND
+ VPWR ringosc.dstage\[1\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[8\].id.delayint0 ringosc.dstage\[8\].id.delayen1/Z VGND VPWR ringosc.dstage\[8\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_5_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__A div[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_324_ _324_/A _324_/B VGND VPWR _325_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_255_ _342_/A _473_/Q VGND VPWR _256_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_307_ _313_/A _316_/A _316_/B _398_/A _325_/A VGND VPWR _309_/A VGND VPWR sky130_fd_sc_hd__a32o_2
X_238_ _461_/Q _476_/Q VGND VPWR _239_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_20_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__361__B dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[1\].id.delayenb1 ringosc.dstage\[1\].id.delayenb1/A _396_/X VGND
+ VPWR ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[5\].id.delaybuf1 ringosc.dstage\[5\].id.delayenb1/A VGND VPWR ringosc.dstage\[5\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_271_ _260_/X _266_/X _267_/X _290_/C VGND VPWR _302_/B VGND VPWR sky130_fd_sc_hd__o31a_2
X_340_ _459_/Q _342_/A VGND VPWR _340_/Y VGND VPWR sky130_fd_sc_hd__xnor2_2
X_469_ _477_/CLK _469_/D _445_/Y VGND VPWR _469_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delayen0 ringosc.dstage\[1\].id.delayen0/A _360_/X VGND VPWR
+ ringosc.dstage\[1\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__389__A2 ext_trim[12] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_323_ _328_/B _322_/Y _465_/Q _291_/X VGND VPWR _465_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_2
XFILLER_13_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_254_ _342_/A _473_/Q VGND VPWR _257_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_306_ _401_/B VGND VPWR _398_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_237_ _461_/Q _476_/Q VGND VPWR _262_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XANTENNA__289__A1 div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_270_ div[4] _266_/B _268_/Y _269_/Y VGND VPWR _290_/C VGND VPWR sky130_fd_sc_hd__o211a_2
X_399_ _379_/X ext_trim[15] _397_/Y _398_/X VGND VPWR _399_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_468_ _477_/CLK _468_/D _444_/Y VGND VPWR _468_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[1\].id.delayen1 ringosc.dstage\[1\].id.delayen1/A _396_/X VGND VPWR
+ ringosc.dstage\[1\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_322_ _322_/A _322_/B VGND VPWR _322_/Y VGND VPWR sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[1\].id.delaybuf0 ringosc.dstage\[0\].id.delayen0/Z VGND VPWR ringosc.dstage\[1\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_253_ _258_/B _253_/B VGND VPWR _288_/B VGND VPWR sky130_fd_sc_hd__nand2b_2
Xringosc.dstage\[4\].id.delayint0 ringosc.dstage\[4\].id.delayen1/Z VGND VPWR ringosc.dstage\[4\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_236_ _251_/A _251_/B _247_/B _235_/X VGND VPWR _240_/B VGND VPWR sky130_fd_sc_hd__a211o_2
X_305_ _301_/Y _322_/A _322_/B _406_/C _325_/A VGND VPWR _316_/B VGND VPWR sky130_fd_sc_hd__a32o_2
X_219_ _461_/Q _476_/Q _345_/S VGND VPWR _220_/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[9\].id.delayen0 ringosc.dstage\[9\].id.delayen0/A _383_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_16_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_398_ _398_/A _398_/B VGND VPWR _398_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_467_ _477_/CLK _467_/D _442_/Y VGND VPWR _467_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_4_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[1\].id.delaybuf1 ringosc.dstage\[1\].id.delayenb1/A VGND VPWR ringosc.dstage\[1\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_321_ _420_/B _321_/B VGND VPWR _466_/D VGND VPWR sky130_fd_sc_hd__xnor2_2
X_252_ div[1] VGND VPWR _253_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_235_ _459_/Q _474_/Q VGND VPWR _235_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_304_ _302_/B _303_/Y _324_/B VGND VPWR _322_/B VGND VPWR sky130_fd_sc_hd__a21o_2
XFILLER_1_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_218_ _218_/A VGND VPWR _477_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_19_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[9\].id.delayen1 ringosc.dstage\[9\].id.delayen1/A _421_/X VGND VPWR
+ ringosc.dstage\[9\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__270__A1 div[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_466_ _477_/CLK _466_/D _441_/Y VGND VPWR _466_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_397_ _397_/A _397_/B VGND VPWR _397_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_251_ _251_/A _251_/B VGND VPWR _258_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_320_ _302_/A _322_/B _319_/X _293_/A VGND VPWR _321_/B VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_13_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_449_ _454_/A _451_/B VGND VPWR _449_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_234_ _460_/Q _475_/Q VGND VPWR _247_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_303_ _324_/A VGND VPWR _303_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[0\].id.delayint0 ringosc.dstage\[0\].id.delayen1/Z VGND VPWR ringosc.dstage\[0\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.iss.reseten0 ringosc.iss.const1/HI _433_/B VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_1
XANTENNA__470__D osc VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_217_ _462_/Q _477_/Q _347_/B VGND VPWR _218_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XANTENNA__419__A1 _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_114 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_396_ _379_/X ext_trim[14] _372_/X _395_/X VGND VPWR _396_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_465_ _477_/CLK _465_/D _440_/Y VGND VPWR _465_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[8\].id.delayenb0 ringosc.dstage\[8\].id.delayenb1/A _380_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_5_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_250_ _250_/A _250_/B VGND VPWR _250_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_379_ dco VGND VPWR _379_/X VGND VPWR sky130_fd_sc_hd__buf_2
X_448_ _454_/A _451_/B VGND VPWR _448_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_1_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_233_ _459_/Q _474_/Q VGND VPWR _251_/B VGND VPWR sky130_fd_sc_hd__xor2_2
X_302_ _302_/A _302_/B VGND VPWR _322_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_1_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_216_ _345_/S VGND VPWR _347_/B VGND VPWR sky130_fd_sc_hd__buf_2
XANTENNA__419__A2 ext_trim[21] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.iss.delayint0 ringosc.iss.delayen1/Z VGND VPWR ringosc.iss.delayen0/A VGND
+ VPWR sky130_fd_sc_hd__clkinv_1
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_464_ _477_/CLK _464_/D _439_/Y VGND VPWR _464_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_395_ _376_/B _395_/B _395_/C VGND VPWR _395_/X VGND VPWR sky130_fd_sc_hd__and3b_2
Xringosc.dstage\[8\].id.delayenb1 ringosc.dstage\[8\].id.delayenb1/A _419_/X VGND
+ VPWR ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_4_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_378_ _352_/X ext_trim[7] _377_/X VGND VPWR _378_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_447_ dco VGND VPWR _454_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_232_ _458_/Q _473_/Q VGND VPWR _251_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_301_ _406_/C _381_/A VGND VPWR _301_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_1_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__373__A2 ext_trim[5] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_215_ _215_/A VGND VPWR _345_/S VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[6\].id.delayen0 ringosc.dstage\[6\].id.delayen0/A _375_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__364__A2 ext_trim[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_394_ _420_/A _278_/D _420_/C VGND VPWR _395_/C VGND VPWR sky130_fd_sc_hd__o21ai_2
X_463_ _477_/CLK _463_/D _437_/Y VGND VPWR _463_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_377_ _406_/C _376_/Y _403_/A VGND VPWR _377_/X VGND VPWR sky130_fd_sc_hd__o21a_2
X_446_ _446_/A _451_/B VGND VPWR _446_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[4\].id.delayenb0 ringosc.dstage\[4\].id.delayenb1/A _369_/X VGND
+ VPWR ringosc.dstage\[4\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[8\].id.delaybuf0 ringosc.dstage\[7\].id.delayen0/Z VGND VPWR ringosc.dstage\[8\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_231_ _460_/Q _231_/B VGND VPWR _240_/A VGND VPWR sky130_fd_sc_hd__nand2b_2
X_300_ _370_/A _465_/Q VGND VPWR _381_/A VGND VPWR sky130_fd_sc_hd__nand2_2
X_429_ _438_/A VGND VPWR _437_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[10\].id.delayen0 ringosc.dstage\[10\].id.delayen0/A _385_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_10_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_214_ _472_/D _472_/Q VGND VPWR _215_/A VGND VPWR sky130_fd_sc_hd__xnor2_2
Xringosc.dstage\[6\].id.delayen1 ringosc.dstage\[6\].id.delayen1/A _411_/X VGND VPWR
+ ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_393_ _468_/Q _406_/C _376_/A _367_/A VGND VPWR _395_/B VGND VPWR sky130_fd_sc_hd__a211o_2
X_462_ _477_/CLK _462_/D _436_/Y VGND VPWR _462_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[4\].id.delayenb1 ringosc.dstage\[4\].id.delayenb1/A _409_/X VGND
+ VPWR ringosc.dstage\[4\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[8\].id.delaybuf1 ringosc.dstage\[8\].id.delayenb1/A VGND VPWR ringosc.dstage\[8\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_376_ _376_/A _376_/B VGND VPWR _376_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_445_ _446_/A _451_/B VGND VPWR _445_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_230_ _475_/Q VGND VPWR _231_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_359_ _359_/A _359_/B VGND VPWR _403_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_428_ _428_/A _433_/B VGND VPWR _428_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[10\].id.delayen1 ringosc.dstage\[10\].id.delayen1/A _422_/X VGND
+ VPWR ringosc.dstage\[10\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_19_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__421__B1 ext_trim[22] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_392_ _428_/A ext_trim[13] _391_/X VGND VPWR _392_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_461_ _477_/CLK _461_/D _435_/Y VGND VPWR _461_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_4_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_375_ _352_/X ext_trim[6] _374_/Y VGND VPWR _375_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_444_ _446_/A _451_/B VGND VPWR _444_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_427_ _428_/A _433_/B VGND VPWR _427_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_358_ dco _358_/B VGND VPWR _359_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_289_ div[3] _242_/Y _249_/X _250_/Y VGND VPWR _290_/D VGND VPWR sky130_fd_sc_hd__o211a_2
Xringosc.dstage\[4\].id.delaybuf0 ringosc.dstage\[3\].id.delayen0/Z VGND VPWR ringosc.dstage\[4\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[0\].id.delayenb0 ringosc.dstage\[0\].id.delayenb1/A _351_/Y VGND
+ VPWR ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delayint0 ringosc.dstage\[7\].id.delayen1/Z VGND VPWR ringosc.dstage\[7\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_10_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__267__A1 div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__425__A enable VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_391_ _370_/A _376_/Y _403_/A VGND VPWR _391_/X VGND VPWR sky130_fd_sc_hd__o21a_2
X_460_ _477_/CLK _460_/D _433_/Y VGND VPWR _460_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_374_ _420_/B _358_/B dco VGND VPWR _374_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
X_443_ _454_/B VGND VPWR _451_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_1_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_288_ _258_/X _288_/B _288_/C _288_/D VGND VPWR _290_/B VGND VPWR sky130_fd_sc_hd__and4b_2
X_426_ _454_/B VGND VPWR _433_/B VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[3\].id.delayen0 ringosc.dstage\[3\].id.delayen0/A _364_/X VGND VPWR
+ ringosc.dstage\[3\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_357_ _469_/Q _398_/A VGND VPWR _358_/B VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[0\].id.delayenb1 ringosc.dstage\[0\].id.delayenb1/A _392_/X VGND
+ VPWR ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[4\].id.delaybuf1 ringosc.dstage\[4\].id.delayenb1/A VGND VPWR ringosc.dstage\[4\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__428__A _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_409_ _405_/Y _407_/X _408_/X ext_trim[17] _348_/X VGND VPWR _409_/X VGND VPWR sky130_fd_sc_hd__a32o_2
Xringosc.iss.delayenb0 ringosc.iss.delayenb1/A ringosc.iss.ctrlen0/X VGND VPWR ringosc.ibufp00/A
+ VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_21_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__425__B resetb VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_ringosc.dstage\[0\].id.delaybuf0_A ringosc.ibufp00/A VGND VPWR VPWR VGND
+ sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_390_ _438_/A VGND VPWR _428_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_13_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_373_ _352_/X ext_trim[5] _372_/X VGND VPWR _373_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_442_ _446_/A _442_/B VGND VPWR _442_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_287_ _251_/A _256_/A div[0] VGND VPWR _288_/D VGND VPWR sky130_fd_sc_hd__o21ai_2
X_425_ enable resetb VGND VPWR _454_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_356_ _386_/B _371_/B VGND VPWR _359_/A VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[3\].id.delayen1 ringosc.dstage\[3\].id.delayen1/A _404_/X VGND VPWR
+ ringosc.dstage\[3\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_408_ _420_/B _365_/Y _401_/Y _406_/B _403_/B VGND VPWR _408_/X VGND VPWR sky130_fd_sc_hd__o221a_2
X_339_ _339_/A VGND VPWR _460_/D VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[0\].id.delaybuf0 ringosc.ibufp00/A VGND VPWR ringosc.dstage\[0\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.iss.delayenb1 ringosc.iss.delayenb1/A _424_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[3\].id.delayint0 ringosc.dstage\[3\].id.delayen1/Z VGND VPWR ringosc.dstage\[3\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XANTENNA__349__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_372_ _301_/Y _367_/Y _359_/B _371_/Y VGND VPWR _372_/X VGND VPWR sky130_fd_sc_hd__o211a_2
X_441_ _446_/A _442_/B VGND VPWR _441_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XANTENNA__447__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_286_ _215_/A _455_/Q _457_/Q _456_/Q VGND VPWR _291_/B VGND VPWR sky130_fd_sc_hd__and4b_2
X_355_ _367_/A _397_/A _467_/Q VGND VPWR _371_/B VGND VPWR sky130_fd_sc_hd__and3_2
X_424_ _379_/X ext_trim[25] _403_/X _407_/C VGND VPWR _424_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_19_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_338_ _347_/B _338_/B VGND VPWR _339_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_407_ _407_/A _407_/B _407_/C VGND VPWR _407_/X VGND VPWR sky130_fd_sc_hd__and3_2
X_269_ _462_/Q _477_/Q VGND VPWR _269_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[0\].id.delaybuf1 ringosc.dstage\[0\].id.delayenb1/A VGND VPWR ringosc.dstage\[0\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.iss.delaybuf0 ringosc.iss.delayenb1/A VGND VPWR ringosc.iss.delayen1/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_371_ _397_/B _371_/B VGND VPWR _371_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_440_ _446_/A _442_/B VGND VPWR _440_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_285_ _302_/B _285_/B _324_/A VGND VPWR _285_/X VGND VPWR sky130_fd_sc_hd__and3_2
X_354_ _467_/Q _376_/B VGND VPWR _386_/B VGND VPWR sky130_fd_sc_hd__and2b_2
X_423_ _379_/X ext_trim[24] _362_/Y _420_/A VGND VPWR _423_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_337_ _331_/B _335_/Y _342_/C VGND VPWR _338_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
X_406_ _401_/Y _406_/B _406_/C VGND VPWR _407_/C VGND VPWR sky130_fd_sc_hd__nand3b_2
X_268_ _268_/A _268_/B VGND VPWR _268_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XANTENNA__424__A2 ext_trim[25] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_8_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_370_ _370_/A _465_/Q VGND VPWR _397_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_422_ _428_/A ext_trim[23] _398_/B VGND VPWR _422_/X VGND VPWR sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[0\].id.delayen0 ringosc.dstage\[0\].id.delayen0/A _351_/Y VGND VPWR
+ ringosc.dstage\[0\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_353_ _469_/Q _397_/A VGND VPWR _376_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_284_ _464_/Q _463_/Q VGND VPWR _324_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_10_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_267_ div[3] _242_/Y _249_/X VGND VPWR _267_/X VGND VPWR sky130_fd_sc_hd__o21ba_2
X_405_ _420_/A _406_/B _420_/C VGND VPWR _405_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
Xringosc.dstage\[7\].id.delayenb0 ringosc.dstage\[7\].id.delayenb1/A _378_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_18_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_336_ _462_/Q _336_/B VGND VPWR _342_/C VGND VPWR sky130_fd_sc_hd__nand2_2
XANTENNA__379__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__409__B1 ext_trim[17] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__360__A2 ext_trim[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_319_ _465_/Q _324_/A _325_/A VGND VPWR _319_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_20_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__260__A1 div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_17_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_421_ _407_/X _408_/X _420_/Y ext_trim[22] _348_/X VGND VPWR _421_/X VGND VPWR sky130_fd_sc_hd__a32o_2
Xringosc.dstage\[0\].id.delayen1 ringosc.dstage\[0\].id.delayen1/A _392_/X VGND VPWR
+ ringosc.dstage\[0\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_352_ _438_/A VGND VPWR _352_/X VGND VPWR sky130_fd_sc_hd__buf_2
X_283_ _298_/A _283_/B VGND VPWR _285_/B VGND VPWR sky130_fd_sc_hd__nor2_2
X_266_ div[4] _266_/B VGND VPWR _266_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_335_ _459_/Q _342_/A _460_/Q VGND VPWR _335_/Y VGND VPWR sky130_fd_sc_hd__a21oi_2
X_404_ _428_/A ext_trim[16] _403_/X VGND VPWR _404_/X VGND VPWR sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[7\].id.delayenb1 ringosc.dstage\[7\].id.delayenb1/A _417_/X VGND
+ VPWR ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_11_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_249_ _243_/Y _242_/A _242_/B _250_/A _250_/B VGND VPWR _249_/X VGND VPWR sky130_fd_sc_hd__o32a_2
X_318_ _318_/A VGND VPWR _467_/D VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[8\].id.delayen0 ringosc.dstage\[8\].id.delayen0/A _380_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_11_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclockp_buffer_0 _477_/CLK VGND VPWR clockp[0] VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_8_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_ringosc.ibufp00_A ringosc.ibufp00/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_5_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_351_ _348_/X _285_/B _350_/Y VGND VPWR _351_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
X_420_ _420_/A _420_/B _420_/C VGND VPWR _420_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
X_282_ _367_/A _401_/B VGND VPWR _283_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_334_ _461_/Q _331_/B _333_/Y _347_/B VGND VPWR _461_/D VGND VPWR sky130_fd_sc_hd__o211a_2
X_403_ _403_/A _403_/B _407_/B VGND VPWR _403_/X VGND VPWR sky130_fd_sc_hd__and3_2
X_265_ _268_/A _268_/B VGND VPWR _266_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_11_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_248_ _248_/A _248_/B VGND VPWR _250_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
X_317_ _376_/A _316_/X _328_/B VGND VPWR _318_/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[3\].id.delayenb0 ringosc.dstage\[3\].id.delayenb1/A _364_/X VGND
+ VPWR ringosc.dstage\[3\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[7\].id.delaybuf0 ringosc.dstage\[6\].id.delayen0/Z VGND VPWR ringosc.dstage\[7\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[11\].id.delayint0 ringosc.dstage\[11\].id.delayen1/Z VGND VPWR ringosc.dstage\[11\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xclockp_buffer_1 ringosc.ibufp11/Y VGND VPWR clockp[1] VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xringosc.dstage\[8\].id.delayen1 ringosc.dstage\[8\].id.delayen1/A _419_/X VGND VPWR
+ ringosc.dstage\[8\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__384__A_N ext_trim[10] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_350_ ext_trim[0] _438_/A VGND VPWR _350_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_281_ _468_/Q _467_/Q VGND VPWR _401_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XANTENNA__257__A_N div[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_264_ _262_/Y _240_/A _240_/B _263_/X VGND VPWR _268_/B VGND VPWR sky130_fd_sc_hd__a31o_2
X_333_ _462_/Q _336_/B VGND VPWR _333_/Y VGND VPWR sky130_fd_sc_hd__nand2b_2
X_402_ _381_/A _376_/Y _401_/Y _406_/C VGND VPWR _407_/B VGND VPWR sky130_fd_sc_hd__o22a_2
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__363__A2 ext_trim[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_316_ _316_/A _316_/B VGND VPWR _316_/X VGND VPWR sky130_fd_sc_hd__xor2_2
XFILLER_14_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_247_ _247_/A _247_/B VGND VPWR _248_/B VGND VPWR sky130_fd_sc_hd__nor2_2
Xringosc.dstage\[3\].id.delayenb1 ringosc.dstage\[3\].id.delayenb1/A _404_/X VGND
+ VPWR ringosc.dstage\[3\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[7\].id.delaybuf1 ringosc.dstage\[7\].id.delayenb1/A VGND VPWR ringosc.dstage\[7\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_11_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_280_ _469_/Q VGND VPWR _367_/A VGND VPWR sky130_fd_sc_hd__inv_2
X_263_ _461_/Q _476_/Q VGND VPWR _263_/X VGND VPWR sky130_fd_sc_hd__and2_2
X_332_ _462_/Q _336_/B _347_/B VGND VPWR _462_/D VGND VPWR sky130_fd_sc_hd__o21a_2
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_401_ _469_/Q _401_/B VGND VPWR _401_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_315_ _315_/A VGND VPWR _468_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_14_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_246_ _460_/Q _475_/Q VGND VPWR _247_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_22_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_229_ _468_/Q VGND VPWR _397_/A VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[3\].id.delaybuf0 ringosc.dstage\[2\].id.delayen0/Z VGND VPWR ringosc.dstage\[3\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xringosc.dstage\[6\].id.delayint0 ringosc.dstage\[6\].id.delayen1/Z VGND VPWR ringosc.dstage\[6\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XFILLER_0_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_477_ _477_/CLK _477_/D _454_/Y VGND VPWR _477_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.ibufp10 ringosc.ibufp10/A VGND VPWR ringosc.ibufp11/A VGND VPWR sky130_fd_sc_hd__clkinv_2
X_331_ _461_/Q _331_/B VGND VPWR _336_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_400_ _376_/Y _406_/B VGND VPWR _403_/B VGND VPWR sky130_fd_sc_hd__nand2b_2
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_262_ _262_/A VGND VPWR _262_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_2_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_245_ _251_/A _251_/B _235_/X VGND VPWR _248_/A VGND VPWR sky130_fd_sc_hd__a21oi_2
X_314_ _468_/Q _313_/Y _328_/B VGND VPWR _315_/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xringosc.dstage\[5\].id.delayen0 ringosc.dstage\[5\].id.delayen0/A _373_/X VGND VPWR
+ ringosc.ibufp10/A VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_22_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_228_ _469_/Q VGND VPWR _420_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[3\].id.delaybuf1 ringosc.dstage\[3\].id.delayenb1/A VGND VPWR ringosc.dstage\[3\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_3_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__375__A2 ext_trim[6] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_476_ _477_/CLK _476_/D _453_/Y VGND VPWR _476_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.ibufp00 ringosc.ibufp00/A VGND VPWR ringosc.ibufp01/A VGND VPWR sky130_fd_sc_hd__clkinv_2
Xringosc.ibufp11 ringosc.ibufp11/A VGND VPWR ringosc.ibufp11/Y VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_14_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_261_ _462_/Q _477_/Q VGND VPWR _268_/A VGND VPWR sky130_fd_sc_hd__xor2_2
X_330_ _460_/Q _459_/Q _342_/A VGND VPWR _331_/B VGND VPWR sky130_fd_sc_hd__and3_2
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_459_ _477_/CLK _459_/D _432_/Y VGND VPWR _459_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_11_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_313_ _313_/A _313_/B VGND VPWR _313_/Y VGND VPWR sky130_fd_sc_hd__xnor2_2
X_244_ div[2] VGND VPWR _250_/A VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[5\].id.delayen1 ringosc.dstage\[5\].id.delayen1/A _410_/X VGND VPWR
+ ringosc.dstage\[5\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XFILLER_22_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_227_ _227_/A VGND VPWR _473_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__387__B1 ext_trim[11] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delayint0 ringosc.dstage\[2\].id.delayen1/Z VGND VPWR ringosc.dstage\[2\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.ibufp01 ringosc.ibufp01/A VGND VPWR _477_/CLK VGND VPWR sky130_fd_sc_hd__clkinv_8
XFILLER_14_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_475_ _477_/CLK _475_/D _452_/Y VGND VPWR _475_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_260_ div[3] _242_/Y _249_/X _250_/Y _259_/X VGND VPWR _260_/X VGND VPWR sky130_fd_sc_hd__o2111a_2
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__243__A div[3] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_389_ _352_/X ext_trim[12] _388_/X VGND VPWR _389_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_458_ _477_/CLK _458_/D _431_/Y VGND VPWR _458_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_312_ _316_/A _316_/B _297_/B VGND VPWR _313_/B VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_14_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_243_ div[3] VGND VPWR _243_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xringosc.dstage\[11\].id.delayenb0 ringosc.dstage\[11\].id.delayenb1/A _387_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvn_8
XFILLER_19_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_226_ _342_/A _473_/Q _345_/S VGND VPWR _227_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_6_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__411__A2 ext_trim[19] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_474_ _477_/CLK _474_/D _451_/Y VGND VPWR _474_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA__287__B1 div[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_388_ _370_/A _367_/Y _359_/B VGND VPWR _388_/X VGND VPWR sky130_fd_sc_hd__o21a_2
X_457_ _477_/CLK _457_/D _430_/Y VGND VPWR _457_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_311_ _420_/A _328_/B _309_/X _310_/Y VGND VPWR _469_/D VGND VPWR sky130_fd_sc_hd__o22a_2
X_242_ _242_/A _242_/B VGND VPWR _242_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_11_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_225_ _458_/Q VGND VPWR _342_/A VGND VPWR sky130_fd_sc_hd__buf_2
Xringosc.dstage\[11\].id.delayenb1 ringosc.dstage\[11\].id.delayenb1/A _423_/X VGND
+ VPWR ringosc.dstage\[11\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
XFILLER_17_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__396__A2 ext_trim[14] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__378__A2 ext_trim[7] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__369__A2 ext_trim[4] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_473_ _477_/CLK _473_/D _450_/Y VGND VPWR _473_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_387_ _367_/Y _359_/B _386_/Y ext_trim[11] _348_/X VGND VPWR _387_/X VGND VPWR sky130_fd_sc_hd__a32o_2
X_456_ _477_/CLK _456_/D _428_/Y VGND VPWR _456_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_310_ _309_/A _309_/B _328_/B VGND VPWR _310_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_14_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_241_ _240_/A _240_/B _240_/C VGND VPWR _242_/B VGND VPWR sky130_fd_sc_hd__a21oi_2
Xringosc.dstage\[2\].id.delayen0 ringosc.dstage\[2\].id.delayen0/A _363_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.iss.const1 VGND VGND VPWR VPWR ringosc.iss.const1/HI ringosc.iss.const1/LO
+ sky130_fd_sc_hd__conb_1
X_439_ _446_/A _442_/B VGND VPWR _439_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_224_ _224_/A VGND VPWR _474_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[6\].id.delayenb0 ringosc.dstage\[6\].id.delayenb1/A _375_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[11\].id.delaybuf0 ringosc.dstage\[10\].id.delayen0/Z VGND VPWR ringosc.dstage\[11\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_472_ _477_/CLK _472_/D _449_/Y VGND VPWR _472_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA__358__A dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_455_ _477_/CLK _455_/D _427_/Y VGND VPWR _455_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_17_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_386_ _406_/B _386_/B VGND VPWR _386_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XANTENNA__423__A2 ext_trim[24] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_240_ _240_/A _240_/B _240_/C VGND VPWR _242_/A VGND VPWR sky130_fd_sc_hd__and3_2
Xringosc.dstage\[2\].id.delayen1 ringosc.dstage\[2\].id.delayen1/A _399_/X VGND VPWR
+ ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
X_369_ _352_/X ext_trim[4] _407_/A VGND VPWR _369_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_438_ _438_/A VGND VPWR _446_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_223_ _459_/Q _474_/Q _345_/S VGND VPWR _224_/A VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_10_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xringosc.dstage\[6\].id.delayenb1 ringosc.dstage\[6\].id.delayenb1/A _411_/X VGND
+ VPWR ringosc.dstage\[6\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[11\].id.delaybuf1 ringosc.dstage\[11\].id.delayenb1/A VGND VPWR ringosc.dstage\[11\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_471_ _477_/CLK _471_/D _448_/Y VGND VPWR _472_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_385_ _348_/X _283_/B _278_/D _384_/Y VGND VPWR _385_/X VGND VPWR sky130_fd_sc_hd__o31a_2
Xringosc.iss.delayen0 ringosc.iss.delayen0/A _389_/X VGND VPWR ringosc.ibufp00/A VGND
+ VPWR sky130_fd_sc_hd__einvp_2
XFILLER_17_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_454_ _454_/A _454_/B VGND VPWR _454_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XANTENNA__417__B1 ext_trim[20] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_299_ _466_/Q VGND VPWR _370_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_368_ _370_/A _365_/Y _367_/Y _359_/B VGND VPWR _407_/A VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_3_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_437_ _437_/A _442_/B VGND VPWR _437_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_222_ _222_/A VGND VPWR _475_/D VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__399__A2 ext_trim[15] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.dstage\[2\].id.delayenb0 ringosc.dstage\[2\].id.delayenb1/A _363_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvn_8
Xringosc.dstage\[6\].id.delaybuf0 ringosc.ibufp10/A VGND VPWR ringosc.dstage\[6\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_14_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_470_ _477_/CLK osc _446_/Y VGND VPWR _471_/D VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xringosc.dstage\[9\].id.delayint0 ringosc.dstage\[9\].id.delayen1/Z VGND VPWR ringosc.dstage\[9\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
Xringosc.dstage\[10\].id.delayint0 ringosc.dstage\[10\].id.delayen1/Z VGND VPWR ringosc.dstage\[10\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_384_ ext_trim[10] _438_/A VGND VPWR _384_/Y VGND VPWR sky130_fd_sc_hd__nand2b_2
Xringosc.iss.delayen1 ringosc.iss.delayen1/A _424_/X VGND VPWR ringosc.iss.delayen1/Z
+ VGND VPWR sky130_fd_sc_hd__einvp_2
X_453_ _454_/A _454_/B VGND VPWR _453_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_298_ _298_/A VGND VPWR _406_/C VGND VPWR sky130_fd_sc_hd__buf_2
X_367_ _367_/A _420_/C VGND VPWR _367_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_436_ _437_/A _442_/B VGND VPWR _436_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_6_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_221_ _460_/Q _475_/Q _345_/S VGND VPWR _222_/A VGND VPWR sky130_fd_sc_hd__mux2_2
X_419_ _428_/A ext_trim[21] _418_/X VGND VPWR _419_/X VGND VPWR sky130_fd_sc_hd__a21o_2
Xringosc.dstage\[2\].id.delayenb1 ringosc.dstage\[2\].id.delayenb1/A _399_/X VGND
+ VPWR ringosc.dstage\[2\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvn_4
Xringosc.dstage\[6\].id.delaybuf1 ringosc.dstage\[6\].id.delayenb1/A VGND VPWR ringosc.dstage\[6\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_383_ _379_/X ext_trim[9] _372_/X _382_/X VGND VPWR _383_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_452_ _454_/A _454_/B VGND VPWR _452_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_366_ _397_/A _376_/A VGND VPWR _420_/C VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_9_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_435_ _437_/A _442_/B VGND VPWR _435_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_297_ _297_/A _297_/B VGND VPWR _316_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_3_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_220_ _220_/A VGND VPWR _476_/D VGND VPWR sky130_fd_sc_hd__buf_2
X_349_ dco VGND VPWR _438_/A VGND VPWR sky130_fd_sc_hd__buf_2
X_418_ _370_/A _302_/A _401_/Y _403_/X VGND VPWR _418_/X VGND VPWR sky130_fd_sc_hd__o31a_2
XFILLER_17_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xringosc.iss.ctrlen0 _433_/B _389_/X VGND VPWR ringosc.iss.ctrlen0/X VGND VPWR sky130_fd_sc_hd__or2_2
XFILLER_9_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__380__A2 ext_trim[8] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delaybuf0 ringosc.dstage\[1\].id.delayen0/Z VGND VPWR ringosc.dstage\[2\].id.delayenb1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_2
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_382_ _406_/C _365_/Y _367_/Y _406_/B VGND VPWR _382_/X VGND VPWR sky130_fd_sc_hd__o22a_2
Xringosc.dstage\[5\].id.delayint0 ringosc.dstage\[5\].id.delayen1/Z VGND VPWR ringosc.dstage\[5\].id.delayen0/A
+ VGND VPWR sky130_fd_sc_hd__clkinv_1
X_451_ _454_/A _451_/B VGND VPWR _451_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_14_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_296_ _467_/Q _302_/B VGND VPWR _297_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_434_ _454_/B VGND VPWR _442_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_22_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_365_ _386_/B VGND VPWR _365_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_348_ dco VGND VPWR _348_/X VGND VPWR sky130_fd_sc_hd__buf_2
X_417_ _374_/Y _414_/X _416_/Y ext_trim[20] _348_/X VGND VPWR _417_/X VGND VPWR sky130_fd_sc_hd__a32o_2
X_279_ _420_/B _302_/A VGND VPWR _298_/A VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[7\].id.delayen0 ringosc.dstage\[7\].id.delayen0/A _378_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen0/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__374__B1 dco VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xringosc.dstage\[2\].id.delaybuf1 ringosc.dstage\[2\].id.delayenb1/A VGND VPWR ringosc.dstage\[2\].id.delayen1/A
+ VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_381_ _381_/A VGND VPWR _406_/B VGND VPWR sky130_fd_sc_hd__buf_2
X_450_ _454_/A _451_/B VGND VPWR _450_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_22_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_433_ _437_/A _433_/B VGND VPWR _433_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_364_ _352_/X ext_trim[3] _359_/B VGND VPWR _364_/X VGND VPWR sky130_fd_sc_hd__a21o_2
X_295_ _376_/A _302_/B VGND VPWR _297_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_278_ _469_/Q _376_/A _324_/B _278_/D VGND VPWR _278_/Y VGND VPWR sky130_fd_sc_hd__nand4_2
X_347_ _455_/Q _347_/B VGND VPWR _455_/D VGND VPWR sky130_fd_sc_hd__nand2b_2
X_416_ _420_/A _416_/B VGND VPWR _416_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xringosc.dstage\[11\].id.delayen0 ringosc.dstage\[11\].id.delayen0/A _387_/X VGND
+ VPWR ringosc.iss.delayenb1/A VGND VPWR sky130_fd_sc_hd__einvp_2
Xringosc.dstage\[7\].id.delayen1 ringosc.dstage\[7\].id.delayen1/A _417_/X VGND VPWR
+ ringosc.dstage\[7\].id.delayen1/Z VGND VPWR sky130_fd_sc_hd__einvp_2
XANTENNA__392__A1 _428_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_380_ _379_/X ext_trim[8] _359_/B _371_/Y VGND VPWR _380_/X VGND VPWR sky130_fd_sc_hd__a22o_2
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_20um abstract view
.subckt sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__gpiov2_pad_wrapped abstract view
.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H
+ OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO
+ ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_1um abstract view
.subckt sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_10um abstract view
.subckt sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for constant_block abstract view
.subckt constant_block one vccd vssd zero
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_5um abstract view
.subckt sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__analog_pad abstract view
.subckt sky130_ef_io__analog_pad P_CORE VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO
+ VSWITCH VSSIO VDDA VCCD VCCHIB VSSIO_Q P_PAD
.ends

* Black-box entry subcircuit for sky130_ef_io__disconnect_vdda_slice_5um abstract view
.subckt sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__corner_pad abstract view
.subckt sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vddio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um abstract view
.subckt sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B
+ VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q VSWITCH VCCHIB
.ends

* Black-box entry subcircuit for sky130_ef_io__vdda_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__top_power_hvc abstract view
.subckt sky130_ef_io__top_power_hvc AMUXBUS_A AMUXBUS_B DRN_HVC P_CORE P_PAD SRC_BDY_HVC
+ VSSA VDDA VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped3_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped3_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q VCCD1 VSSD1
.ends

* Black-box entry subcircuit for sky130_ef_io__vssa_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_fd_io__top_xres4v2 abstract view
.subckt sky130_fd_io__top_xres4v2 PAD_A_ESD_H XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H
+ ENABLE_H PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H
+ VSSIO VSSA VSSD AMUXBUS_B AMUXBUS_A VDDIO_Q VDDIO VSWITCH VDDA VCCD VCCHIB VSSIO_Q
+ PAD
.ends

.subckt chip_io_alt clock clock_core por flash_clk flash_csb flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_ieb_core flash_io0_oeb_core flash_io1 flash_io1_di_core
+ flash_io1_do_core flash_io1_ieb_core flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core
+ gpio_mode0_core gpio_out_core gpio_outenb_core vccd_pad vdda_pad vddio_pad vddio_pad2
+ vssa_pad vssd_pad vssio_pad vssio_pad2 mprj_io[0] mprj_io_analog_en[0] mprj_io_analog_pol[0]
+ mprj_io_analog_sel[0] mprj_io_dm[0] mprj_io_dm[1] mprj_io_dm[2] mprj_io_holdover[0]
+ mprj_io_ib_mode_sel[0] mprj_io_inp_dis[0] mprj_io_oeb[0] mprj_io_out[0] mprj_io_slow_sel[0]
+ mprj_io_vtrip_sel[0] mprj_io_in[0] mprj_io_in_3v3[0] mprj_gpio_analog[3] mprj_gpio_noesd[3]
+ mprj_io[10] mprj_io_analog_en[10] mprj_io_analog_pol[10] mprj_io_analog_sel[10]
+ mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_ib_mode_sel[10]
+ mprj_io_inp_dis[10] mprj_io_oeb[10] mprj_io_out[10] mprj_io_slow_sel[10] mprj_io_vtrip_sel[10]
+ mprj_io_in[10] mprj_io_in_3v3[10] mprj_gpio_analog[4] mprj_gpio_noesd[4] mprj_io[11]
+ mprj_io_analog_en[11] mprj_io_analog_pol[11] mprj_io_analog_sel[11] mprj_io_dm[33]
+ mprj_io_dm[34] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_ib_mode_sel[11] mprj_io_inp_dis[11]
+ mprj_io_oeb[11] mprj_io_out[11] mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_in[11]
+ mprj_io_in_3v3[11] mprj_gpio_analog[5] mprj_gpio_noesd[5] mprj_io[12] mprj_io_analog_en[12]
+ mprj_io_analog_pol[12] mprj_io_analog_sel[12] mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38]
+ mprj_io_holdover[12] mprj_io_ib_mode_sel[12] mprj_io_inp_dis[12] mprj_io_oeb[12]
+ mprj_io_out[12] mprj_io_slow_sel[12] mprj_io_vtrip_sel[12] mprj_io_in[12] mprj_io_in_3v3[12]
+ mprj_gpio_analog[6] mprj_gpio_noesd[6] mprj_io[13] mprj_io_analog_en[13] mprj_io_analog_pol[13]
+ mprj_io_analog_sel[13] mprj_io_dm[39] mprj_io_dm[40] mprj_io_dm[41] mprj_io_holdover[13]
+ mprj_io_ib_mode_sel[13] mprj_io_inp_dis[13] mprj_io_oeb[13] mprj_io_out[13] mprj_io_slow_sel[13]
+ mprj_io_vtrip_sel[13] mprj_io_in[13] mprj_io_in_3v3[13] mprj_io[1] mprj_io_analog_en[1]
+ mprj_io_analog_pol[1] mprj_io_analog_sel[1] mprj_io_dm[3] mprj_io_dm[4] mprj_io_dm[5]
+ mprj_io_holdover[1] mprj_io_ib_mode_sel[1] mprj_io_inp_dis[1] mprj_io_oeb[1] mprj_io_out[1]
+ mprj_io_slow_sel[1] mprj_io_vtrip_sel[1] mprj_io_in[1] mprj_io_in_3v3[1] mprj_io[2]
+ mprj_io_analog_en[2] mprj_io_analog_pol[2] mprj_io_analog_sel[2] mprj_io_dm[6] mprj_io_dm[7]
+ mprj_io_dm[8] mprj_io_holdover[2] mprj_io_ib_mode_sel[2] mprj_io_inp_dis[2] mprj_io_oeb[2]
+ mprj_io_out[2] mprj_io_slow_sel[2] mprj_io_vtrip_sel[2] mprj_io_in[2] mprj_io_in_3v3[2]
+ mprj_io[3] mprj_io_analog_en[3] mprj_io_analog_pol[3] mprj_io_analog_sel[3] mprj_io_dm[10]
+ mprj_io_dm[11] mprj_io_dm[9] mprj_io_holdover[3] mprj_io_ib_mode_sel[3] mprj_io_inp_dis[3]
+ mprj_io_oeb[3] mprj_io_out[3] mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_in[3]
+ mprj_io_in_3v3[3] mprj_io[4] mprj_io_analog_en[4] mprj_io_analog_pol[4] mprj_io_analog_sel[4]
+ mprj_io_dm[12] mprj_io_dm[13] mprj_io_dm[14] mprj_io_holdover[4] mprj_io_ib_mode_sel[4]
+ mprj_io_inp_dis[4] mprj_io_oeb[4] mprj_io_out[4] mprj_io_slow_sel[4] mprj_io_vtrip_sel[4]
+ mprj_io_in[4] mprj_io_in_3v3[4] mprj_io[5] mprj_io_analog_en[5] mprj_io_analog_pol[5]
+ mprj_io_analog_sel[5] mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17] mprj_io_holdover[5]
+ mprj_io_ib_mode_sel[5] mprj_io_inp_dis[5] mprj_io_oeb[5] mprj_io_out[5] mprj_io_slow_sel[5]
+ mprj_io_vtrip_sel[5] mprj_io_in[5] mprj_io_in_3v3[5] mprj_io[6] mprj_io_analog_en[6]
+ mprj_io_analog_pol[6] mprj_io_analog_sel[6] mprj_io_dm[18] mprj_io_dm[19] mprj_io_dm[20]
+ mprj_io_holdover[6] mprj_io_ib_mode_sel[6] mprj_io_inp_dis[6] mprj_io_oeb[6] mprj_io_out[6]
+ mprj_io_slow_sel[6] mprj_io_vtrip_sel[6] mprj_io_in[6] mprj_io_in_3v3[6] mprj_gpio_analog[0]
+ mprj_gpio_noesd[0] mprj_io[7] mprj_io_analog_en[7] mprj_io_analog_pol[7] mprj_io_analog_sel[7]
+ mprj_io_dm[21] mprj_io_dm[22] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_ib_mode_sel[7]
+ mprj_io_inp_dis[7] mprj_io_oeb[7] mprj_io_out[7] mprj_io_slow_sel[7] mprj_io_vtrip_sel[7]
+ mprj_io_in[7] mprj_io_in_3v3[7] mprj_gpio_analog[1] mprj_gpio_noesd[1] mprj_io[8]
+ mprj_io_analog_en[8] mprj_io_analog_pol[8] mprj_io_analog_sel[8] mprj_io_dm[24]
+ mprj_io_dm[25] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_ib_mode_sel[8] mprj_io_inp_dis[8]
+ mprj_io_oeb[8] mprj_io_out[8] mprj_io_slow_sel[8] mprj_io_vtrip_sel[8] mprj_io_in[8]
+ mprj_io_in_3v3[8] mprj_gpio_analog[2] mprj_gpio_noesd[2] mprj_io[9] mprj_io_analog_en[9]
+ mprj_io_analog_pol[9] mprj_io_analog_sel[9] mprj_io_dm[27] mprj_io_dm[28] mprj_io_dm[29]
+ mprj_io_holdover[9] mprj_io_ib_mode_sel[9] mprj_io_inp_dis[9] mprj_io_oeb[9] mprj_io_out[9]
+ mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_in[9] mprj_io_in_3v3[9] mprj_gpio_analog[7]
+ mprj_gpio_noesd[7] mprj_io[25] mprj_io_analog_en[14] mprj_io_analog_pol[14] mprj_io_analog_sel[14]
+ mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_ib_mode_sel[14]
+ mprj_io_inp_dis[14] mprj_io_oeb[14] mprj_io_out[14] mprj_io_slow_sel[14] mprj_io_vtrip_sel[14]
+ mprj_io_in[14] mprj_io_in_3v3[14] mprj_gpio_analog[17] mprj_gpio_noesd[17] mprj_io[35]
+ mprj_io_analog_en[24] mprj_io_analog_pol[24] mprj_io_analog_sel[24] mprj_io_dm[72]
+ mprj_io_dm[73] mprj_io_dm[74] mprj_io_holdover[24] mprj_io_ib_mode_sel[24] mprj_io_inp_dis[24]
+ mprj_io_oeb[24] mprj_io_out[24] mprj_io_slow_sel[24] mprj_io_vtrip_sel[24] mprj_io_in[24]
+ mprj_io_in_3v3[24] mprj_io[36] mprj_io_analog_en[25] mprj_io_analog_pol[25] mprj_io_analog_sel[25]
+ mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77] mprj_io_holdover[25] mprj_io_ib_mode_sel[25]
+ mprj_io_inp_dis[25] mprj_io_oeb[25] mprj_io_out[25] mprj_io_slow_sel[25] mprj_io_vtrip_sel[25]
+ mprj_io_in[25] mprj_io_in_3v3[25] mprj_io[37] mprj_io_analog_en[26] mprj_io_analog_pol[26]
+ mprj_io_analog_sel[26] mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[80] mprj_io_holdover[26]
+ mprj_io_ib_mode_sel[26] mprj_io_inp_dis[26] mprj_io_oeb[26] mprj_io_out[26] mprj_io_slow_sel[26]
+ mprj_io_vtrip_sel[26] mprj_io_in[26] mprj_io_in_3v3[26] mprj_gpio_analog[8] mprj_gpio_noesd[8]
+ mprj_io[26] mprj_io_analog_en[15] mprj_io_analog_pol[15] mprj_io_analog_sel[15]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_holdover[15] mprj_io_ib_mode_sel[15]
+ mprj_io_inp_dis[15] mprj_io_oeb[15] mprj_io_out[15] mprj_io_slow_sel[15] mprj_io_vtrip_sel[15]
+ mprj_io_in[15] mprj_io_in_3v3[15] mprj_gpio_analog[9] mprj_gpio_noesd[9] mprj_io[27]
+ mprj_io_analog_en[16] mprj_io_analog_pol[16] mprj_io_analog_sel[16] mprj_io_dm[48]
+ mprj_io_dm[49] mprj_io_dm[50] mprj_io_holdover[16] mprj_io_ib_mode_sel[16] mprj_io_inp_dis[16]
+ mprj_io_oeb[16] mprj_io_out[16] mprj_io_slow_sel[16] mprj_io_vtrip_sel[16] mprj_io_in[16]
+ mprj_io_in_3v3[16] mprj_gpio_analog[10] mprj_gpio_noesd[10] mprj_io[28] mprj_io_analog_en[17]
+ mprj_io_analog_pol[17] mprj_io_analog_sel[17] mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53]
+ mprj_io_holdover[17] mprj_io_ib_mode_sel[17] mprj_io_inp_dis[17] mprj_io_oeb[17]
+ mprj_io_out[17] mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_in[17] mprj_io_in_3v3[17]
+ mprj_gpio_analog[11] mprj_gpio_noesd[11] mprj_io[29] mprj_io_analog_en[18] mprj_io_analog_pol[18]
+ mprj_io_analog_sel[18] mprj_io_dm[54] mprj_io_dm[55] mprj_io_dm[56] mprj_io_holdover[18]
+ mprj_io_ib_mode_sel[18] mprj_io_inp_dis[18] mprj_io_oeb[18] mprj_io_out[18] mprj_io_slow_sel[18]
+ mprj_io_vtrip_sel[18] mprj_io_in[18] mprj_io_in_3v3[18] mprj_gpio_analog[12] mprj_gpio_noesd[12]
+ mprj_io[30] mprj_io_analog_en[19] mprj_io_analog_pol[19] mprj_io_analog_sel[19]
+ mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_holdover[19] mprj_io_ib_mode_sel[19]
+ mprj_io_inp_dis[19] mprj_io_oeb[19] mprj_io_out[19] mprj_io_slow_sel[19] mprj_io_vtrip_sel[19]
+ mprj_io_in[19] mprj_io_in_3v3[19] mprj_gpio_analog[13] mprj_gpio_noesd[13] mprj_io[31]
+ mprj_io_analog_en[20] mprj_io_analog_pol[20] mprj_io_analog_sel[20] mprj_io_dm[60]
+ mprj_io_dm[61] mprj_io_dm[62] mprj_io_holdover[20] mprj_io_ib_mode_sel[20] mprj_io_inp_dis[20]
+ mprj_io_oeb[20] mprj_io_out[20] mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_in[20]
+ mprj_io_in_3v3[20] mprj_gpio_analog[14] mprj_gpio_noesd[14] mprj_io[32] mprj_io_analog_en[21]
+ mprj_io_analog_pol[21] mprj_io_analog_sel[21] mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65]
+ mprj_io_holdover[21] mprj_io_ib_mode_sel[21] mprj_io_inp_dis[21] mprj_io_oeb[21]
+ mprj_io_out[21] mprj_io_slow_sel[21] mprj_io_vtrip_sel[21] mprj_io_in[21] mprj_io_in_3v3[21]
+ mprj_gpio_analog[15] mprj_gpio_noesd[15] mprj_io[33] mprj_io_analog_en[22] mprj_io_analog_pol[22]
+ mprj_io_analog_sel[22] mprj_io_dm[66] mprj_io_dm[67] mprj_io_dm[68] mprj_io_holdover[22]
+ mprj_io_ib_mode_sel[22] mprj_io_inp_dis[22] mprj_io_oeb[22] mprj_io_out[22] mprj_io_slow_sel[22]
+ mprj_io_vtrip_sel[22] mprj_io_in[22] mprj_io_in_3v3[22] mprj_gpio_analog[16] mprj_gpio_noesd[16]
+ mprj_io[34] mprj_io_analog_en[23] mprj_io_analog_pol[23] mprj_io_analog_sel[23]
+ mprj_io_dm[69] mprj_io_dm[70] mprj_io_dm[71] mprj_io_holdover[23] mprj_io_ib_mode_sel[23]
+ mprj_io_inp_dis[23] mprj_io_oeb[23] mprj_io_out[23] mprj_io_slow_sel[23] mprj_io_vtrip_sel[23]
+ mprj_io_in[23] mprj_io_in_3v3[23] resetb resetb_core_h vdda mprj_analog[1] mprj_io[15]
+ mprj_analog[2] mprj_io[16] mprj_analog[3] mprj_io[17] mprj_analog[0] mprj_io[14]
+ mprj_clamp_high[0] mprj_io[18] vccd1_pad vdda1_pad vdda1_pad2 vssa1_pad vssa1_pad2
+ vccd1 vdda1 vssd1 vssd1_pad mprj_analog[7] mprj_io[21] mprj_analog[8] mprj_io[22]
+ mprj_analog[9] mprj_io[23] mprj_analog[10] mprj_io[24] mprj_analog[5] mprj_clamp_high[1]
+ mprj_clamp_low[1] mprj_io[19] mprj_io[20] vccd2_pad vdda2_pad vssa2_pad vccd2 vdda2
+ vssd2 vssd2_pad flash_csb_core flash_clk_oeb_core flash_clk_core flash_csb_oeb_core
+ mprj_io_one[0] mprj_io_one[1] mprj_io_one[2] mprj_io_one[3] mprj_io_one[4] mprj_io_one[5]
+ mprj_io_one[6] mprj_io_one[7] mprj_io_one[8] mprj_io_one[9] mprj_io_one[10] mprj_io_one[11]
+ mprj_io_one[12] mprj_io_one[13] mprj_io_one[14] mprj_io_one[15] mprj_io_one[16]
+ mprj_io_one[17] mprj_io_one[18] mprj_io_one[19] mprj_io_one[20] mprj_io_one[21]
+ mprj_io_one[22] mprj_io_one[23] mprj_io_one[24] mprj_io_one[25] mprj_io_one[26]
+ porb_h gpio_mode1_core vssa mprj_analog[6] mprj_clamp_low[0] mprj_clamp_high[2]
+ mprj_clamp_low[2] vssa2 vddio vssa1 vssd mprj_analog[4] vccd vssio
XFILLER_570 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xclock_pad clock_pad/IN_H clock_pad/PAD_A_NOESD_H clock_pad/PAD_A_ESD_0_H clock_pad/PAD_A_ESD_1_H
+ clock clock_pad/OUT clock_pad/OUT clock_pad/OE_N clock_pad/HLD_H_N clock_core por
+ clock_pad/OUT porb_h porb_h clock_pad/TIE_LO_ESD clock_pad/OE_N clock_pad/HLD_H_N
+ clock_pad/TIE_LO_ESD clock_pad/OUT clock_pad/OUT clock_pad/OUT clock_pad/OUT clock_pad/OUT
+ clock_pad/OE_N clock_pad/TIE_LO_ESD clock_pad/OUT clock_pad/OUT gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q
+ sky130_ef_io__gpiov2_pad_wrapped
XFILLER_581 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_592 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vccd_lvc_clamped_pad
Xmprj_pads.area2_io_pad\[7\] mprj_io_in_3v3[21] mprj_gpio_noesd[14] mprj_gpio_analog[14]
+ mprj_pads.area2_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[32] mprj_io_dm[65] mprj_io_dm[64]
+ mprj_io_dm[63] mprj_pads.area2_io_pad\[7\]/HLD_H_N mprj_io_in[21] mprj_io_inp_dis[21]
+ mprj_io_ib_mode_sel[21] porb_h porb_h mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD mprj_io_oeb[21]
+ mprj_pads.area2_io_pad\[7\]/HLD_H_N mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD mprj_io_slow_sel[21]
+ mprj_io_vtrip_sel[21] mprj_io_holdover[21] mprj_io_analog_en[21] mprj_io_analog_sel[21]
+ mprj_io_one[21] mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD mprj_io_analog_pol[21] mprj_io_out[21]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_2 flash_csb_pad/DM[2] vccd vssd flash_csb_pad/SLOW constant_block
XFILLER_229 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_218 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_785 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_774 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_763 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_752 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_741 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_analog_pad\[2\] mprj_analog[9] vssa2 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda2 vccd vccd gpio_pad/VSSIO_Q mprj_io[23]
+ sky130_ef_io__analog_pad
XFILLER_571 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_582 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_593 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[7\] mprj_io_in_3v3[7] mprj_gpio_noesd[0] mprj_gpio_analog[0]
+ mprj_pads.area1_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[7] mprj_io_dm[23] mprj_io_dm[22]
+ mprj_io_dm[21] mprj_pads.area1_io_pad\[7\]/HLD_H_N mprj_io_in[7] mprj_io_inp_dis[7]
+ mprj_io_ib_mode_sel[7] mprj_pads.area1_io_pad\[7\]/ENABLE_H mprj_pads.area1_io_pad\[7\]/ENABLE_H
+ mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD mprj_io_oeb[7] mprj_pads.area1_io_pad\[7\]/HLD_H_N
+ mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD mprj_io_slow_sel[7] mprj_io_vtrip_sel[7]
+ mprj_io_holdover[7] mprj_io_analog_en[7] mprj_io_analog_sel[7] mprj_io_one[7] mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD
+ mprj_io_analog_pol[7] mprj_io_out[7] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xconstant_block_3 flash_clk_pad/DM[2] vccd vssd flash_clk_pad/SLOW constant_block
XFILLER_219 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_786 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_775 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_764 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_753 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_742 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_731 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_720 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_572 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_561 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_583 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_594 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_380 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_391 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[11\] mprj_io_in_3v3[11] mprj_gpio_noesd[4] mprj_gpio_analog[4]
+ mprj_pads.area1_io_pad\[11\]/PAD_A_ESD_1_H mprj_io[11] mprj_io_dm[35] mprj_io_dm[34]
+ mprj_io_dm[33] mprj_pads.area1_io_pad\[11\]/HLD_H_N mprj_io_in[11] mprj_io_inp_dis[11]
+ mprj_io_ib_mode_sel[11] mprj_pads.area1_io_pad\[11\]/ENABLE_H mprj_pads.area1_io_pad\[11\]/ENABLE_H
+ mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD mprj_io_oeb[11] mprj_pads.area1_io_pad\[11\]/HLD_H_N
+ mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD mprj_io_slow_sel[11] mprj_io_vtrip_sel[11]
+ mprj_io_holdover[11] mprj_io_analog_en[11] mprj_io_analog_sel[11] mprj_io_one[11]
+ mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD mprj_io_analog_pol[11] mprj_io_out[11] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xconstant_block_4 constant_block_4/one vccd vssd flash_io0_pad/SLOW constant_block
XFILLER_776 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_765 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_754 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_743 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_732 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_710 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_573 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_562 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_551 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_584 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_595 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_370 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_381 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_392 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_17 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xconstant_block_5 constant_block_5/one vccd vssd flash_io1_pad/SLOW constant_block
Xmprj_pads.area2_io_pad\[5\] mprj_io_in_3v3[19] mprj_gpio_noesd[12] mprj_gpio_analog[12]
+ mprj_pads.area2_io_pad\[5\]/PAD_A_ESD_1_H mprj_io[30] mprj_io_dm[59] mprj_io_dm[58]
+ mprj_io_dm[57] mprj_pads.area2_io_pad\[5\]/HLD_H_N mprj_io_in[19] mprj_io_inp_dis[19]
+ mprj_io_ib_mode_sel[19] porb_h porb_h mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD mprj_io_oeb[19]
+ mprj_pads.area2_io_pad\[5\]/HLD_H_N mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD mprj_io_slow_sel[19]
+ mprj_io_vtrip_sel[19] mprj_io_holdover[19] mprj_io_analog_en[19] mprj_io_analog_sel[19]
+ mprj_io_one[19] mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD mprj_io_analog_pol[19] mprj_io_out[19]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_777 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_766 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_755 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_744 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_733 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_722 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_700 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_574 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_563 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_552 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_541 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_585 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_596 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_analog_pad\[0\] mprj_analog[7] vssa2 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda2 vccd vccd gpio_pad/VSSIO_Q mprj_io[21]
+ sky130_ef_io__analog_pad
XFILLER_360 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_382 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_393 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[5\] mprj_io_in_3v3[5] mprj_pads.area1_io_pad\[5\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_1_H
+ mprj_io[5] mprj_io_dm[17] mprj_io_dm[16] mprj_io_dm[15] mprj_pads.area1_io_pad\[5\]/HLD_H_N
+ mprj_io_in[5] mprj_io_inp_dis[5] mprj_io_ib_mode_sel[5] porb_h porb_h mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_oeb[5] mprj_pads.area1_io_pad\[5\]/HLD_H_N mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_slow_sel[5] mprj_io_vtrip_sel[5] mprj_io_holdover[5] mprj_io_analog_en[5]
+ mprj_io_analog_sel[5] mprj_io_one[5] mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD mprj_io_analog_pol[5]
+ mprj_io_out[5] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xdisconnect_vdda_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
Xconstant_block_6 constant_block_6/one vccd vssd gpio_pad/SLOW constant_block
XFILLER_734 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_723 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_712 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_701 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_767 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_756 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_745 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_575 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_564 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_553 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_542 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_531 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_586 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_597 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_350 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_383 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_394 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_180 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xdisconnect_vdda_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
XFILLER_779 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_757 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_746 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_735 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_724 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_713 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_576 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_565 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_554 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_543 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_532 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_521 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_587 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xuser2_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xmgmt_vddio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_351 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_362 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_384 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_395 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xdisconnect_vdda_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
Xmgmt_vssio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_769 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_747 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_736 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_725 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_714 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_703 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[3\] mprj_io_in_3v3[17] mprj_gpio_noesd[10] mprj_gpio_analog[10]
+ mprj_pads.area2_io_pad\[3\]/PAD_A_ESD_1_H mprj_io[28] mprj_io_dm[53] mprj_io_dm[52]
+ mprj_io_dm[51] mprj_pads.area2_io_pad\[3\]/HLD_H_N mprj_io_in[17] mprj_io_inp_dis[17]
+ mprj_io_ib_mode_sel[17] porb_h porb_h mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD mprj_io_oeb[17]
+ mprj_pads.area2_io_pad\[3\]/HLD_H_N mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD mprj_io_slow_sel[17]
+ mprj_io_vtrip_sel[17] mprj_io_holdover[17] mprj_io_analog_en[17] mprj_io_analog_sel[17]
+ mprj_io_one[17] mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD mprj_io_analog_pol[17] mprj_io_out[17]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_577 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_566 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_555 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_544 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_533 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_522 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_511 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_599 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_352 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_330 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_363 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_374 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_385 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_396 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xsky130_ef_io__com_bus_slice_5um_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_193 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_182 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_160 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xbus_tie_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[3\] mprj_io_in_3v3[3] mprj_pads.area1_io_pad\[3\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_1_H
+ mprj_io[3] mprj_io_dm[11] mprj_io_dm[10] mprj_io_dm[9] mprj_pads.area1_io_pad\[3\]/HLD_H_N
+ mprj_io_in[3] mprj_io_inp_dis[3] mprj_io_ib_mode_sel[3] porb_h porb_h mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_oeb[3] mprj_pads.area1_io_pad\[3\]/HLD_H_N mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_holdover[3] mprj_io_analog_en[3]
+ mprj_io_analog_sel[3] mprj_io_one[3] mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD mprj_io_analog_pol[3]
+ mprj_io_out[3] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_759 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_748 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_737 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_726 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_715 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_704 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_578 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_567 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_556 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_545 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_534 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_523 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_512 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_501 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_320 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_331 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_353 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_364 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_375 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_386 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xsky130_ef_io__com_bus_slice_5um_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_397 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_194 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_183 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_161 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_150 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xbus_tie_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_738 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_727 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_716 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_705 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
XFILLER_579 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_568 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_557 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_546 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_535 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_524 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_513 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_502 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xsky130_ef_io__com_bus_slice_5um_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_321 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_332 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_354 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_365 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_376 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_387 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_398 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_140 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_analog_pad_with_clamp\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B mprj_clamp_high[2]
+ mprj_analog[6] mprj_io[20] mprj_clamp_low[2] vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__top_power_hvc
XFILLER_195 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_184 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_162 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_151 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_70 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[11\] mprj_io_in_3v3[25] mprj_pads.area2_io_pad\[11\]/PAD_A_NOESD_H
+ mprj_pads.area2_io_pad\[11\]/PAD_A_ESD_0_H mprj_pads.area2_io_pad\[11\]/PAD_A_ESD_1_H
+ mprj_io[36] mprj_io_dm[77] mprj_io_dm[76] mprj_io_dm[75] mprj_pads.area2_io_pad\[11\]/HLD_H_N
+ mprj_io_in[25] mprj_io_inp_dis[25] mprj_io_ib_mode_sel[25] porb_h porb_h mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_oeb[25] mprj_pads.area2_io_pad\[11\]/HLD_H_N mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_slow_sel[25] mprj_io_vtrip_sel[25] mprj_io_holdover[25] mprj_io_analog_en[25]
+ mprj_io_analog_sel[25] mprj_io_one[25] mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD mprj_io_analog_pol[25]
+ mprj_io_out[25] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_728 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_717 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_706 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_558 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_547 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_536 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_525 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_514 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_503 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[1\] mprj_io_in_3v3[15] mprj_gpio_noesd[8] mprj_gpio_analog[8]
+ mprj_pads.area2_io_pad\[1\]/PAD_A_ESD_1_H mprj_io[26] mprj_io_dm[47] mprj_io_dm[46]
+ mprj_io_dm[45] mprj_pads.area2_io_pad\[1\]/HLD_H_N mprj_io_in[15] mprj_io_inp_dis[15]
+ mprj_io_ib_mode_sel[15] porb_h porb_h mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD mprj_io_oeb[15]
+ mprj_pads.area2_io_pad\[1\]/HLD_H_N mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD mprj_io_slow_sel[15]
+ mprj_io_vtrip_sel[15] mprj_io_holdover[15] mprj_io_analog_en[15] mprj_io_analog_sel[15]
+ mprj_io_one[15] mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD mprj_io_analog_pol[15] mprj_io_out[15]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xsky130_ef_io__com_bus_slice_5um_3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_322 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_333 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_355 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_366 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_377 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_388 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_399 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_141 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_130 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_196 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_185 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_163 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_152 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser1_analog_pad\[3\] mprj_analog[0] vssa1 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda1 vccd vccd gpio_pad/VSSIO_Q mprj_io[14]
+ sky130_ef_io__analog_pad
Xbus_tie_4 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_729 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_718 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_707 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[1\] mprj_io_in_3v3[1] mprj_pads.area1_io_pad\[1\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_1_H
+ mprj_io[1] mprj_io_dm[5] mprj_io_dm[4] mprj_io_dm[3] mprj_pads.area1_io_pad\[1\]/HLD_H_N
+ mprj_io_in[1] mprj_io_inp_dis[1] mprj_io_ib_mode_sel[1] porb_h porb_h mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_oeb[1] mprj_pads.area1_io_pad\[1\]/HLD_H_N mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_slow_sel[1] mprj_io_vtrip_sel[1] mprj_io_holdover[1] mprj_io_analog_en[1]
+ mprj_io_analog_sel[1] mprj_io_one[1] mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD mprj_io_analog_pol[1]
+ mprj_io_out[1] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_559 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_548 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_537 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_526 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_515 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_504 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_301 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_312 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_356 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_367 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_378 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_389 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_142 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_131 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_120 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser1_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd1 vssd1 sky130_ef_io__vssd_lvc_clamped3_pad
XFILLER_197 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_186 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xgpio_pad gpio_pad/IN_H gpio_pad/PAD_A_NOESD_H gpio_pad/PAD_A_ESD_0_H gpio_pad/PAD_A_ESD_1_H
+ gpio gpio_mode1_core gpio_mode1_core gpio_mode0_core gpio_pad/HLD_H_N gpio_in_core
+ gpio_inenb_core gpio_pad/SLOW porb_h porb_h gpio_pad/TIE_LO_ESD gpio_outenb_core
+ gpio_pad/HLD_H_N gpio_pad/TIE_LO_ESD gpio_pad/SLOW gpio_pad/SLOW gpio_pad/SLOW gpio_pad/SLOW
+ gpio_pad/SLOW constant_block_6/one gpio_pad/TIE_LO_ESD gpio_pad/SLOW gpio_out_core
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_719 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_708 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_516 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_505 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_549 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_538 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_527 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_302 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_313 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_335 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_346 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_357 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_368 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_379 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_143 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_132 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_121 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_110 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_176 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_165 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vdda_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xbus_tie_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_40 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_709 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssd_lvc_clamped_pad
XFILLER_539 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_528 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_517 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_506 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_303 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_314 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_336 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_347 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_358 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_369 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_144 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_133 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_111 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_100 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_199 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_177 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_166 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser2_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd2 vssd2 sky130_ef_io__vccd_lvc_clamped3_pad
Xbus_tie_30 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xuser1_analog_pad\[1\] mprj_analog[2] vssa1 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda1 vccd vccd gpio_pad/VSSIO_Q mprj_io[16]
+ sky130_ef_io__analog_pad
Xbus_tie_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_529 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_518 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_507 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_304 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_315 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_337 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_348 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_359 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmgmt_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
XFILLER_145 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_123 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_112 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_101 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_178 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_167 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_SB1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_690 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_corner\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xuser1_vssa_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xbus_tie_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_519 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_508 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xsky130_ef_io__com_bus_slice_10um_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_305 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_316 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_338 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_349 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_146 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_135 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_124 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_113 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_102 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_SB2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_691 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_680 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_179 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_168 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_43 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_509 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xsky130_ef_io__com_bus_slice_10um_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_339 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_SB3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_147 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_136 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_125 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_114 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_103 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_169 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_681 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_670 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[8\] mprj_io_in_3v3[22] mprj_gpio_noesd[15] mprj_gpio_analog[15]
+ mprj_pads.area2_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[33] mprj_io_dm[68] mprj_io_dm[67]
+ mprj_io_dm[66] mprj_pads.area2_io_pad\[8\]/HLD_H_N mprj_io_in[22] mprj_io_inp_dis[22]
+ mprj_io_ib_mode_sel[22] porb_h porb_h mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD mprj_io_oeb[22]
+ mprj_pads.area2_io_pad\[8\]/HLD_H_N mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD mprj_io_slow_sel[22]
+ mprj_io_vtrip_sel[22] mprj_io_holdover[22] mprj_io_analog_en[22] mprj_io_analog_sel[22]
+ mprj_io_one[22] mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD mprj_io_analog_pol[22] mprj_io_out[22]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_318 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_329 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_137 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_126 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_115 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_104 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_analog_pad\[3\] mprj_analog[10] vssa2 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda2 vccd vccd gpio_pad/VSSIO_Q mprj_io[24]
+ sky130_ef_io__analog_pad
XFILLER_159 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_148 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_693 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_682 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_671 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_660 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_56 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_67 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[8\] mprj_io_in_3v3[8] mprj_gpio_noesd[1] mprj_gpio_analog[1]
+ mprj_pads.area1_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[8] mprj_io_dm[26] mprj_io_dm[25]
+ mprj_io_dm[24] mprj_pads.area1_io_pad\[8\]/HLD_H_N mprj_io_in[8] mprj_io_inp_dis[8]
+ mprj_io_ib_mode_sel[8] mprj_pads.area1_io_pad\[8\]/ENABLE_H mprj_pads.area1_io_pad\[8\]/ENABLE_H
+ mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD mprj_io_oeb[8] mprj_pads.area1_io_pad\[8\]/HLD_H_N
+ mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD mprj_io_slow_sel[8] mprj_io_vtrip_sel[8]
+ mprj_io_holdover[8] mprj_io_analog_en[8] mprj_io_analog_sel[8] mprj_io_one[8] mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD
+ mprj_io_analog_pol[8] mprj_io_out[8] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xresetb_pad xresloop resetb_core_h xres_vss_loop constant_block_0/one xresloop porb_h
+ xres_vss_loop xres_vss_loop xres_vss_loop resetb_pad/TIE_HI_ESD xres_vss_loop xres_vss_loop
+ vssio vssa vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A gpio_pad/VDDIO_Q vddio vddio
+ vdda vccd vccd gpio_pad/VSSIO_Q resetb sky130_fd_io__top_xres4v2
XFILLER_319 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_138 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_127 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_116 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_105 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_149 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_694 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_672 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_661 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_650 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_491 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[12\] mprj_io_in_3v3[12] mprj_gpio_noesd[5] mprj_gpio_analog[5]
+ mprj_pads.area1_io_pad\[12\]/PAD_A_ESD_1_H mprj_io[12] mprj_io_dm[38] mprj_io_dm[37]
+ mprj_io_dm[36] mprj_pads.area1_io_pad\[12\]/HLD_H_N mprj_io_in[12] mprj_io_inp_dis[12]
+ mprj_io_ib_mode_sel[12] mprj_pads.area1_io_pad\[12\]/ENABLE_H mprj_pads.area1_io_pad\[12\]/ENABLE_H
+ mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD mprj_io_oeb[12] mprj_pads.area1_io_pad\[12\]/HLD_H_N
+ mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD mprj_io_slow_sel[12] mprj_io_vtrip_sel[12]
+ mprj_io_holdover[12] mprj_io_analog_en[12] mprj_io_analog_sel[12] mprj_io_one[12]
+ mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD mprj_io_analog_pol[12] mprj_io_out[12] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_139 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_128 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_117 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_106 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_695 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_684 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_673 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_662 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_640 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_651 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_492 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_481 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_58 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[6\] mprj_io_in_3v3[20] mprj_gpio_noesd[13] mprj_gpio_analog[13]
+ mprj_pads.area2_io_pad\[6\]/PAD_A_ESD_1_H mprj_io[31] mprj_io_dm[62] mprj_io_dm[61]
+ mprj_io_dm[60] mprj_pads.area2_io_pad\[6\]/HLD_H_N mprj_io_in[20] mprj_io_inp_dis[20]
+ mprj_io_ib_mode_sel[20] porb_h porb_h mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD mprj_io_oeb[20]
+ mprj_pads.area2_io_pad\[6\]/HLD_H_N mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD mprj_io_slow_sel[20]
+ mprj_io_vtrip_sel[20] mprj_io_holdover[20] mprj_io_analog_en[20] mprj_io_analog_sel[20]
+ mprj_io_one[20] mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD mprj_io_analog_pol[20] mprj_io_out[20]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xflash_csb_pad flash_csb_pad/IN_H flash_csb_pad/PAD_A_NOESD_H flash_csb_pad/PAD_A_ESD_0_H
+ flash_csb_pad/PAD_A_ESD_1_H flash_csb flash_csb_pad/DM[2] flash_csb_pad/DM[2] flash_csb_pad/SLOW
+ flash_csb_pad/HLD_H_N flash_csb_pad/IN flash_csb_pad/SLOW flash_csb_pad/SLOW porb_h
+ porb_h flash_csb_pad/TIE_LO_ESD flash_csb_oeb_core flash_csb_pad/HLD_H_N flash_csb_pad/TIE_LO_ESD
+ flash_csb_pad/SLOW flash_csb_pad/SLOW flash_csb_pad/SLOW flash_csb_pad/SLOW flash_csb_pad/SLOW
+ flash_csb_pad/DM[2] flash_csb_pad/TIE_LO_ESD flash_csb_pad/SLOW flash_csb_core gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q
+ sky130_ef_io__gpiov2_pad_wrapped
XFILLER_129 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_118 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_107 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_696 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_685 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_663 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_630 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_641 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_652 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_analog_pad\[1\] mprj_analog[8] vssa2 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda2 vccd vccd gpio_pad/VSSIO_Q mprj_io[22]
+ sky130_ef_io__analog_pad
XFILLER_493 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_482 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_471 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_48 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_59 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[6\] mprj_io_in_3v3[6] mprj_pads.area1_io_pad\[6\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_1_H
+ mprj_io[6] mprj_io_dm[20] mprj_io_dm[19] mprj_io_dm[18] mprj_pads.area1_io_pad\[6\]/HLD_H_N
+ mprj_io_in[6] mprj_io_inp_dis[6] mprj_io_ib_mode_sel[6] porb_h porb_h mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_oeb[6] mprj_pads.area1_io_pad\[6\]/HLD_H_N mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_slow_sel[6] mprj_io_vtrip_sel[6] mprj_io_holdover[6] mprj_io_analog_en[6]
+ mprj_io_analog_sel[6] mprj_io_one[6] mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD mprj_io_analog_pol[6]
+ mprj_io_out[6] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_119 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_108 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_697 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_686 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_675 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_620 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_631 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_642 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_653 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_494 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_483 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_472 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_461 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_16 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_280 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[10\] mprj_io_in_3v3[10] mprj_gpio_noesd[3] mprj_gpio_analog[3]
+ mprj_pads.area1_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[10] mprj_io_dm[32] mprj_io_dm[31]
+ mprj_io_dm[30] mprj_pads.area1_io_pad\[10\]/HLD_H_N mprj_io_in[10] mprj_io_inp_dis[10]
+ mprj_io_ib_mode_sel[10] mprj_pads.area1_io_pad\[10\]/ENABLE_H mprj_pads.area1_io_pad\[10\]/ENABLE_H
+ mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD mprj_io_oeb[10] mprj_pads.area1_io_pad\[10\]/HLD_H_N
+ mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD mprj_io_slow_sel[10] mprj_io_vtrip_sel[10]
+ mprj_io_holdover[10] mprj_io_analog_en[10] mprj_io_analog_sel[10] mprj_io_one[10]
+ mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD mprj_io_analog_pol[10] mprj_io_out[10] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xflash_io1_pad flash_io1_pad/IN_H flash_io1_pad/PAD_A_NOESD_H flash_io1_pad/PAD_A_ESD_0_H
+ flash_io1_pad/PAD_A_ESD_1_H flash_io1 flash_io1_ieb_core flash_io1_ieb_core flash_io1_oeb_core
+ flash_io1_pad/HLD_H_N flash_io1_di_core flash_io1_ieb_core flash_io1_pad/SLOW porb_h
+ porb_h flash_io1_pad/TIE_LO_ESD flash_io1_oeb_core flash_io1_pad/HLD_H_N flash_io1_pad/TIE_LO_ESD
+ flash_io1_pad/SLOW flash_io1_pad/SLOW flash_io1_pad/SLOW flash_io1_pad/SLOW flash_io1_pad/SLOW
+ constant_block_5/one flash_io1_pad/TIE_LO_ESD flash_io1_pad/SLOW flash_io1_do_core
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_698 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_687 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_676 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_665 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_610 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_621 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_632 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_643 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_654 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmgmt_vddio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_495 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_484 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_473 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_462 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_451 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_28 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_17 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_270 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_281 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[4\] mprj_io_in_3v3[18] mprj_gpio_noesd[11] mprj_gpio_analog[11]
+ mprj_pads.area2_io_pad\[4\]/PAD_A_ESD_1_H mprj_io[29] mprj_io_dm[56] mprj_io_dm[55]
+ mprj_io_dm[54] mprj_pads.area2_io_pad\[4\]/HLD_H_N mprj_io_in[18] mprj_io_inp_dis[18]
+ mprj_io_ib_mode_sel[18] porb_h porb_h mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD mprj_io_oeb[18]
+ mprj_pads.area2_io_pad\[4\]/HLD_H_N mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD mprj_io_slow_sel[18]
+ mprj_io_vtrip_sel[18] mprj_io_holdover[18] mprj_io_analog_en[18] mprj_io_analog_sel[18]
+ mprj_io_one[18] mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD mprj_io_analog_pol[18] mprj_io_out[18]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xuser1_analog_pad_with_clamp gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B mprj_clamp_high[0]
+ mprj_analog[4] mprj_io[18] mprj_clamp_low[0] vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__top_power_hvc
XFILLER_699 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_688 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_677 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_666 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_600 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_611 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_622 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_633 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_644 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_496 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_485 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_474 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_463 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_452 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_441 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_271 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_282 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[4\] mprj_io_in_3v3[4] mprj_pads.area1_io_pad\[4\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_1_H
+ mprj_io[4] mprj_io_dm[14] mprj_io_dm[13] mprj_io_dm[12] mprj_pads.area1_io_pad\[4\]/HLD_H_N
+ mprj_io_in[4] mprj_io_inp_dis[4] mprj_io_ib_mode_sel[4] porb_h porb_h mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_oeb[4] mprj_pads.area1_io_pad\[4\]/HLD_H_N mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_slow_sel[4] mprj_io_vtrip_sel[4] mprj_io_holdover[4] mprj_io_analog_en[4]
+ mprj_io_analog_sel[4] mprj_io_one[4] mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD mprj_io_analog_pol[4]
+ mprj_io_out[4] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_689 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_678 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_667 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_656 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_601 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_612 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_623 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_634 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_90 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_497 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_486 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_475 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_464 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_453 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_442 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_431 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_250 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_261 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_679 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_668 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_657 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_602 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_613 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_624 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_635 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_646 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_91 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_80 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_498 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_487 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_476 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_465 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_454 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_443 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_421 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_432 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_251 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_262 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_284 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_295 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vssd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd2 vssd2 sky130_ef_io__vssd_lvc_clamped3_pad
Xmprj_pads.area2_io_pad\[12\] mprj_io_in_3v3[26] mprj_pads.area2_io_pad\[12\]/PAD_A_NOESD_H
+ mprj_pads.area2_io_pad\[12\]/PAD_A_ESD_0_H mprj_pads.area2_io_pad\[12\]/PAD_A_ESD_1_H
+ mprj_io[37] mprj_io_dm[80] mprj_io_dm[79] mprj_io_dm[78] mprj_pads.area2_io_pad\[12\]/HLD_H_N
+ mprj_io_in[26] mprj_io_inp_dis[26] mprj_io_ib_mode_sel[26] porb_h porb_h mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_oeb[26] mprj_pads.area2_io_pad\[12\]/HLD_H_N mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_slow_sel[26] mprj_io_vtrip_sel[26] mprj_io_holdover[26] mprj_io_analog_en[26]
+ mprj_io_analog_sel[26] mprj_io_one[26] mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD mprj_io_analog_pol[26]
+ mprj_io_out[26] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vssio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_603 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_614 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_625 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_669 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_658 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_647 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_92 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_81 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_70 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[2\] mprj_io_in_3v3[16] mprj_gpio_noesd[9] mprj_gpio_analog[9]
+ mprj_pads.area2_io_pad\[2\]/PAD_A_ESD_1_H mprj_io[27] mprj_io_dm[50] mprj_io_dm[49]
+ mprj_io_dm[48] mprj_pads.area2_io_pad\[2\]/HLD_H_N mprj_io_in[16] mprj_io_inp_dis[16]
+ mprj_io_ib_mode_sel[16] porb_h porb_h mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD mprj_io_oeb[16]
+ mprj_pads.area2_io_pad\[2\]/HLD_H_N mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD mprj_io_slow_sel[16]
+ mprj_io_vtrip_sel[16] mprj_io_holdover[16] mprj_io_analog_en[16] mprj_io_analog_sel[16]
+ mprj_io_one[16] mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD mprj_io_analog_pol[16] mprj_io_out[16]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_499 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_488 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_477 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_466 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_455 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_444 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_411 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_422 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_433 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_230 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_252 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_263 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_285 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_296 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser2_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[2\] mprj_io_in_3v3[2] mprj_pads.area1_io_pad\[2\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_1_H
+ mprj_io[2] mprj_io_dm[8] mprj_io_dm[7] mprj_io_dm[6] mprj_pads.area1_io_pad\[2\]/HLD_H_N
+ mprj_io_in[2] mprj_io_inp_dis[2] mprj_io_ib_mode_sel[2] porb_h porb_h mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_oeb[2] mprj_pads.area1_io_pad\[2\]/HLD_H_N mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_slow_sel[2] mprj_io_vtrip_sel[2] mprj_io_holdover[2] mprj_io_analog_en[2]
+ mprj_io_analog_sel[2] mprj_io_one[2] mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD mprj_io_analog_pol[2]
+ mprj_io_out[2] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_659 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_604 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_615 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_626 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_637 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_648 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_93 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_82 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_489 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_478 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_467 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_456 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_445 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_401 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_412 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_423 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_434 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_231 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_220 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_253 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_264 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_286 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_297 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_605 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_616 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_638 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_649 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_94 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_83 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_479 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_468 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_457 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_446 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_435 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_402 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_413 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_424 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_210 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_254 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_265 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_287 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_298 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser2_analog_pad_with_clamp\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B mprj_clamp_high[1]
+ mprj_analog[5] mprj_io[19] mprj_clamp_low[1] vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__top_power_hvc
Xuser1_vdda_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[10\] mprj_io_in_3v3[24] mprj_gpio_noesd[17] mprj_gpio_analog[17]
+ mprj_pads.area2_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[35] mprj_io_dm[74] mprj_io_dm[73]
+ mprj_io_dm[72] mprj_pads.area2_io_pad\[10\]/HLD_H_N mprj_io_in[24] mprj_io_inp_dis[24]
+ mprj_io_ib_mode_sel[24] porb_h porb_h mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD mprj_io_oeb[24]
+ mprj_pads.area2_io_pad\[10\]/HLD_H_N mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD mprj_io_slow_sel[24]
+ mprj_io_vtrip_sel[24] mprj_io_holdover[24] mprj_io_analog_en[24] mprj_io_analog_sel[24]
+ mprj_io_one[24] mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD mprj_io_analog_pol[24] mprj_io_out[24]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_606 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_628 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_639 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_95 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_84 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_73 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_469 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_458 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_447 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_436 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_403 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_414 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_425 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[0\] mprj_io_in_3v3[14] mprj_gpio_noesd[7] mprj_gpio_analog[7]
+ mprj_pads.area2_io_pad\[0\]/PAD_A_ESD_1_H mprj_io[25] mprj_io_dm[44] mprj_io_dm[43]
+ mprj_io_dm[42] mprj_pads.area2_io_pad\[0\]/HLD_H_N mprj_io_in[14] mprj_io_inp_dis[14]
+ mprj_io_ib_mode_sel[14] porb_h porb_h mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD mprj_io_oeb[14]
+ mprj_pads.area2_io_pad\[0\]/HLD_H_N mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD mprj_io_slow_sel[14]
+ mprj_io_vtrip_sel[14] mprj_io_holdover[14] mprj_io_analog_en[14] mprj_io_analog_sel[14]
+ mprj_io_one[14] mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD mprj_io_analog_pol[14] mprj_io_out[14]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_233 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_211 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_200 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_244 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_288 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_299 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser1_analog_pad\[2\] mprj_analog[3] vssa1 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda1 vccd vccd gpio_pad/VSSIO_Q mprj_io[17]
+ sky130_ef_io__analog_pad
XFILLER_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_607 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_618 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_629 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_96 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_85 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_30 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[0\] mprj_io_in_3v3[0] mprj_pads.area1_io_pad\[0\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_1_H
+ mprj_io[0] mprj_io_dm[2] mprj_io_dm[1] mprj_io_dm[0] mprj_pads.area1_io_pad\[0\]/HLD_H_N
+ mprj_io_in[0] mprj_io_inp_dis[0] mprj_io_ib_mode_sel[0] porb_h porb_h mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_oeb[0] mprj_pads.area1_io_pad\[0\]/HLD_H_N mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_slow_sel[0] mprj_io_vtrip_sel[0] mprj_io_holdover[0] mprj_io_analog_en[0]
+ mprj_io_analog_sel[0] mprj_io_one[0] mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD mprj_io_analog_pol[0]
+ mprj_io_out[0] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_459 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_448 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_437 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_404 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_415 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_426 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_234 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_212 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_201 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_245 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_267 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_278 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_619 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_86 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_449 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_438 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_405 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_416 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_427 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_235 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_213 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_202 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_246 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_268 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_279 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_780 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
XFILLER_609 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_98 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_87 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_43 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_439 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_406 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_417 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_428 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_236 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_214 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_203 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_247 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_269 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_781 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_770 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_analog_pad\[0\] mprj_analog[1] vssa1 vssd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ gpio_pad/VDDIO_Q vddio vddio vssio vdda1 vccd vccd gpio_pad/VSSIO_Q mprj_io[15]
+ sky130_ef_io__analog_pad
Xflash_io0_pad flash_io0_pad/IN_H flash_io0_pad/PAD_A_NOESD_H flash_io0_pad/PAD_A_ESD_0_H
+ flash_io0_pad/PAD_A_ESD_1_H flash_io0 flash_io0_ieb_core flash_io0_ieb_core flash_io0_oeb_core
+ flash_io0_pad/HLD_H_N flash_io0_di_core flash_io0_ieb_core flash_io0_pad/SLOW porb_h
+ porb_h flash_io0_pad/TIE_LO_ESD flash_io0_oeb_core flash_io0_pad/HLD_H_N flash_io0_pad/TIE_LO_ESD
+ flash_io0_pad/SLOW flash_io0_pad/SLOW flash_io0_pad/SLOW flash_io0_pad/SLOW flash_io0_pad/SLOW
+ constant_block_4/one flash_io0_pad/TIE_LO_ESD flash_io0_pad/SLOW flash_io0_do_core
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[9\] mprj_io_in_3v3[23] mprj_gpio_noesd[16] mprj_gpio_analog[16]
+ mprj_pads.area2_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[34] mprj_io_dm[71] mprj_io_dm[70]
+ mprj_io_dm[69] mprj_pads.area2_io_pad\[9\]/HLD_H_N mprj_io_in[23] mprj_io_inp_dis[23]
+ mprj_io_ib_mode_sel[23] porb_h porb_h mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD mprj_io_oeb[23]
+ mprj_pads.area2_io_pad\[9\]/HLD_H_N mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD mprj_io_slow_sel[23]
+ mprj_io_vtrip_sel[23] mprj_io_holdover[23] mprj_io_analog_en[23] mprj_io_analog_sel[23]
+ mprj_io_one[23] mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD mprj_io_analog_pol[23] mprj_io_out[23]
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_99 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_88 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_407 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_418 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_429 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_237 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_248 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_782 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_771 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_760 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_corner\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
XFILLER_590 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vssa_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[9\] mprj_io_in_3v3[9] mprj_gpio_noesd[2] mprj_gpio_analog[2]
+ mprj_pads.area1_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[9] mprj_io_dm[29] mprj_io_dm[28]
+ mprj_io_dm[27] mprj_pads.area1_io_pad\[9\]/HLD_H_N mprj_io_in[9] mprj_io_inp_dis[9]
+ mprj_io_ib_mode_sel[9] mprj_pads.area1_io_pad\[9\]/ENABLE_H mprj_pads.area1_io_pad\[9\]/ENABLE_H
+ mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD mprj_io_oeb[9] mprj_pads.area1_io_pad\[9\]/HLD_H_N
+ mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD mprj_io_slow_sel[9] mprj_io_vtrip_sel[9]
+ mprj_io_holdover[9] mprj_io_analog_en[9] mprj_io_analog_sel[9] mprj_io_one[9] mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD
+ mprj_io_analog_pol[9] mprj_io_out[9] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_89 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_78 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_56 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xconstant_block_0 constant_block_0/one vccd vssd constant_block_0/zero constant_block
Xflash_clk_pad flash_clk_pad/IN_H flash_clk_pad/PAD_A_NOESD_H flash_clk_pad/PAD_A_ESD_0_H
+ flash_clk_pad/PAD_A_ESD_1_H flash_clk flash_clk_pad/DM[2] flash_clk_pad/DM[2] flash_clk_pad/SLOW
+ flash_clk_pad/HLD_H_N flash_clk_pad/IN flash_clk_pad/SLOW flash_clk_pad/SLOW porb_h
+ porb_h flash_clk_pad/TIE_LO_ESD flash_clk_oeb_core flash_clk_pad/HLD_H_N flash_clk_pad/TIE_LO_ESD
+ flash_clk_pad/SLOW flash_clk_pad/SLOW flash_clk_pad/SLOW flash_clk_pad/SLOW flash_clk_pad/SLOW
+ flash_clk_pad/DM[2] flash_clk_pad/TIE_LO_ESD flash_clk_pad/SLOW flash_clk_core gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q
+ sky130_ef_io__gpiov2_pad_wrapped
XFILLER_408 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_419 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_227 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_216 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_783 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_772 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_761 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_750 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q vccd1 vssd1 sky130_ef_io__vccd_lvc_clamped3_pad
XFILLER_580 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_591 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[13\] mprj_io_in_3v3[13] mprj_gpio_noesd[6] mprj_gpio_analog[6]
+ mprj_pads.area1_io_pad\[13\]/PAD_A_ESD_1_H mprj_io[13] mprj_io_dm[41] mprj_io_dm[40]
+ mprj_io_dm[39] mprj_pads.area1_io_pad\[13\]/HLD_H_N mprj_io_in[13] mprj_io_inp_dis[13]
+ mprj_io_ib_mode_sel[13] mprj_pads.area1_io_pad\[13\]/ENABLE_H mprj_pads.area1_io_pad\[13\]/ENABLE_H
+ mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD mprj_io_oeb[13] mprj_pads.area1_io_pad\[13\]/HLD_H_N
+ mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD mprj_io_slow_sel[13] mprj_io_vtrip_sel[13]
+ mprj_io_holdover[13] mprj_io_analog_en[13] mprj_io_analog_sel[13] mprj_io_one[13]
+ mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD mprj_io_analog_pol[13] mprj_io_out[13] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_79 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
XFILLER_409 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xconstant_block_1 clock_pad/OE_N vccd vssd clock_pad/OUT constant_block
XFILLER_228 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_217 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_784 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_773 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_762 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_751 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_740 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VGND VPWR clk_in clk_out core_clk core_rstn debug_in debug_mode
+ debug_oeb debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb
+ flash_io1_di flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb
+ flash_io3_di flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad
+ gpio_mode1_pad gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10]
+ hk_dat_i[11] hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17]
+ hk_dat_i[18] hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23]
+ hk_dat_i[24] hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2]
+ hk_dat_i[30] hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7]
+ hk_dat_i[8] hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0]
+ la_iena[100] la_iena[101] la_iena[102] la_iena[103] la_iena[104] la_iena[105] la_iena[106]
+ la_iena[107] la_iena[108] la_iena[109] la_iena[10] la_iena[110] la_iena[111] la_iena[112]
+ la_iena[113] la_iena[114] la_iena[115] la_iena[116] la_iena[117] la_iena[118] la_iena[119]
+ la_iena[11] la_iena[120] la_iena[121] la_iena[122] la_iena[123] la_iena[124] la_iena[125]
+ la_iena[126] la_iena[127] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16]
+ la_iena[17] la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22]
+ la_iena[23] la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29]
+ la_iena[2] la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35]
+ la_iena[36] la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41]
+ la_iena[42] la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48]
+ la_iena[49] la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54]
+ la_iena[55] la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60]
+ la_iena[61] la_iena[62] la_iena[63] la_iena[64] la_iena[65] la_iena[66] la_iena[67]
+ la_iena[68] la_iena[69] la_iena[6] la_iena[70] la_iena[71] la_iena[72] la_iena[73]
+ la_iena[74] la_iena[75] la_iena[76] la_iena[77] la_iena[78] la_iena[79] la_iena[7]
+ la_iena[80] la_iena[81] la_iena[82] la_iena[83] la_iena[84] la_iena[85] la_iena[86]
+ la_iena[87] la_iena[88] la_iena[89] la_iena[8] la_iena[90] la_iena[91] la_iena[92]
+ la_iena[93] la_iena[94] la_iena[95] la_iena[96] la_iena[97] la_iena[98] la_iena[99]
+ la_iena[9] la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105]
+ la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124]
+ la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66]
+ la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72]
+ la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79]
+ la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85]
+ la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91]
+ la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98]
+ la_oenb[99] la_oenb[9] la_output[0] la_output[100] la_output[101] la_output[102]
+ la_output[103] la_output[104] la_output[105] la_output[106] la_output[107] la_output[108]
+ la_output[109] la_output[10] la_output[110] la_output[111] la_output[112] la_output[113]
+ la_output[114] la_output[115] la_output[116] la_output[117] la_output[118] la_output[119]
+ la_output[11] la_output[120] la_output[121] la_output[122] la_output[123] la_output[124]
+ la_output[125] la_output[126] la_output[127] la_output[12] la_output[13] la_output[14]
+ la_output[15] la_output[16] la_output[17] la_output[18] la_output[19] la_output[1]
+ la_output[20] la_output[21] la_output[22] la_output[23] la_output[24] la_output[25]
+ la_output[26] la_output[27] la_output[28] la_output[29] la_output[2] la_output[30]
+ la_output[31] la_output[32] la_output[33] la_output[34] la_output[35] la_output[36]
+ la_output[37] la_output[38] la_output[39] la_output[3] la_output[40] la_output[41]
+ la_output[42] la_output[43] la_output[44] la_output[45] la_output[46] la_output[47]
+ la_output[48] la_output[49] la_output[4] la_output[50] la_output[51] la_output[52]
+ la_output[53] la_output[54] la_output[55] la_output[56] la_output[57] la_output[58]
+ la_output[59] la_output[5] la_output[60] la_output[61] la_output[62] la_output[63]
+ la_output[64] la_output[65] la_output[66] la_output[67] la_output[68] la_output[69]
+ la_output[6] la_output[70] la_output[71] la_output[72] la_output[73] la_output[74]
+ la_output[75] la_output[76] la_output[77] la_output[78] la_output[79] la_output[7]
+ la_output[80] la_output[81] la_output[82] la_output[83] la_output[84] la_output[85]
+ la_output[86] la_output[87] la_output[88] la_output[89] la_output[8] la_output[90]
+ la_output[91] la_output[92] la_output[93] la_output[94] la_output[95] la_output[96]
+ la_output[97] la_output[98] la_output[99] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o por_l_in por_l_out porb_h_in porb_h_out qspi_enabled resetn_in resetn_out
+ rstb_l_in rstb_l_out ser_rx ser_tx serial_clock_in serial_clock_out serial_data_2_in
+ serial_data_2_out serial_load_in serial_load_out serial_resetn_in serial_resetn_out
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb trap uart_enabled user_irq_ena[0]
+ user_irq_ena[1] user_irq_ena[2]
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_sc_hvl__buf_8 A VGND VPWR X VNB VPB
X0 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X3 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X5 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X7 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X9 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X10 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X11 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X12 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X14 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X15 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X16 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X17 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X18 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X21 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_n1806_2500# a_n4122_n2932# a_n5280_2500#
+ a_2054_n2932# a_896_n2932# a_4756_2500# a_3598_n2932# a_3212_2500# a_n3736_n2932#
+ a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_896_2500# a_510_n2932# a_n3350_2500#
+ a_n4508_2500# a_3212_n2932# a_n4894_2500# a_n5410_n3062# a_1282_2500# a_4756_n2932#
+ a_2826_2500# a_2826_n2932# a_n2192_n2932# a_n1034_2500# a_n2578_2500# a_n1420_2500#
+ a_n2964_2500# a_n648_n2932# a_n648_2500# a_n5280_n2932# a_n3350_n2932# a_4370_2500#
+ a_1282_n2932# a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_124_2500# a_n2964_n2932#
+ a_n4122_2500# a_2054_2500# a_510_2500# a_n4508_n2932# a_4370_n2932# a_3598_2500#
+ a_3984_2500# a_2440_n2932# a_2440_2500# a_3984_n2932# a_n2192_2500# a_n3736_2500#
+ a_1668_2500# a_n262_n2932# a_n262_2500# a_n1034_n2932# a_5142_2500# a_n2578_n2932#
X0 a_n2578_n2932# a_n2578_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X1 a_n1420_n2932# a_n1420_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X2 a_n1806_n2932# a_n1806_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X3 a_3212_n2932# a_3212_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X4 a_3598_n2932# a_3598_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X5 a_n2964_n2932# a_n2964_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X6 a_2826_n2932# a_2826_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X7 a_4370_n2932# a_4370_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X8 a_3984_n2932# a_3984_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X9 a_n262_n2932# a_n262_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X10 a_n3350_n2932# a_n3350_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X11 a_n4122_n2932# a_n4122_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X12 a_n3736_n2932# a_n3736_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X13 a_5142_n2932# a_5142_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X14 a_n4894_n2932# a_n4894_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X15 a_1282_n2932# a_1282_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X16 a_4756_n2932# a_4756_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X17 a_124_n2932# a_124_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X18 a_510_n2932# a_510_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X19 a_896_n2932# a_896_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X20 a_n648_n2932# a_n648_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X21 a_n5280_n2932# a_n5280_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X22 a_n4508_n2932# a_n4508_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X23 a_n1034_n2932# a_n1034_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X24 a_n2192_n2932# a_n2192_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X25 a_2054_n2932# a_2054_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X26 a_1668_n2932# a_1668_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
X27 a_2440_n2932# a_2440_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=2.5e+07u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VPWR X VNB VPB
X0 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X1 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X4 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=290000u l=1.355e+06u
X5 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=290000u l=3.11e+06u
X6 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X7 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PKVMTM a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=800000u
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X15 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
.ends

.subckt simple_por vdd3v3 vdd1v8 porb_h por_l porb_l vss1v8 vss3v3
Xsky130_fd_pr__cap_mim_m3_2_W5U4AW_0 vss3v3 sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_W5U4AW
Xsky130_fd_sc_hvl__buf_8_1 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vdd1v8 porb_l vss1v8
+ vdd1v8 sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss3v3 m1_721_6815# vss3v3 vss3v3
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815#
+ vss3v3 m1_721_6815# vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 li_3322_5813# li_1391_165# vss3v3 li_7567_165#
+ li_6023_165# vdd3v3 li_9111_165# li_8726_5813# li_1391_165# li_6795_165# li_3707_165#
+ vss3v3 li_6410_5813# li_6023_165# li_1778_5813# li_1006_5813# li_8339_165# vss3v3
+ vss3v3 li_6410_5813# li_9883_165# li_7954_5813# li_8339_165# li_2935_165# li_4094_5813#
+ li_2550_5813# li_4094_5813# li_2550_5813# li_4479_165# li_4866_5813# vss3v3 li_2163_165#
+ li_9498_5813# li_6795_165# li_5251_165# li_3707_165# li_619_165# li_5638_5813# li_2163_165#
+ li_1006_5813# li_7182_5813# li_5638_5813# li_619_165# li_9883_165# li_8726_5813#
+ li_9498_5813# li_7567_165# li_7954_5813# li_9111_165# li_3322_5813# li_1778_5813#
+ li_7182_5813# li_5251_165# li_4866_5813# li_4479_165# vss3v3 li_2935_165# sky130_fd_pr__res_xhigh_po_0p69_S5N9F3
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_2756_6573# m1_4283_8081# vdd3v3 m1_2756_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 vdd3v3
+ sky130_fd_sc_hvl__inv_8_0/A vss3v3 vdd3v3 sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6573# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 m1_6249_7690# sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 m1_2756_6573# vss3v3 vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_PKVMTM
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 m1_185_6573# vss3v3 vss3v3 li_2550_5813# sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_1_WRT4AW_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 sky130_fd_pr__cap_mim_m3_1_WRT4AW
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__buf_8_0 sky130_fd_sc_hvl__inv_8_0/A vss3v3 vdd3v3 porb_h vss3v3
+ vdd3v3 sky130_fd_sc_hvl__buf_8
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vdd1v8 por_l vss1v8
+ vdd1v8 sky130_fd_sc_hvl__inv_8
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 A B VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VPWR Y VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_531_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C_N a_531_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_281_297# a_531_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y a_531_21# a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND C_N a_531_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y a_531_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X5 a_1228_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_1602_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1028_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND a_1602_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1028_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X25 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1300_47# a_1178_261# a_1228_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X30 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VGND SET_B a_1300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VPWR Y VNB VPB
X0 VGND A_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y a_27_93# a_206_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_206_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VPWR Y VNB VPB
X0 VGND B_N a_27_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_496_21# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 Y a_496_21# a_426_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_496_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_426_47# a_27_93# a_326_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B_N a_27_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_496_21# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y a_27_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_218_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_326_47# C a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VPWR Q VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VPWR X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VPWR Y VNB VPB
X0 VPWR A2_N a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y a_112_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B2 a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_112_297# A2_N a_112_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_112_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_112_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B1 a_478_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_394_47# a_112_297# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_394_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_478_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VPWR Y VNB VPB
X0 VPWR A a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_193_297# B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_12 A VGND VPWR X VNB VPB
X0 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VPWR Y VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VPWR Y VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_298_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_664_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_298_47# B1 a_497_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_497_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_497_47# B1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y A2 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_27_47# C1 a_298_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_497_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR A1 a_664_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_664_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 a_281_297# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y A3 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A2 a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VPWR X VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VPWR Y VNB VPB
X0 a_236_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_428_47# A2 a_336_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A1 a_428_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_336_47# A3 a_236_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR A4 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VPWR Q VNB VPB
X0 a_1217_47# a_193_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_27_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_193_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_193_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_193_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_27_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_27_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_235_47# C1 a_163_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_343_47# B1 a_235_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_454_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_454_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_163_47# D1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND A2 a_343_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_343_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VPWR Y VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VPWR Y VNB VPB
X0 Y C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_281_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VPWR X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VPWR Y VNB VPB
X0 a_388_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_105_352# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_297_47# a_105_352# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_388_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1_N a_105_352# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 Y a_105_352# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4 A VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VPWR Q VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VPWR Y VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 Y B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A3 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VPWR Y VNB VPB
X0 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_806_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# B1 a_1314_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y A2 a_110_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y C1 a_978_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 Y C1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_27_47# B1 a_806_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_110_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_806_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 a_978_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_1314_47# C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VPWR X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VPWR Y VNB VPB
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_191_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_297_297# B a_191_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt caravel_clocking core_clk ext_clk ext_clk_sel ext_reset pll_clk pll_clk90
+ resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk VGND VPWR
XFILLER_26_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_432_ _204_/A1 _432_/D _372_/S VGND VPWR _432_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_294_ _429_/Q _430_/Q VGND VPWR _294_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_363_ _365_/A _429_/Q VGND VPWR _363_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_8_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_415_ _204_/A1 _440_/Q _372_/S VGND VPWR _415_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_346_ _416_/D _292_/Y _419_/Q VGND VPWR _347_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_277_ _422_/Q _423_/Q _421_/Q VGND VPWR _277_/Y VGND VPWR sky130_fd_sc_hd__nor3b_2
XFILLER_23_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_329_ _329_/A _329_/B VGND VPWR _329_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_6_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__037_ clkbuf_0__037_/X VGND VPWR _208_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_431_ _204_/A1 _431_/D _372_/S VGND VPWR _431_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_13_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_293_ _223_/S _365_/A VGND VPWR _293_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_9_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_362_ _295_/C _293_/Y _361_/Y VGND VPWR _428_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
XANTENNA__265__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_345_ _311_/C _419_/Q _345_/C _431_/Q VGND VPWR _347_/A VGND VPWR sky130_fd_sc_hd__nand4bb_1
X_414_ _207_/A1 _414_/D fanout27/X VGND VPWR _414_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_276_ _426_/Q _210_/X _360_/S VGND VPWR _426_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_328_ _442_/D _441_/D _327_/A VGND VPWR _329_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA__395__B1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_29_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_292_ _431_/Q _345_/C VGND VPWR _292_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_13_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_430_ _456_/CLK _430_/D fanout26/X VGND VPWR _430_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_361_ _223_/S _280_/X _219_/X VGND VPWR _361_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_413_ _204_/A1 _413_/D _372_/S VGND VPWR _413_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_344_ _414_/Q _342_/Y _343_/Y VGND VPWR _414_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_275_ _232_/X _273_/Y _274_/Y _234_/S VGND VPWR _447_/D VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
XFILLER_5_131 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_258_ _258_/A VGND VPWR _258_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_9_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_327_ _327_/A _442_/D _441_/D VGND VPWR _329_/A VGND VPWR sky130_fd_sc_hd__nor3_1
XANTENNA__452__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput11 _341_/Y VGND VPWR resetb_sync VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_16_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_291_ _432_/Q _433_/Q VGND VPWR _345_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_26_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_360_ _427_/Q _211_/X _360_/S VGND VPWR _427_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_412_ _456_/CLK _412_/D fanout26/X VGND VPWR _413_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_343_ _342_/Y _414_/Q _234_/S VGND VPWR _343_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_274_ _385_/B _447_/Q VGND VPWR _274_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_5_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_326_ _451_/Q _450_/Q VGND VPWR _326_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_257_ _257_/A VGND VPWR _257_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_18_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__395__A2 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_309_ _311_/B _311_/C VGND VPWR _309_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
Xclkbuf_0_divider.out _304_/Y VGND VPWR clkbuf_0_divider.out/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_6_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_131 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input8_A sel[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_7_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_290_ _215_/X _288_/Y _289_/Y _219_/S VGND VPWR _422_/D VGND VPWR sky130_fd_sc_hd__o2bb2ai_1
Xclkbuf_0_pll_clk pll_clk VGND VPWR clkbuf_0_pll_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_12_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_411_ _411_/CLK _411_/D _372_/S VGND VPWR _411_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_273_ _234_/S _385_/B VGND VPWR _273_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
X_342_ _327_/A _442_/D _441_/D _453_/Q _299_/Y VGND VPWR _342_/Y VGND VPWR sky130_fd_sc_hd__o2111ai_2
XANTENNA__446__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_23_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_325_ _442_/D _441_/D VGND VPWR _325_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_308_ _307_/Y _298_/B _306_/X _305_/Y VGND VPWR _308_/Y VGND VPWR sky130_fd_sc_hd__o31ai_2
XFILLER_1_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_239_ _339_/Y _327_/A _300_/Y VGND VPWR _239_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__451__SET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_31_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VPWR _455_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_12_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_341_ _341_/A _409_/Q VGND VPWR _341_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_410_ _410_/CLK _411_/Q _372_/S VGND VPWR _410_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_272_ _263_/Y _265_/X _234_/S VGND VPWR _272_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_4_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_324_ _432_/Q _431_/Q VGND VPWR _324_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_9_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_255_ _255_/A VGND VPWR _255_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_18_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_307_ _449_/Q _414_/Q VGND VPWR _307_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_238_ _237_/X _442_/D _240_/S VGND VPWR _238_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_340_ _458_/Q _457_/Q VGND VPWR _340_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_271_ _271_/A _271_/B VGND VPWR _449_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_5_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__455__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_9_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_323_ _321_/Y _323_/B VGND VPWR _323_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_2_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA__240__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_306_ _449_/Q _414_/Q VGND VPWR _306_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_237_ _336_/Y _442_/D _300_/Y VGND VPWR _237_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__213__A1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input6_A sel2[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_270_ _262_/Y _263_/Y _265_/X _243_/Y _234_/S VGND VPWR _271_/B VGND VPWR sky130_fd_sc_hd__a41oi_1
X_399_ _242_/X _458_/Q _400_/A VGND VPWR _458_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_322_ _428_/Q _429_/Q _430_/Q VGND VPWR _323_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_2_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_net10 clkbuf_0_net10/X VGND VPWR core_clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_1_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_253_ _253_/A VGND VPWR _412_/D VGND VPWR sky130_fd_sc_hd__clkinv_4
X_305_ _441_/D _305_/B VGND VPWR _305_/Y VGND VPWR sky130_fd_sc_hd__nand2b_2
X_236_ _235_/X _441_/D _240_/S VGND VPWR _236_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout27_A fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_219_ _218_/X _311_/C _219_/S VGND VPWR _219_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_398_ _241_/X _457_/Q _400_/A VGND VPWR _457_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_252_ _453_/Q VGND VPWR _300_/C VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_1_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_321_ _428_/Q _429_/Q _430_/Q VGND VPWR _321_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_304_ _303_/Y _365_/A _302_/X _301_/Y VGND VPWR _304_/Y VGND VPWR sky130_fd_sc_hd__o31ai_2
X_235_ _300_/C _441_/D _300_/Y VGND VPWR _235_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_218_ _295_/C _311_/C _295_/Y VGND VPWR _218_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xuser_clk_out_buffer _208_/X VGND VPWR user_clk VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_21_186 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_397_ _456_/Q _395_/Y _396_/Y VGND VPWR _456_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_251_ _446_/Q VGND VPWR _251_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_320_ _428_/Q _429_/Q VGND VPWR _320_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_449_ _449_/CLK _449_/D fanout27/X VGND VPWR _449_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XANTENNA__234__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider.out clkbuf_0_divider.out/X VGND VPWR _206_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_303_ _424_/Q _456_/Q VGND VPWR _303_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_234_ _233_/X _327_/A _234_/S VGND VPWR _260_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_217_ _216_/X _351_/A _223_/S VGND VPWR _257_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__328__B1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_465_ _208_/A1 _465_/D fanout27/X VGND VPWR _465_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_396_ _395_/Y _456_/Q _223_/S VGND VPWR _396_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
Xfanout20 _437_/Q VGND VPWR _416_/D VGND VPWR sky130_fd_sc_hd__clkbuf_2
XANTENNA_input4_A sel2[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_13_63 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_250_ _450_/Q VGND VPWR _250_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_379_ _465_/Q _443_/Q VGND VPWR _379_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_448_ _455_/CLK _448_/D fanout28/X VGND VPWR _448_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_24_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_302_ _424_/Q _456_/Q VGND VPWR _302_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_233_ _335_/Y _327_/A _262_/Y VGND VPWR _233_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_216_ _319_/Y _351_/A _277_/Y VGND VPWR _216_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__282__B1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_12_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_259__1 _455_/CLK VGND VPWR _447_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_464_ _464_/CLK _464_/D fanout27/X VGND VPWR _464_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_395_ _351_/A _311_/B _311_/C _428_/Q _294_/Y VGND VPWR _395_/Y VGND VPWR sky130_fd_sc_hd__o2111ai_1
XFILLER_4_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout21 _234_/S VGND VPWR _240_/S VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_447_ _447_/CLK _447_/D fanout28/X VGND VPWR _447_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_378_ _378_/A _378_/B _441_/Q VGND VPWR _378_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_1_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_301_ _416_/D _301_/B VGND VPWR _301_/Y VGND VPWR sky130_fd_sc_hd__nand2b_2
X_232_ _231_/X _442_/D _234_/S VGND VPWR _232_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__037_ clkbuf_0__037_/X VGND VPWR _206_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_28_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_215_ _214_/X _311_/B _219_/S VGND VPWR _215_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_463_ _464_/CLK _463_/D fanout27/X VGND VPWR _463_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_394_ _240_/S _455_/Q _265_/X _393_/Y VGND VPWR _455_/D VGND VPWR sky130_fd_sc_hd__o31a_1
Xfanout22 _445_/Q VGND VPWR _234_/S VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_1__f_pll_clk90 clkbuf_0_pll_clk90/X VGND VPWR _207_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_377_ _442_/Q _464_/Q VGND VPWR _378_/B VGND VPWR sky130_fd_sc_hd__nand2b_1
X_446_ _455_/CLK _446_/D fanout28/X VGND VPWR _446_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__219__A1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_406__6 _204_/A1 VGND VPWR _426_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
Xclkbuf_0_ext_clk ext_clk VGND VPWR clkbuf_0_ext_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_231_ _332_/Y _442_/D _262_/Y VGND VPWR _231_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_300_ _454_/Q _455_/Q _300_/C VGND VPWR _300_/Y VGND VPWR sky130_fd_sc_hd__nor3_2
X_429_ _456_/CLK _429_/D fanout26/X VGND VPWR _429_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_19_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput1 ext_clk_sel VGND VPWR _253_/A VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_214_ _316_/Y _311_/B _277_/Y VGND VPWR _214_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__282__A2 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_462_ _208_/A1 _462_/D fanout27/X VGND VPWR _465_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_27_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_393_ _240_/S _265_/X _240_/X VGND VPWR _393_/Y VGND VPWR sky130_fd_sc_hd__o21bai_1
Xfanout23 _223_/S VGND VPWR _219_/S VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_445_ _207_/A1 _445_/D fanout28/X VGND VPWR _445_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_376_ _464_/Q _442_/Q VGND VPWR _378_/A VGND VPWR sky130_fd_sc_hd__nand2b_1
X_256__4 _456_/CLK VGND VPWR _422_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XANTENNA_input2_A ext_reset VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_230_ _229_/X _441_/D _234_/S VGND VPWR _258_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_359_ _425_/Q _209_/X _360_/S VGND VPWR _425_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_428_ _456_/CLK _428_/D fanout26/X VGND VPWR _428_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xinput2 ext_reset VGND VPWR _341_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_27_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_213_ _212_/X _311_/C _219_/S VGND VPWR _255_/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_403__8 _403__8/A VGND VPWR _410_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_18_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_net10 _206_/X VGND VPWR clkbuf_0_net10/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_21_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_461_ _464_/CLK _461_/D fanout27/X VGND VPWR _464_/D VGND VPWR sky130_fd_sc_hd__dfstp_1
X_392_ _240_/S _454_/Q _265_/X _391_/Y VGND VPWR _454_/D VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_4_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout13 _465_/Q VGND VPWR _327_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout24 _420_/Q VGND VPWR _223_/S VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_1_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_444_ _207_/A1 _444_/D fanout27/X VGND VPWR _444_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_375_ _375_/A _375_/B VGND VPWR _444_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_24_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_427_ _456_/CLK _427_/D fanout26/X VGND VPWR _427_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_358_ _257_/Y _287_/Y _357_/Y VGND VPWR _423_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
Xinput3 resetb VGND VPWR input3/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__327__A _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_289_ _357_/B _422_/Q VGND VPWR _289_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_212_ _247_/Y _311_/C _277_/Y VGND VPWR _212_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__267__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_411__30 VGND VGND VPWR VPWR _411__30/HI _411_/D sky130_fd_sc_hd__conb_1
XANTENNA__445__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_460_ _464_/CLK _460_/D fanout27/X VGND VPWR _463_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_391_ _240_/S _265_/X _238_/X VGND VPWR _391_/Y VGND VPWR sky130_fd_sc_hd__o21bai_1
XFILLER_4_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout25 fanout29/X VGND VPWR _372_/S VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout14 _464_/Q VGND VPWR _442_/D VGND VPWR sky130_fd_sc_hd__buf_4
X_374_ _400_/A _297_/Y _444_/Q VGND VPWR _375_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_443_ _207_/A1 _465_/Q VGND VPWR _443_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput4 sel2[0] VGND VPWR _460_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_426_ _426_/CLK _426_/D fanout26/X VGND VPWR _426_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_288_ _219_/S _357_/B VGND VPWR _288_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
X_357_ _219_/S _357_/B _423_/Q VGND VPWR _357_/Y VGND VPWR sky130_fd_sc_hd__nand3b_1
X_211_ _315_/X _313_/B _223_/S VGND VPWR _211_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_409_ _409_/CLK _410_/Q fanout27/X VGND VPWR _409_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_24_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_390_ _300_/C _298_/Y _389_/Y VGND VPWR _453_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_4_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout15 _463_/Q VGND VPWR _441_/D VGND VPWR sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f_pll_clk clkbuf_0_pll_clk/X VGND VPWR _204_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xfanout26 fanout29/X VGND VPWR fanout26/X VGND VPWR sky130_fd_sc_hd__buf_4
X_373_ _400_/A _444_/Q _373_/C _457_/Q VGND VPWR _375_/A VGND VPWR sky130_fd_sc_hd__nand4bb_1
XANTENNA__312__A1 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_442_ _455_/CLK _442_/D VGND VPWR _442_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_0_170 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA__345__A_N _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__447__SET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput5 sel2[1] VGND VPWR _461_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_425_ _456_/CLK _425_/D fanout26/X VGND VPWR _425_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_287_ _278_/Y _280_/X _219_/S VGND VPWR _287_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_356_ _255_/Y _287_/Y _355_/Y VGND VPWR _421_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_19_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_210_ _310_/Y _313_/Y _223_/S VGND VPWR _210_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f_divider2.out clkbuf_0_divider2.out/X VGND VPWR _464_/CLK VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
X_339_ _337_/Y _339_/B VGND VPWR _339_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_2_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__264__A _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout16 _463_/Q VGND VPWR _400_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xfanout27 fanout28/X VGND VPWR fanout27/X VGND VPWR sky130_fd_sc_hd__buf_4
X_372_ _440_/Q _372_/A1 _372_/S VGND VPWR _440_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_441_ _455_/CLK _441_/D VGND VPWR _441_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_13_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__312__A2 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_24_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_424_ _424_/CLK _424_/D fanout26/X VGND VPWR _424_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_286_ _286_/A _286_/B VGND VPWR _424_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_355_ _219_/S _357_/B _421_/Q VGND VPWR _355_/Y VGND VPWR sky130_fd_sc_hd__nand3b_1
Xinput6 sel2[2] VGND VPWR _462_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__221__A1 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__212__A1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_269_ _262_/Y _263_/Y _265_/X _243_/Y VGND VPWR _271_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_338_ _454_/Q _453_/Q _455_/Q VGND VPWR _339_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_32_170 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__037_ _205_/X VGND VPWR clkbuf_0__037_/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_4_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout28 fanout29/X VGND VPWR fanout28/X VGND VPWR sky130_fd_sc_hd__buf_4
X_371_ _369_/Y _371_/B VGND VPWR _433_/D VGND VPWR sky130_fd_sc_hd__nand2b_1
X_440_ _204_/A1 _440_/D VGND VPWR _440_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
Xfanout17 _439_/Q VGND VPWR _351_/A VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_0_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_354_ _223_/S _280_/X _352_/Y _353_/Y VGND VPWR _420_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_14_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_285_ _277_/Y _278_/Y _280_/X _244_/Y _223_/S VGND VPWR _286_/B VGND VPWR sky130_fd_sc_hd__a41oi_1
X_423_ _456_/CLK _423_/D fanout26/X VGND VPWR _423_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XANTENNA__448__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xinput7 sel[0] VGND VPWR _434_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_268_ _385_/B VGND VPWR _268_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_337_ _454_/Q _453_/Q _455_/Q VGND VPWR _337_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_15_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_138 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_divider.out clkbuf_0_divider.out/X VGND VPWR _439_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_11_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__342__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xfanout29 input3/X VGND VPWR fanout29/X VGND VPWR sky130_fd_sc_hd__buf_2
Xfanout18 _438_/Q VGND VPWR _311_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_370_ _416_/D _432_/Q _431_/Q _433_/Q VGND VPWR _371_/B VGND VPWR sky130_fd_sc_hd__o31ai_1
XANTENNA__242__A0 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_353_ _353_/A _353_/B _416_/Q VGND VPWR _353_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_284_ _277_/Y _278_/Y _280_/X _244_/Y VGND VPWR _286_/A VGND VPWR sky130_fd_sc_hd__a31o_1
X_422_ _422_/CLK _422_/D fanout26/X VGND VPWR _422_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
Xclkbuf_1_0__f_pll_clk clkbuf_0_pll_clk/X VGND VPWR _456_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xinput8 sel[1] VGND VPWR _435_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_267_ _327_/A _442_/D _441_/D _263_/Y VGND VPWR _385_/B VGND VPWR sky130_fd_sc_hd__o211ai_4
X_336_ _454_/Q _453_/Q VGND VPWR _336_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_32_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_319_ _317_/Y _319_/B VGND VPWR _319_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_11_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout19 _437_/Q VGND VPWR _311_/C VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_12_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input9_A sel[2] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__233__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA__215__A1 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_421_ _456_/CLK _421_/D fanout26/X VGND VPWR _421_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_352_ _350_/Y _351_/X _280_/X VGND VPWR _352_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
Xinput9 sel[2] VGND VPWR _436_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_283_ _357_/B VGND VPWR _283_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_407__2 _207_/A1 VGND VPWR _449_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XPHY_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_266_ _327_/A _464_/Q _400_/A VGND VPWR _298_/B VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_18_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_335_ _333_/Y _335_/B VGND VPWR _335_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_24_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_249_ _457_/Q VGND VPWR _249_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_318_ _422_/Q _421_/Q _423_/Q VGND VPWR _319_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_22_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_divider2.out _308_/Y VGND VPWR clkbuf_0_divider2.out/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_351_ _351_/A _418_/Q VGND VPWR _351_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_420_ _204_/A1 _420_/D _372_/S VGND VPWR _420_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_282_ _351_/A _311_/B _311_/C _278_/Y VGND VPWR _357_/B VGND VPWR sky130_fd_sc_hd__o211ai_4
XFILLER_27_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_334_ _447_/Q _446_/Q _448_/Q VGND VPWR _335_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_265_ _327_/A _442_/D _441_/D VGND VPWR _265_/X VGND VPWR sky130_fd_sc_hd__o21a_2
XFILLER_14_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_248_ _428_/Q VGND VPWR _295_/C VGND VPWR sky130_fd_sc_hd__clkinv_4
X_317_ _422_/Q _421_/Q _423_/Q VGND VPWR _317_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__281__B1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_281_ _351_/A _311_/B _311_/C VGND VPWR _365_/A VGND VPWR sky130_fd_sc_hd__o21ai_2
X_350_ _351_/A _418_/Q VGND VPWR _350_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_14_74 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_402_ _400_/Y _402_/B VGND VPWR _459_/D VGND VPWR sky130_fd_sc_hd__nand2b_1
X_264_ _327_/A _464_/Q VGND VPWR _264_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_333_ _447_/Q _446_/Q _448_/Q VGND VPWR _333_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_2_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_316_ _422_/Q _421_/Q VGND VPWR _316_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
X_247_ _421_/Q VGND VPWR _247_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_28_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_167 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA__218__A1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_280_ _351_/A _311_/B _311_/C VGND VPWR _280_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_14_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input7_A sel[0] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
Xclkbuf_1_1__f_divider2.out clkbuf_0_divider2.out/X VGND VPWR _208_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_401_ _400_/A _458_/Q _457_/Q _459_/Q VGND VPWR _402_/B VGND VPWR sky130_fd_sc_hd__o31ai_1
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_332_ _447_/Q _446_/Q VGND VPWR _332_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_18_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_263_ _451_/Q _452_/Q VGND VPWR _263_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_11_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__281__A2 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_315_ _246_/Y _278_/Y _314_/X VGND VPWR _315_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_246_ _425_/Q VGND VPWR _246_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_11_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__454__SET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_229_ _251_/Y _441_/D _262_/Y VGND VPWR _229_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__450__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_17_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_ext_clk clkbuf_0_ext_clk/X VGND VPWR _205_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_26_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_400_ _400_/A _458_/Q _457_/Q _459_/Q VGND VPWR _400_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_25_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_262_ _447_/Q _448_/Q _446_/Q VGND VPWR _262_/Y VGND VPWR sky130_fd_sc_hd__nor3b_2
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_331_ _250_/Y _263_/Y _330_/X VGND VPWR _331_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_32_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_245_ _431_/Q VGND VPWR _245_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_14_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_314_ _426_/Q _425_/Q _427_/Q VGND VPWR _314_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__309__A _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_228_ _331_/X _329_/B _240_/S VGND VPWR _228_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__311__B _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_0_157 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_330_ _451_/Q _450_/Q _452_/Q VGND VPWR _330_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_261_ _451_/Q _227_/X _388_/S VGND VPWR _451_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_459_ _207_/A1 _459_/D fanout28/X VGND VPWR _459_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_313_ _313_/A _313_/B VGND VPWR _313_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_14_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_244_ _424_/Q VGND VPWR _244_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
XFILLER_20_126 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__309__B _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_227_ _326_/Y _329_/Y _240_/S VGND VPWR _227_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__239__A1 _327_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__311__C _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_28_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A sel2[1] VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_260_ _260_/A VGND VPWR _260_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_157 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_458_ _207_/A1 _458_/D fanout27/X VGND VPWR _458_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_17_143 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_389_ _234_/S _265_/X _236_/X VGND VPWR _389_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_243_ _449_/Q VGND VPWR _243_/Y VGND VPWR sky130_fd_sc_hd__clkinv_4
X_312_ _311_/B _311_/C _351_/A VGND VPWR _313_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_404__9 core_clk VGND VPWR _411_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_20_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_226_ _250_/Y _325_/Y _240_/S VGND VPWR _226_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_209_ _246_/Y _309_/Y _219_/S VGND VPWR _209_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__453__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_457_ _207_/A1 _457_/D fanout27/X VGND VPWR _457_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_388_ _452_/Q _228_/X _388_/S VGND VPWR _452_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_242_ _327_/A _340_/Y _297_/Y VGND VPWR _242_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_311_ _351_/A _311_/B _311_/C VGND VPWR _313_/A VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_14_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_254__7 _403__8/A VGND VPWR _409_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_9_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_ext_clk clkbuf_0_ext_clk/X VGND VPWR _372_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_225_ _439_/Q _324_/Y _292_/Y VGND VPWR _225_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_208_ _208_/A0 _208_/A1 _413_/Q VGND VPWR _208_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA__220__A1 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XPHY_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_17 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_456_ _456_/CLK _456_/D fanout26/X VGND VPWR _456_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_387_ _450_/Q _226_/X _388_/S VGND VPWR _450_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_310_ _426_/Q _425_/Q VGND VPWR _310_/Y VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_14_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_241_ _442_/D _249_/Y _297_/Y VGND VPWR _241_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_439_ _439_/CLK _439_/D fanout29/X VGND VPWR _439_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_9_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_224_ _438_/Q _245_/Y _292_/Y VGND VPWR _224_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_207_ _444_/Q _207_/A1 _264_/Y VGND VPWR _305_/B VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_157 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_386_ _260_/Y _272_/Y _385_/Y VGND VPWR _448_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_455_ _455_/CLK _455_/D fanout28/X VGND VPWR _455_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA_input3_A resetb VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_31_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_240_ _239_/X _327_/A _240_/S VGND VPWR _240_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_369_ _416_/D _432_/Q _431_/Q _433_/Q VGND VPWR _369_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_438_ _206_/A1 _438_/D fanout29/X VGND VPWR _438_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_13_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_223_ _222_/X _351_/A _223_/S VGND VPWR _223_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_206_ _206_/A0 _206_/A1 _413_/Q VGND VPWR _206_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__434__D _434_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_385_ _234_/S _385_/B _448_/Q VGND VPWR _385_/Y VGND VPWR sky130_fd_sc_hd__nand3b_1
X_454_ _455_/CLK _454_/D fanout28/X VGND VPWR _454_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_368_ _225_/X _432_/Q _416_/D VGND VPWR _432_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_437_ _206_/A1 _437_/D fanout29/X VGND VPWR _437_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_299_ _454_/Q _455_/Q VGND VPWR _299_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_12_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_222_ _323_/Y _351_/A _295_/Y VGND VPWR _222_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_102 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_205_ _205_/A0 _415_/Q _413_/D VGND VPWR _205_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_pll_clk90 pll_clk90 VGND VPWR clkbuf_0_pll_clk90/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_18_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__214__A1 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_25_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_51 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_384_ _258_/Y _272_/Y _383_/Y VGND VPWR _446_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
X_453_ _455_/CLK _453_/D fanout28/X VGND VPWR _453_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_16_170 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_22_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_367_ _224_/X _431_/Q _416_/D VGND VPWR _431_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__279__B _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_436_ _439_/CLK _436_/D fanout29/X VGND VPWR _439_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_298_ _240_/S _298_/B VGND VPWR _298_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_3_30 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_221_ _220_/X _311_/B _223_/S VGND VPWR _221_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_419_ _204_/A1 _419_/D _372_/S VGND VPWR _419_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_5_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_204_ _419_/Q _204_/A1 _279_/Y VGND VPWR _301_/B VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f_net10 clkbuf_0_net10/X VGND VPWR _403__8/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_383_ _234_/S _385_/B _446_/Q VGND VPWR _383_/Y VGND VPWR sky130_fd_sc_hd__nand3b_1
X_452_ _455_/CLK _452_/D fanout28/X VGND VPWR _452_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_31_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_297_ _457_/Q _373_/C VGND VPWR _297_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_435_ _439_/CLK _435_/D _372_/S VGND VPWR _438_/D VGND VPWR sky130_fd_sc_hd__dfstp_1
X_366_ _219_/S _365_/Y _293_/Y _223_/X VGND VPWR _430_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_1
XANTENNA__280__B1 _311_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_3_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input1_A ext_clk_sel VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_220_ _320_/Y _311_/B _295_/Y VGND VPWR _220_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_6_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_418_ _204_/A1 _439_/Q VGND VPWR _418_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_349_ _417_/Q _438_/Q VGND VPWR _353_/B VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_23_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_203_ _298_/Y _240_/S _268_/Y VGND VPWR _388_/S VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_382_ _445_/Q _265_/X _378_/Y _381_/Y VGND VPWR _445_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_451_ _451_/CLK _451_/D fanout28/X VGND VPWR _451_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_408__3 _455_/CLK VGND VPWR _451_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
X_296_ _458_/Q _459_/Q VGND VPWR _373_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_434_ _206_/A1 _434_/D _372_/S VGND VPWR _437_/D VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_13_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_365_ _365_/A _430_/Q VGND VPWR _365_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_9_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_279_ _439_/Q _311_/B VGND VPWR _279_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_417_ _204_/A1 _438_/Q VGND VPWR _417_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_348_ _438_/Q _417_/Q VGND VPWR _353_/A VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_5_160 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_202_ _293_/Y _219_/S _283_/Y VGND VPWR _360_/S VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_381_ _379_/Y _380_/X _265_/X VGND VPWR _381_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_450_ _455_/CLK _450_/D fanout28/X VGND VPWR _450_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_433_ _204_/A1 _433_/D _372_/S VGND VPWR _433_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_26_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__280__A2 _311_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_364_ _219_/S _363_/Y _293_/Y _221_/X VGND VPWR _429_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_295_ _429_/Q _430_/Q _295_/C VGND VPWR _295_/Y VGND VPWR sky130_fd_sc_hd__nor3_2
X_347_ _347_/A _347_/B VGND VPWR _419_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XANTENNA__459__RESET_B fanout28/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_416_ _204_/A1 _416_/D VGND VPWR _416_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_278_ _426_/Q _427_/Q VGND VPWR _278_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_5_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_405__5 _456_/CLK VGND VPWR _424_/CLK VGND VPWR sky130_fd_sc_hd__inv_4
XFILLER_29_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_380_ _465_/Q _443_/Q VGND VPWR _380_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_16_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
.ends

.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VPWR Q Q_N VNB VPB
X0 a_788_47# a_942_21# a_648_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR RESET_B a_942_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_942_21# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1429_21# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_474_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X8 a_1545_47# a_942_21# a_1429_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR a_1429_21# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_582_47# a_193_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X11 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_648_21# a_474_413# a_788_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 a_1341_413# a_193_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1663_329# a_1255_47# a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1160_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1255_47# a_27_47# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_648_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_788_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q_N a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND RESET_B a_942_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR a_942_21# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 a_558_413# a_27_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND a_648_21# a_582_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_892_329# a_474_413# a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 VGND a_1429_21# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 a_474_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_1364_47# a_27_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X32 a_1255_47# a_193_47# a_1160_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X33 Q_N a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 a_1545_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 VPWR a_648_21# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 a_1113_329# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 a_1429_21# a_1255_47# a_1545_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_8 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt spare_logic_block spare_xfq[0] spare_xfq[1] spare_xfqn[0] spare_xfqn[1] spare_xi[0]
+ spare_xi[1] spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0]
+ spare_xna[1] spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12]
+ spare_xz[13] spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19]
+ spare_xz[1] spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25]
+ spare_xz[26] spare_xz[2] spare_xz[3] spare_xz[4] spare_xz[5] spare_xz[6] spare_xz[7]
+ spare_xz[8] spare_xz[9] vccd vssd
XFILLER_0_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[8\] vssd vssd vccd vccd spare_logic_const\[8\]/HI spare_xz[8]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_nor\[0\] spare_xz[9] spare_xz[11] vssd vccd spare_xno[0] vssd vccd sky130_fd_sc_hd__nor2_2
XFILLER_0_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[22\] vssd vssd vccd vccd spare_logic_const\[22\]/HI spare_xz[22]
+ sky130_fd_sc_hd__conb_1
XFILLER_3_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[15\] vssd vssd vccd vccd spare_logic_const\[15\]/HI spare_xz[15]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[6\] vssd vssd vccd vccd spare_logic_const\[6\]/HI spare_xz[6]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[20\] vssd vssd vccd vccd spare_logic_const\[20\]/HI spare_xz[20]
+ sky130_fd_sc_hd__conb_1
XFILLER_9_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[13\] vssd vssd vccd vccd spare_logic_const\[13\]/HI spare_xz[13]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[4\] vssd vssd vccd vccd spare_logic_const\[4\]/HI spare_xz[4]
+ sky130_fd_sc_hd__conb_1
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_flop\[0\] spare_xz[21] spare_xz[19] spare_xz[25] spare_xz[23] vssd vccd
+ spare_xfq[0] spare_xfqn[0] vssd vccd sky130_fd_sc_hd__dfbbp_1
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_mux\[1\] spare_xz[14] spare_xz[16] spare_xz[18] vssd vccd spare_xmx[1]
+ vssd vccd sky130_fd_sc_hd__mux2_2
Xspare_logic_const\[11\] vssd vssd vccd vccd spare_logic_const\[11\]/HI spare_xz[11]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[2\] vssd vssd vccd vccd spare_logic_const\[2\]/HI spare_xz[2]
+ sky130_fd_sc_hd__conb_1
XFILLER_1_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[3\] spare_xz[3] vssd vccd spare_xi[3] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[0\] vssd vssd vccd vccd spare_logic_const\[0\]/HI spare_xz[0]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[1\] spare_xz[1] vssd vccd spare_xi[1] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_46 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[25\] vssd vssd vccd vccd spare_logic_const\[25\]/HI spare_xz[25]
+ sky130_fd_sc_hd__conb_1
Xspare_logic_nand\[1\] spare_xz[6] spare_xz[8] vssd vccd spare_xna[1] vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_1_38 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[18\] vssd vssd vccd vccd spare_logic_const\[18\]/HI spare_xz[18]
+ sky130_fd_sc_hd__conb_1
XFILLER_10_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[9\] vssd vssd vccd vccd spare_logic_const\[9\]/HI spare_xz[9]
+ sky130_fd_sc_hd__conb_1
XFILLER_8_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_nor\[1\] spare_xz[10] spare_xz[12] vssd vccd spare_xno[1] vssd vccd sky130_fd_sc_hd__nor2_2
XFILLER_7_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[23\] vssd vssd vccd vccd spare_logic_const\[23\]/HI spare_xz[23]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[16\] vssd vssd vccd vccd spare_logic_const\[16\]/HI spare_xz[16]
+ sky130_fd_sc_hd__conb_1
XFILLER_2_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_const\[7\] vssd vssd vccd vccd spare_logic_const\[7\]/HI spare_xz[7]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_biginv spare_xz[4] vssd vccd spare_xib vssd vccd sky130_fd_sc_hd__inv_8
XFILLER_8_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[21\] vssd vssd vccd vccd spare_logic_const\[21\]/HI spare_xz[21]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[14\] vssd vssd vccd vccd spare_logic_const\[14\]/HI spare_xz[14]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_43 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[5\] vssd vssd vccd vccd spare_logic_const\[5\]/HI spare_xz[5]
+ sky130_fd_sc_hd__conb_1
XFILLER_4_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_flop\[1\] spare_xz[22] spare_xz[20] spare_xz[26] spare_xz[24] vssd vccd
+ spare_xfq[1] spare_xfqn[1] vssd vccd sky130_fd_sc_hd__dfbbp_1
XFILLER_0_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[12\] vssd vssd vccd vccd spare_logic_const\[12\]/HI spare_xz[12]
+ sky130_fd_sc_hd__conb_1
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[3\] vssd vssd vccd vccd spare_logic_const\[3\]/HI spare_xz[3]
+ sky130_fd_sc_hd__conb_1
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_mux\[0\] spare_xz[13] spare_xz[15] spare_xz[17] vssd vccd spare_xmx[0]
+ vssd vccd sky130_fd_sc_hd__mux2_2
Xspare_logic_const\[10\] vssd vssd vccd vccd spare_logic_const\[10\]/HI spare_xz[10]
+ sky130_fd_sc_hd__conb_1
XFILLER_11_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[1\] vssd vssd vccd vccd spare_logic_const\[1\]/HI spare_xz[1]
+ sky130_fd_sc_hd__conb_1
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[2\] spare_xz[2] vssd vccd spare_xi[2] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_8_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[26\] vssd vssd vccd vccd spare_logic_const\[26\]/HI spare_xz[26]
+ sky130_fd_sc_hd__conb_1
XFILLER_5_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
Xspare_logic_const\[19\] vssd vssd vccd vccd spare_logic_const\[19\]/HI spare_xz[19]
+ sky130_fd_sc_hd__conb_1
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xspare_logic_inv\[0\] spare_xz[0] vssd vccd spare_xi[0] vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_0_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_const\[24\] vssd vssd vccd vccd spare_logic_const\[24\]/HI spare_xz[24]
+ sky130_fd_sc_hd__conb_1
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xspare_logic_nand\[0\] spare_xz[5] spare_xz[7] vssd vccd spare_xna[0] vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_3_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xspare_logic_const\[17\] vssd vssd vccd vccd spare_logic_const\[17\]/HI spare_xz[17]
+ sky130_fd_sc_hd__conb_1
XFILLER_6_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
.ends

.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VPWR VGND
Xmask_rev_value\[1\] VGND VGND VPWR VPWR mask_rev_value\[1\]/HI mask_rev[1] sky130_fd_sc_hd__conb_1
XFILLER_6_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[30\] VGND VGND VPWR VPWR mask_rev_value\[30\]/HI mask_rev[30] sky130_fd_sc_hd__conb_1
XFILLER_0_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[23\] VGND VGND VPWR VPWR mask_rev_value\[23\]/HI mask_rev[23] sky130_fd_sc_hd__conb_1
XFILLER_0_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[16\] VGND VGND VPWR VPWR mask_rev_value\[16\]/HI mask_rev[16] sky130_fd_sc_hd__conb_1
XFILLER_0_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[21\] VGND VGND VPWR VPWR mask_rev_value\[21\]/HI mask_rev[21] sky130_fd_sc_hd__conb_1
XFILLER_3_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[14\] VGND VGND VPWR VPWR mask_rev_value\[14\]/HI mask_rev[14] sky130_fd_sc_hd__conb_1
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[8\] VGND VGND VPWR VPWR mask_rev_value\[8\]/HI mask_rev[8] sky130_fd_sc_hd__conb_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[12\] VGND VGND VPWR VPWR mask_rev_value\[12\]/HI mask_rev[12] sky130_fd_sc_hd__conb_1
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[6\] VGND VGND VPWR VPWR mask_rev_value\[6\]/HI mask_rev[6] sky130_fd_sc_hd__conb_1
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[28\] VGND VGND VPWR VPWR mask_rev_value\[28\]/HI mask_rev[28] sky130_fd_sc_hd__conb_1
XFILLER_8_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[10\] VGND VGND VPWR VPWR mask_rev_value\[10\]/HI mask_rev[10] sky130_fd_sc_hd__conb_1
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[4\] VGND VGND VPWR VPWR mask_rev_value\[4\]/HI mask_rev[4] sky130_fd_sc_hd__conb_1
XFILLER_7_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[26\] VGND VGND VPWR VPWR mask_rev_value\[26\]/HI mask_rev[26] sky130_fd_sc_hd__conb_1
XFILLER_4_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[19\] VGND VGND VPWR VPWR mask_rev_value\[19\]/HI mask_rev[19] sky130_fd_sc_hd__conb_1
XFILLER_7_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[2\] VGND VGND VPWR VPWR mask_rev_value\[2\]/HI mask_rev[2] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[31\] VGND VGND VPWR VPWR mask_rev_value\[31\]/HI mask_rev[31] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[24\] VGND VGND VPWR VPWR mask_rev_value\[24\]/HI mask_rev[24] sky130_fd_sc_hd__conb_1
XFILLER_5_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[17\] VGND VGND VPWR VPWR mask_rev_value\[17\]/HI mask_rev[17] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[0\] VGND VGND VPWR VPWR mask_rev_value\[0\]/HI mask_rev[11] sky130_fd_sc_hd__conb_1
XFILLER_5_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[22\] VGND VGND VPWR VPWR mask_rev_value\[22\]/HI mask_rev[22] sky130_fd_sc_hd__conb_1
XFILLER_2_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[15\] VGND VGND VPWR VPWR mask_rev_value\[15\]/HI mask_rev[15] sky130_fd_sc_hd__conb_1
XFILLER_2_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[9\] VGND VGND VPWR VPWR mask_rev_value\[9\]/HI mask_rev[9] sky130_fd_sc_hd__conb_1
XFILLER_8_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[20\] VGND VGND VPWR VPWR mask_rev_value\[20\]/HI mask_rev[20] sky130_fd_sc_hd__conb_1
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[13\] VGND VGND VPWR VPWR mask_rev_value\[13\]/HI mask_rev[13] sky130_fd_sc_hd__conb_1
XFILLER_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[7\] VGND VGND VPWR VPWR mask_rev_value\[7\]/HI mask_rev[7] sky130_fd_sc_hd__conb_1
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[29\] VGND VGND VPWR VPWR mask_rev_value\[29\]/HI mask_rev[29] sky130_fd_sc_hd__conb_1
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[11\] VGND VGND VPWR VPWR mask_rev_value\[11\]/HI mask_rev[0] sky130_fd_sc_hd__conb_1
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[5\] VGND VGND VPWR VPWR mask_rev_value\[5\]/HI mask_rev[5] sky130_fd_sc_hd__conb_1
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[27\] VGND VGND VPWR VPWR mask_rev_value\[27\]/HI mask_rev[27] sky130_fd_sc_hd__conb_1
XFILLER_6_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[3\] VGND VGND VPWR VPWR mask_rev_value\[3\]/HI mask_rev[3] sky130_fd_sc_hd__conb_1
XFILLER_6_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[25\] VGND VGND VPWR VPWR mask_rev_value\[25\]/HI mask_rev[25] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[18\] VGND VGND VPWR VPWR mask_rev_value\[18\]/HI mask_rev[18] sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt gpio_signal_buffering_alt mgmt_io_in_unbuf[6] mgmt_io_out_buf[6] mgmt_io_in_unbuf[5]
+ mgmt_io_in_unbuf[4] mgmt_io_in_unbuf[3] mgmt_io_in_unbuf[2] mgmt_io_in_unbuf[1]
+ mgmt_io_in_unbuf[0] mgmt_io_out_buf[0] mgmt_io_out_buf[1] mgmt_io_out_buf[2] mgmt_io_out_buf[3]
+ mgmt_io_out_buf[4] mgmt_io_out_buf[5] mgmt_io_out_unbuf[0] mgmt_io_out_unbuf[1]
+ mgmt_io_out_unbuf[2] mgmt_io_out_unbuf[3] mgmt_io_out_unbuf[4] mgmt_io_out_unbuf[5]
+ mgmt_io_out_unbuf[6] mgmt_io_in_buf[6] mgmt_io_in_buf[5] mgmt_io_in_buf[4] mgmt_io_in_buf[3]
+ mgmt_io_in_buf[2] mgmt_io_in_buf[1] mgmt_io_in_buf[0] mgmt_io_out_buf[10] mgmt_io_out_buf[11]
+ mgmt_io_in_unbuf[11] mgmt_io_in_unbuf[10] mgmt_io_out_buf[12] mgmt_io_out_buf[13]
+ mgmt_io_out_buf[14] mgmt_io_out_buf[15] mgmt_io_in_unbuf[15] mgmt_io_in_unbuf[14]
+ mgmt_io_in_unbuf[13] mgmt_io_in_unbuf[12] mgmt_io_out_buf[16] mgmt_io_out_buf[17]
+ mgmt_io_out_buf[18] mgmt_io_out_buf[19] mgmt_io_in_unbuf[19] mgmt_io_in_unbuf[18]
+ mgmt_io_in_unbuf[17] mgmt_io_in_unbuf[16] mgmt_io_oeb_buf[0] mgmt_io_oeb_buf[1]
+ mgmt_io_oeb_buf[2] mgmt_io_oeb_unbuf[2] mgmt_io_oeb_unbuf[1] mgmt_io_oeb_unbuf[0]
+ mgmt_io_in_buf[19] mgmt_io_in_buf[18] mgmt_io_in_buf[17] mgmt_io_in_buf[16] mgmt_io_out_unbuf[16]
+ mgmt_io_out_unbuf[17] mgmt_io_out_unbuf[18] mgmt_io_out_unbuf[19] mgmt_io_out_unbuf[15]
+ mgmt_io_out_unbuf[14] mgmt_io_out_unbuf[13] mgmt_io_out_unbuf[12] mgmt_io_out_unbuf[11]
+ mgmt_io_out_unbuf[10] mgmt_io_out_unbuf[9] mgmt_io_out_unbuf[8] mgmt_io_out_unbuf[7]
+ mgmt_io_in_buf[7] mgmt_io_in_buf[8] mgmt_io_in_buf[9] mgmt_io_in_buf[10] mgmt_io_in_buf[11]
+ mgmt_io_in_buf[12] mgmt_io_in_buf[13] mgmt_io_in_buf[14] mgmt_io_in_buf[15] vccd
+ mgmt_io_out_buf[9] mgmt_io_in_unbuf[9] mgmt_io_out_buf[8] mgmt_io_in_unbuf[8] mgmt_io_out_buf[7]
+ mgmt_io_in_unbuf[7] vssd
Xsky130_fd_sc_hd__buf_8_1 sky130_fd_sc_hd__buf_8_1/A vssd vccd sky130_fd_sc_hd__buf_8_1/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_2 mgmt_io_in_unbuf[16] vssd vccd sky130_fd_sc_hd__buf_8_2/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_3 sky130_fd_sc_hd__buf_8_3/A vssd vccd mgmt_io_out_buf[17]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_4 mgmt_io_in_unbuf[18] vssd vccd sky130_fd_sc_hd__buf_8_4/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_5 sky130_fd_sc_hd__buf_8_5/A vssd vccd mgmt_io_out_buf[19]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_6 mgmt_io_in_unbuf[19] vssd vccd sky130_fd_sc_hd__buf_8_6/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_7 sky130_fd_sc_hd__buf_8_7/A vssd vccd mgmt_io_oeb_buf[0]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_8 sky130_fd_sc_hd__buf_8_8/A vssd vccd mgmt_io_oeb_buf[1]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_0 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_9 sky130_fd_sc_hd__buf_8_9/A vssd vccd mgmt_io_oeb_buf[2]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_1 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_2 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_50 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_4 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_90 sky130_fd_sc_hd__buf_8_90/A vssd vccd mgmt_io_in_buf[14]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_40 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_51 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_5 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_170 sky130_fd_sc_hd__buf_8_170/A vssd vccd mgmt_io_out_buf[7]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_91 mgmt_io_out_unbuf[13] vssd vccd sky130_fd_sc_hd__buf_8_91/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_80 sky130_fd_sc_hd__buf_8_80/A vssd vccd sky130_fd_sc_hd__buf_8_90/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_6 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_30 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_52 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_171 mgmt_io_in_unbuf[7] vssd vccd sky130_fd_sc_hd__buf_8_171/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_20 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_31 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_42 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_92 mgmt_io_out_unbuf[12] vssd vccd sky130_fd_sc_hd__buf_8_92/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_81 sky130_fd_sc_hd__buf_8_91/X vssd vccd sky130_fd_sc_hd__buf_8_81/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_7 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_70 sky130_fd_sc_hd__buf_8_70/A vssd vccd sky130_fd_sc_hd__buf_8_70/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_172 mgmt_io_in_unbuf[8] vssd vccd sky130_fd_sc_hd__buf_8_172/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_93 sky130_fd_sc_hd__buf_8_93/A vssd vccd mgmt_io_in_buf[13]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_82 sky130_fd_sc_hd__buf_8_82/A vssd vccd sky130_fd_sc_hd__buf_8_89/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_8 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_10 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_21 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_32 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_43 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_54 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_71 sky130_fd_sc_hd__buf_8_71/A vssd vccd sky130_fd_sc_hd__buf_8_71/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_173 sky130_fd_sc_hd__buf_8_173/A vssd vccd mgmt_io_out_buf[8]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_140 sky130_fd_sc_hd__buf_8_71/X vssd vccd sky130_fd_sc_hd__buf_8_173/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_11 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_22 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_33 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_44 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_55 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_94 mgmt_io_out_unbuf[11] vssd vccd sky130_fd_sc_hd__buf_8_94/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_83 sky130_fd_sc_hd__buf_8_88/X vssd vccd sky130_fd_sc_hd__buf_8_83/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_9 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_50 mgmt_io_out_unbuf[3] vssd vccd mgmt_io_out_buf[3] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_72 sky130_fd_sc_hd__buf_8_72/A vssd vccd sky130_fd_sc_hd__buf_8_97/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_141 sky130_fd_sc_hd__buf_8_172/X vssd vccd sky130_fd_sc_hd__buf_8_68/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_130 mgmt_io_in_unbuf[14] vssd vccd sky130_fd_sc_hd__buf_8_80/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_174 sky130_fd_sc_hd__buf_8_174/A vssd vccd mgmt_io_out_buf[9]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_95 sky130_fd_sc_hd__buf_8_95/A vssd vccd mgmt_io_in_buf[12]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_84 sky130_fd_sc_hd__buf_8_84/A vssd vccd mgmt_io_out_buf[18]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_12 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_23 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_34 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_45 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_56 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_51 mgmt_io_in_unbuf[3] vssd vccd mgmt_io_in_buf[3] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_73 sky130_fd_sc_hd__buf_8_99/X vssd vccd sky130_fd_sc_hd__buf_8_73/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_175 mgmt_io_in_unbuf[9] vssd vccd sky130_fd_sc_hd__buf_8_175/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_142 sky130_fd_sc_hd__buf_8_73/X vssd vccd sky130_fd_sc_hd__buf_8_174/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_131 sky130_fd_sc_hd__buf_8_83/X vssd vccd mgmt_io_out_buf[14]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_120 mgmt_io_out_unbuf[18] vssd vccd sky130_fd_sc_hd__buf_8_84/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_13 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_24 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_35 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_46 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_96 sky130_fd_sc_hd__buf_8_96/A vssd vccd mgmt_io_in_buf[11]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_85 mgmt_io_in_unbuf[17] vssd vccd sky130_fd_sc_hd__buf_8_85/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_52 mgmt_io_out_unbuf[4] vssd vccd mgmt_io_out_buf[4] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_74 sky130_fd_sc_hd__buf_8_74/A vssd vccd sky130_fd_sc_hd__buf_8_96/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_176 sky130_fd_sc_hd__buf_8_176/A vssd vccd mgmt_io_out_buf[10]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_143 sky130_fd_sc_hd__buf_8_175/X vssd vccd sky130_fd_sc_hd__buf_8_70/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_132 mgmt_io_in_unbuf[13] vssd vccd sky130_fd_sc_hd__buf_8_79/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_121 sky130_fd_sc_hd__buf_8_85/X vssd vccd mgmt_io_in_buf[17]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_97 sky130_fd_sc_hd__buf_8_97/A vssd vccd mgmt_io_in_buf[10]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_86 mgmt_io_out_unbuf[15] vssd vccd sky130_fd_sc_hd__buf_8_1/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_14 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_25 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_36 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_47 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_58 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_53 mgmt_io_in_unbuf[4] vssd vccd mgmt_io_in_buf[4] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_75 sky130_fd_sc_hd__buf_8_98/X vssd vccd sky130_fd_sc_hd__buf_8_75/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_177 mgmt_io_in_unbuf[10] vssd vccd sky130_fd_sc_hd__buf_8_177/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_133 sky130_fd_sc_hd__buf_8_81/X vssd vccd mgmt_io_out_buf[13]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_122 sky130_fd_sc_hd__buf_8_4/X vssd vccd mgmt_io_in_buf[18]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_100 sky130_fd_sc_hd__buf_8_70/X vssd vccd mgmt_io_in_buf[9]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_26 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_37 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_48 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_59 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_98 mgmt_io_out_unbuf[10] vssd vccd sky130_fd_sc_hd__buf_8_98/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_76 sky130_fd_sc_hd__buf_8_76/A vssd vccd sky130_fd_sc_hd__buf_8_95/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_178 sky130_fd_sc_hd__buf_8_178/A vssd vccd mgmt_io_out_buf[11]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_134 sky130_fd_sc_hd__buf_8_177/X vssd vccd sky130_fd_sc_hd__buf_8_72/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_123 mgmt_io_out_unbuf[19] vssd vccd sky130_fd_sc_hd__buf_8_5/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_101 sky130_fd_sc_hd__buf_8_68/X vssd vccd mgmt_io_in_buf[8]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_99 mgmt_io_out_unbuf[9] vssd vccd sky130_fd_sc_hd__buf_8_99/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_88 mgmt_io_out_unbuf[14] vssd vccd sky130_fd_sc_hd__buf_8_88/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_77 sky130_fd_sc_hd__buf_8_94/X vssd vccd sky130_fd_sc_hd__buf_8_77/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_16 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_38 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_49 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_55 sky130_fd_sc_hd__buf_8_55/A vssd vccd mgmt_io_out_buf[16]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_179 mgmt_io_in_unbuf[11] vssd vccd sky130_fd_sc_hd__buf_8_179/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_135 sky130_fd_sc_hd__buf_8_75/X vssd vccd sky130_fd_sc_hd__buf_8_176/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_124 sky130_fd_sc_hd__buf_8_6/X vssd vccd mgmt_io_in_buf[19]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_102 sky130_fd_sc_hd__buf_8_67/X vssd vccd mgmt_io_in_buf[7]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_17 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_28 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_89 sky130_fd_sc_hd__buf_8_89/A vssd vccd mgmt_io_in_buf[15]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_78 sky130_fd_sc_hd__buf_8_92/X vssd vccd sky130_fd_sc_hd__buf_8_78/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_12 mgmt_io_out_unbuf[0] vssd vccd mgmt_io_out_buf[0] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_34 mgmt_io_in_unbuf[5] vssd vccd mgmt_io_in_buf[5] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_67 sky130_fd_sc_hd__buf_8_67/A vssd vccd sky130_fd_sc_hd__buf_8_67/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_136 sky130_fd_sc_hd__buf_8_179/X vssd vccd sky130_fd_sc_hd__buf_8_74/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_125 mgmt_io_oeb_unbuf[1] vssd vccd sky130_fd_sc_hd__buf_8_8/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_103 mgmt_io_out_unbuf[8] vssd vccd sky130_fd_sc_hd__buf_8_71/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_18 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_13 mgmt_io_in_unbuf[0] vssd vccd mgmt_io_in_buf[0] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_24 sky130_fd_sc_hd__buf_8_37/X vssd vccd mgmt_io_out_buf[6]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_79 sky130_fd_sc_hd__buf_8_79/A vssd vccd sky130_fd_sc_hd__buf_8_93/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_35 mgmt_io_out_unbuf[5] vssd vccd mgmt_io_out_buf[5] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_46 mgmt_io_in_unbuf[1] vssd vccd mgmt_io_in_buf[1] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_68 sky130_fd_sc_hd__buf_8_68/A vssd vccd sky130_fd_sc_hd__buf_8_68/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_148 sky130_fd_sc_hd__buf_8_69/X vssd vccd sky130_fd_sc_hd__buf_8_170/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_137 sky130_fd_sc_hd__buf_8_77/X vssd vccd sky130_fd_sc_hd__buf_8_178/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_126 mgmt_io_oeb_unbuf[0] vssd vccd sky130_fd_sc_hd__buf_8_7/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_104 mgmt_io_out_unbuf[7] vssd vccd sky130_fd_sc_hd__buf_8_69/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_19 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_25 mgmt_io_in_unbuf[6] vssd vccd sky130_fd_sc_hd__buf_8_36/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_36 sky130_fd_sc_hd__buf_8_36/A vssd vccd mgmt_io_in_buf[6]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_47 mgmt_io_out_unbuf[1] vssd vccd mgmt_io_out_buf[1] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_69 sky130_fd_sc_hd__buf_8_69/A vssd vccd sky130_fd_sc_hd__buf_8_69/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_149 sky130_fd_sc_hd__buf_8_171/X vssd vccd sky130_fd_sc_hd__buf_8_67/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_138 sky130_fd_sc_hd__buf_8_78/X vssd vccd mgmt_io_out_buf[12]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_127 mgmt_io_oeb_unbuf[2] vssd vccd sky130_fd_sc_hd__buf_8_9/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_37 mgmt_io_out_unbuf[6] vssd vccd sky130_fd_sc_hd__buf_8_37/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_48 mgmt_io_out_unbuf[2] vssd vccd mgmt_io_out_buf[2] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_139 mgmt_io_in_unbuf[12] vssd vccd sky130_fd_sc_hd__buf_8_76/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_128 mgmt_io_in_unbuf[15] vssd vccd sky130_fd_sc_hd__buf_8_82/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_117 mgmt_io_out_unbuf[16] vssd vccd sky130_fd_sc_hd__buf_8_55/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_49 mgmt_io_in_unbuf[2] vssd vccd mgmt_io_in_buf[2] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_129 sky130_fd_sc_hd__buf_8_1/X vssd vccd mgmt_io_out_buf[15]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_118 mgmt_io_out_unbuf[17] vssd vccd sky130_fd_sc_hd__buf_8_3/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_119 sky130_fd_sc_hd__buf_8_2/X vssd vccd mgmt_io_in_buf[16]
+ vssd vccd sky130_fd_sc_hd__buf_8
.ends

.subckt sky130_fd_sc_hd__buf_6 A VGND VPWR X VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_4 A B VGND VPWR X VNB VPB
X0 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VPWR X VNB VPB
X0 a_98_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_98_199# a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_56_297# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_56_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_257_47# B a_152_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_56_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_152_47# a_98_199# a_56_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C a_56_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_98_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_56_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND C a_257_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 X a_56_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_4 A B VGND VPWR Y VNB VPB
X0 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_8 A B VGND VPWR Y VNB VPB
X0 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VPWR X VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VPWR X VNB VPB
X0 a_109_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_209_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_296_53# a_109_93# a_209_311# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR C a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_368_53# B a_296_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_209_311# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_209_311# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR a_109_93# a_209_311# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND C a_368_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt mprj2_logic_high HI vccd2 vssd2
XFILLER_0_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_95 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XPHY_0 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_1 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_6
XFILLER_1_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_2 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XPHY_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_209 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_69 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_15 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_181 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_193 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_1_29 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_1_107 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_197 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_153 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_165 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_113 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_169 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_125 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_137 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_81 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
Xinst vssd2 vssd2 vccd2 vccd2 HI inst/LO sky130_fd_sc_hd__conb_1
XFILLER_0_85 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_41 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_109 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
XFILLER_0_97 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd2 vccd2 vssd2 vccd2 sky130_fd_sc_hd__decap_3
.ends

.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[462] HI[46]
+ HI[47] HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57]
+ HI[58] HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79]
+ HI[7] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8]
+ HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1
+ vssd1
Xinsts\[210\] vssd1 vssd1 vccd1 vccd1 HI[210] insts\[210\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[308\] vssd1 vssd1 vccd1 vccd1 HI[308] insts\[308\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[425\] vssd1 vssd1 vccd1 vccd1 HI[425] insts\[425\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[160\] vssd1 vssd1 vccd1 vccd1 HI[160] insts\[160\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_357 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_302 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[258\] vssd1 vssd1 vccd1 vccd1 HI[258] insts\[258\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[40\] vssd1 vssd1 vccd1 vccd1 HI[40] insts\[40\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[375\] vssd1 vssd1 vccd1 vccd1 HI[375] insts\[375\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[88\] vssd1 vssd1 vccd1 vccd1 HI[88] insts\[88\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_165 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[123\] vssd1 vssd1 vccd1 vccd1 HI[123] insts\[123\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[338\] vssd1 vssd1 vccd1 vccd1 HI[338] insts\[338\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[240\] vssd1 vssd1 vccd1 vccd1 HI[240] insts\[240\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[9\] vssd1 vssd1 vccd1 vccd1 HI[9] insts\[9\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[455\] vssd1 vssd1 vccd1 vccd1 HI[455] insts\[455\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[288\] vssd1 vssd1 vccd1 vccd1 HI[288] insts\[288\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[190\] vssd1 vssd1 vccd1 vccd1 HI[190] insts\[190\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[70\] vssd1 vssd1 vccd1 vccd1 HI[70] insts\[70\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[203\] vssd1 vssd1 vccd1 vccd1 HI[203] insts\[203\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_561 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[418\] vssd1 vssd1 vccd1 vccd1 HI[418] insts\[418\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[153\] vssd1 vssd1 vccd1 vccd1 HI[153] insts\[153\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[320\] vssd1 vssd1 vccd1 vccd1 HI[320] insts\[320\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[33\] vssd1 vssd1 vccd1 vccd1 HI[33] insts\[33\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[368\] vssd1 vssd1 vccd1 vccd1 HI[368] insts\[368\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[270\] vssd1 vssd1 vccd1 vccd1 HI[270] insts\[270\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_177 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_486 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[116\] vssd1 vssd1 vccd1 vccd1 HI[116] insts\[116\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[400\] vssd1 vssd1 vccd1 vccd1 HI[400] insts\[400\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[233\] vssd1 vssd1 vccd1 vccd1 HI[233] insts\[233\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[183\] vssd1 vssd1 vccd1 vccd1 HI[183] insts\[183\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[350\] vssd1 vssd1 vccd1 vccd1 HI[350] insts\[350\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[448\] vssd1 vssd1 vccd1 vccd1 HI[448] insts\[448\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_721 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[63\] vssd1 vssd1 vccd1 vccd1 HI[63] insts\[63\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[398\] vssd1 vssd1 vccd1 vccd1 HI[398] insts\[398\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_573 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[146\] vssd1 vssd1 vccd1 vccd1 HI[146] insts\[146\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[313\] vssd1 vssd1 vccd1 vccd1 HI[313] insts\[313\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[26\] vssd1 vssd1 vccd1 vccd1 HI[26] insts\[26\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[430\] vssd1 vssd1 vccd1 vccd1 HI[430] insts\[430\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_189 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[263\] vssd1 vssd1 vccd1 vccd1 HI[263] insts\[263\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[380\] vssd1 vssd1 vccd1 vccd1 HI[380] insts\[380\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[109\] vssd1 vssd1 vccd1 vccd1 HI[109] insts\[109\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[93\] vssd1 vssd1 vccd1 vccd1 HI[93] insts\[93\]/LO sky130_fd_sc_hd__conb_1
XFILLER_3_498 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_80 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[226\] vssd1 vssd1 vccd1 vccd1 HI[226] insts\[226\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[343\] vssd1 vssd1 vccd1 vccd1 HI[343] insts\[343\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[176\] vssd1 vssd1 vccd1 vccd1 HI[176] insts\[176\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[56\] vssd1 vssd1 vccd1 vccd1 HI[56] insts\[56\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[460\] vssd1 vssd1 vccd1 vccd1 HI[460] insts\[460\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[293\] vssd1 vssd1 vccd1 vccd1 HI[293] insts\[293\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_541 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[139\] vssd1 vssd1 vccd1 vccd1 HI[139] insts\[139\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[306\] vssd1 vssd1 vccd1 vccd1 HI[306] insts\[306\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[19\] vssd1 vssd1 vccd1 vccd1 HI[19] insts\[19\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_393 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[423\] vssd1 vssd1 vccd1 vccd1 HI[423] insts\[423\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[256\] vssd1 vssd1 vccd1 vccd1 HI[256] insts\[256\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[373\] vssd1 vssd1 vccd1 vccd1 HI[373] insts\[373\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[86\] vssd1 vssd1 vccd1 vccd1 HI[86] insts\[86\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[121\] vssd1 vssd1 vccd1 vccd1 HI[121] insts\[121\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[219\] vssd1 vssd1 vccd1 vccd1 HI[219] insts\[219\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[336\] vssd1 vssd1 vccd1 vccd1 HI[336] insts\[336\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[169\] vssd1 vssd1 vccd1 vccd1 HI[169] insts\[169\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[49\] vssd1 vssd1 vccd1 vccd1 HI[49] insts\[49\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[286\] vssd1 vssd1 vccd1 vccd1 HI[286] insts\[286\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[7\] vssd1 vssd1 vccd1 vccd1 HI[7] insts\[7\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[453\] vssd1 vssd1 vccd1 vccd1 HI[453] insts\[453\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_597 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[201\] vssd1 vssd1 vccd1 vccd1 HI[201] insts\[201\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[416\] vssd1 vssd1 vccd1 vccd1 HI[416] insts\[416\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[151\] vssd1 vssd1 vccd1 vccd1 HI[151] insts\[151\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[249\] vssd1 vssd1 vccd1 vccd1 HI[249] insts\[249\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_681 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[31\] vssd1 vssd1 vccd1 vccd1 HI[31] insts\[31\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[366\] vssd1 vssd1 vccd1 vccd1 HI[366] insts\[366\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[199\] vssd1 vssd1 vccd1 vccd1 HI[199] insts\[199\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[79\] vssd1 vssd1 vccd1 vccd1 HI[79] insts\[79\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[114\] vssd1 vssd1 vccd1 vccd1 HI[114] insts\[114\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[329\] vssd1 vssd1 vccd1 vccd1 HI[329] insts\[329\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[231\] vssd1 vssd1 vccd1 vccd1 HI[231] insts\[231\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[446\] vssd1 vssd1 vccd1 vccd1 HI[446] insts\[446\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[181\] vssd1 vssd1 vccd1 vccd1 HI[181] insts\[181\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[279\] vssd1 vssd1 vccd1 vccd1 HI[279] insts\[279\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[61\] vssd1 vssd1 vccd1 vccd1 HI[61] insts\[61\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[396\] vssd1 vssd1 vccd1 vccd1 HI[396] insts\[396\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[144\] vssd1 vssd1 vccd1 vccd1 HI[144] insts\[144\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[409\] vssd1 vssd1 vccd1 vccd1 HI[409] insts\[409\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[311\] vssd1 vssd1 vccd1 vccd1 HI[311] insts\[311\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[24\] vssd1 vssd1 vccd1 vccd1 HI[24] insts\[24\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[359\] vssd1 vssd1 vccd1 vccd1 HI[359] insts\[359\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[261\] vssd1 vssd1 vccd1 vccd1 HI[261] insts\[261\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[107\] vssd1 vssd1 vccd1 vccd1 HI[107] insts\[107\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[91\] vssd1 vssd1 vccd1 vccd1 HI[91] insts\[91\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[224\] vssd1 vssd1 vccd1 vccd1 HI[224] insts\[224\]/LO sky130_fd_sc_hd__conb_1
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[439\] vssd1 vssd1 vccd1 vccd1 HI[439] insts\[439\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[174\] vssd1 vssd1 vccd1 vccd1 HI[174] insts\[174\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[341\] vssd1 vssd1 vccd1 vccd1 HI[341] insts\[341\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[54\] vssd1 vssd1 vccd1 vccd1 HI[54] insts\[54\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[389\] vssd1 vssd1 vccd1 vccd1 HI[389] insts\[389\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[291\] vssd1 vssd1 vccd1 vccd1 HI[291] insts\[291\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[137\] vssd1 vssd1 vccd1 vccd1 HI[137] insts\[137\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[304\] vssd1 vssd1 vccd1 vccd1 HI[304] insts\[304\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[17\] vssd1 vssd1 vccd1 vccd1 HI[17] insts\[17\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[421\] vssd1 vssd1 vccd1 vccd1 HI[421] insts\[421\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[254\] vssd1 vssd1 vccd1 vccd1 HI[254] insts\[254\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[371\] vssd1 vssd1 vccd1 vccd1 HI[371] insts\[371\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[84\] vssd1 vssd1 vccd1 vccd1 HI[84] insts\[84\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[217\] vssd1 vssd1 vccd1 vccd1 HI[217] insts\[217\]/LO sky130_fd_sc_hd__conb_1
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[334\] vssd1 vssd1 vccd1 vccd1 HI[334] insts\[334\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[167\] vssd1 vssd1 vccd1 vccd1 HI[167] insts\[167\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[47\] vssd1 vssd1 vccd1 vccd1 HI[47] insts\[47\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_309 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[5\] vssd1 vssd1 vccd1 vccd1 HI[5] insts\[5\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[451\] vssd1 vssd1 vccd1 vccd1 HI[451] insts\[451\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[284\] vssd1 vssd1 vccd1 vccd1 HI[284] insts\[284\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_331 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[247\] vssd1 vssd1 vccd1 vccd1 HI[247] insts\[247\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[414\] vssd1 vssd1 vccd1 vccd1 HI[414] insts\[414\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_470 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_96 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[364\] vssd1 vssd1 vccd1 vccd1 HI[364] insts\[364\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[197\] vssd1 vssd1 vccd1 vccd1 HI[197] insts\[197\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[77\] vssd1 vssd1 vccd1 vccd1 HI[77] insts\[77\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[112\] vssd1 vssd1 vccd1 vccd1 HI[112] insts\[112\]/LO sky130_fd_sc_hd__conb_1
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[327\] vssd1 vssd1 vccd1 vccd1 HI[327] insts\[327\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[444\] vssd1 vssd1 vccd1 vccd1 HI[444] insts\[444\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[277\] vssd1 vssd1 vccd1 vccd1 HI[277] insts\[277\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_343 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[394\] vssd1 vssd1 vccd1 vccd1 HI[394] insts\[394\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_118 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[407\] vssd1 vssd1 vccd1 vccd1 HI[407] insts\[407\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[142\] vssd1 vssd1 vccd1 vccd1 HI[142] insts\[142\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[22\] vssd1 vssd1 vccd1 vccd1 HI[22] insts\[22\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[357\] vssd1 vssd1 vccd1 vccd1 HI[357] insts\[357\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[105\] vssd1 vssd1 vccd1 vccd1 HI[105] insts\[105\]/LO sky130_fd_sc_hd__conb_1
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[222\] vssd1 vssd1 vccd1 vccd1 HI[222] insts\[222\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[437\] vssd1 vssd1 vccd1 vccd1 HI[437] insts\[437\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[172\] vssd1 vssd1 vccd1 vccd1 HI[172] insts\[172\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_355 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[52\] vssd1 vssd1 vccd1 vccd1 HI[52] insts\[52\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[387\] vssd1 vssd1 vccd1 vccd1 HI[387] insts\[387\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_196 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[135\] vssd1 vssd1 vccd1 vccd1 HI[135] insts\[135\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[302\] vssd1 vssd1 vccd1 vccd1 HI[302] insts\[302\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[15\] vssd1 vssd1 vccd1 vccd1 HI[15] insts\[15\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[252\] vssd1 vssd1 vccd1 vccd1 HI[252] insts\[252\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[82\] vssd1 vssd1 vccd1 vccd1 HI[82] insts\[82\]/LO sky130_fd_sc_hd__conb_1
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[215\] vssd1 vssd1 vccd1 vccd1 HI[215] insts\[215\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[165\] vssd1 vssd1 vccd1 vccd1 HI[165] insts\[165\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[332\] vssd1 vssd1 vccd1 vccd1 HI[332] insts\[332\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_301 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_367 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[45\] vssd1 vssd1 vccd1 vccd1 HI[45] insts\[45\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_109 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[3\] vssd1 vssd1 vccd1 vccd1 HI[3] insts\[3\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[282\] vssd1 vssd1 vccd1 vccd1 HI[282] insts\[282\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_142 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[128\] vssd1 vssd1 vccd1 vccd1 HI[128] insts\[128\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[412\] vssd1 vssd1 vccd1 vccd1 HI[412] insts\[412\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[245\] vssd1 vssd1 vccd1 vccd1 HI[245] insts\[245\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[362\] vssd1 vssd1 vccd1 vccd1 HI[362] insts\[362\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[195\] vssd1 vssd1 vccd1 vccd1 HI[195] insts\[195\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[75\] vssd1 vssd1 vccd1 vccd1 HI[75] insts\[75\]/LO sky130_fd_sc_hd__conb_1
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[110\] vssd1 vssd1 vccd1 vccd1 HI[110] insts\[110\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[208\] vssd1 vssd1 vccd1 vccd1 HI[208] insts\[208\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_505 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[158\] vssd1 vssd1 vccd1 vccd1 HI[158] insts\[158\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[325\] vssd1 vssd1 vccd1 vccd1 HI[325] insts\[325\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_379 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[38\] vssd1 vssd1 vccd1 vccd1 HI[38] insts\[38\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[442\] vssd1 vssd1 vccd1 vccd1 HI[442] insts\[442\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[275\] vssd1 vssd1 vccd1 vccd1 HI[275] insts\[275\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_121 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_154 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[392\] vssd1 vssd1 vccd1 vccd1 HI[392] insts\[392\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[405\] vssd1 vssd1 vccd1 vccd1 HI[405] insts\[405\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[140\] vssd1 vssd1 vccd1 vccd1 HI[140] insts\[140\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[238\] vssd1 vssd1 vccd1 vccd1 HI[238] insts\[238\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[20\] vssd1 vssd1 vccd1 vccd1 HI[20] insts\[20\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[355\] vssd1 vssd1 vccd1 vccd1 HI[355] insts\[355\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[188\] vssd1 vssd1 vccd1 vccd1 HI[188] insts\[188\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_709 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[68\] vssd1 vssd1 vccd1 vccd1 HI[68] insts\[68\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_517 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[103\] vssd1 vssd1 vccd1 vccd1 HI[103] insts\[103\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[318\] vssd1 vssd1 vccd1 vccd1 HI[318] insts\[318\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[220\] vssd1 vssd1 vccd1 vccd1 HI[220] insts\[220\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[170\] vssd1 vssd1 vccd1 vccd1 HI[170] insts\[170\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[435\] vssd1 vssd1 vccd1 vccd1 HI[435] insts\[435\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_689 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[268\] vssd1 vssd1 vccd1 vccd1 HI[268] insts\[268\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[50\] vssd1 vssd1 vccd1 vccd1 HI[50] insts\[50\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[385\] vssd1 vssd1 vccd1 vccd1 HI[385] insts\[385\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[98\] vssd1 vssd1 vccd1 vccd1 HI[98] insts\[98\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_442 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_68 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[133\] vssd1 vssd1 vccd1 vccd1 HI[133] insts\[133\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[300\] vssd1 vssd1 vccd1 vccd1 HI[300] insts\[300\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[13\] vssd1 vssd1 vccd1 vccd1 HI[13] insts\[13\]/LO sky130_fd_sc_hd__conb_1
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[348\] vssd1 vssd1 vccd1 vccd1 HI[348] insts\[348\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[250\] vssd1 vssd1 vccd1 vccd1 HI[250] insts\[250\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[298\] vssd1 vssd1 vccd1 vccd1 HI[298] insts\[298\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_529 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[80\] vssd1 vssd1 vccd1 vccd1 HI[80] insts\[80\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[213\] vssd1 vssd1 vccd1 vccd1 HI[213] insts\[213\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_337 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[428\] vssd1 vssd1 vccd1 vccd1 HI[428] insts\[428\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[330\] vssd1 vssd1 vccd1 vccd1 HI[330] insts\[330\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[163\] vssd1 vssd1 vccd1 vccd1 HI[163] insts\[163\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[43\] vssd1 vssd1 vccd1 vccd1 HI[43] insts\[43\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[378\] vssd1 vssd1 vccd1 vccd1 HI[378] insts\[378\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[280\] vssd1 vssd1 vccd1 vccd1 HI[280] insts\[280\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[1\] vssd1 vssd1 vccd1 vccd1 HI[1] insts\[1\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_454 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[126\] vssd1 vssd1 vccd1 vccd1 HI[126] insts\[126\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[410\] vssd1 vssd1 vccd1 vccd1 HI[410] insts\[410\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[243\] vssd1 vssd1 vccd1 vccd1 HI[243] insts\[243\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[458\] vssd1 vssd1 vccd1 vccd1 HI[458] insts\[458\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[360\] vssd1 vssd1 vccd1 vccd1 HI[360] insts\[360\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[193\] vssd1 vssd1 vccd1 vccd1 HI[193] insts\[193\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[73\] vssd1 vssd1 vccd1 vccd1 HI[73] insts\[73\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[206\] vssd1 vssd1 vccd1 vccd1 HI[206] insts\[206\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_669 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[156\] vssd1 vssd1 vccd1 vccd1 HI[156] insts\[156\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[323\] vssd1 vssd1 vccd1 vccd1 HI[323] insts\[323\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[36\] vssd1 vssd1 vccd1 vccd1 HI[36] insts\[36\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[273\] vssd1 vssd1 vccd1 vccd1 HI[273] insts\[273\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[440\] vssd1 vssd1 vccd1 vccd1 HI[440] insts\[440\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_433 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[390\] vssd1 vssd1 vccd1 vccd1 HI[390] insts\[390\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[119\] vssd1 vssd1 vccd1 vccd1 HI[119] insts\[119\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[403\] vssd1 vssd1 vccd1 vccd1 HI[403] insts\[403\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[236\] vssd1 vssd1 vccd1 vccd1 HI[236] insts\[236\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_701 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[353\] vssd1 vssd1 vccd1 vccd1 HI[353] insts\[353\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[186\] vssd1 vssd1 vccd1 vccd1 HI[186] insts\[186\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[66\] vssd1 vssd1 vccd1 vccd1 HI[66] insts\[66\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[101\] vssd1 vssd1 vccd1 vccd1 HI[101] insts\[101\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[149\] vssd1 vssd1 vccd1 vccd1 HI[149] insts\[149\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_637 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[316\] vssd1 vssd1 vccd1 vccd1 HI[316] insts\[316\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[29\] vssd1 vssd1 vccd1 vccd1 HI[29] insts\[29\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[433\] vssd1 vssd1 vccd1 vccd1 HI[433] insts\[433\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[266\] vssd1 vssd1 vccd1 vccd1 HI[266] insts\[266\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[383\] vssd1 vssd1 vccd1 vccd1 HI[383] insts\[383\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[96\] vssd1 vssd1 vccd1 vccd1 HI[96] insts\[96\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_253 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[131\] vssd1 vssd1 vccd1 vccd1 HI[131] insts\[131\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[229\] vssd1 vssd1 vccd1 vccd1 HI[229] insts\[229\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_713 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[11\] vssd1 vssd1 vccd1 vccd1 HI[11] insts\[11\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[346\] vssd1 vssd1 vccd1 vccd1 HI[346] insts\[346\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[179\] vssd1 vssd1 vccd1 vccd1 HI[179] insts\[179\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[59\] vssd1 vssd1 vccd1 vccd1 HI[59] insts\[59\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_307 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[296\] vssd1 vssd1 vccd1 vccd1 HI[296] insts\[296\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[309\] vssd1 vssd1 vccd1 vccd1 HI[309] insts\[309\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[211\] vssd1 vssd1 vccd1 vccd1 HI[211] insts\[211\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[426\] vssd1 vssd1 vccd1 vccd1 HI[426] insts\[426\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[161\] vssd1 vssd1 vccd1 vccd1 HI[161] insts\[161\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[259\] vssd1 vssd1 vccd1 vccd1 HI[259] insts\[259\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[41\] vssd1 vssd1 vccd1 vccd1 HI[41] insts\[41\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_490 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[376\] vssd1 vssd1 vccd1 vccd1 HI[376] insts\[376\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_265 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[89\] vssd1 vssd1 vccd1 vccd1 HI[89] insts\[89\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_60 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[124\] vssd1 vssd1 vccd1 vccd1 HI[124] insts\[124\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_725 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[241\] vssd1 vssd1 vccd1 vccd1 HI[241] insts\[241\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[339\] vssd1 vssd1 vccd1 vccd1 HI[339] insts\[339\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_319 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[456\] vssd1 vssd1 vccd1 vccd1 HI[456] insts\[456\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[289\] vssd1 vssd1 vccd1 vccd1 HI[289] insts\[289\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[191\] vssd1 vssd1 vccd1 vccd1 HI[191] insts\[191\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[71\] vssd1 vssd1 vccd1 vccd1 HI[71] insts\[71\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[204\] vssd1 vssd1 vccd1 vccd1 HI[204] insts\[204\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[419\] vssd1 vssd1 vccd1 vccd1 HI[419] insts\[419\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[154\] vssd1 vssd1 vccd1 vccd1 HI[154] insts\[154\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[321\] vssd1 vssd1 vccd1 vccd1 HI[321] insts\[321\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[34\] vssd1 vssd1 vccd1 vccd1 HI[34] insts\[34\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[369\] vssd1 vssd1 vccd1 vccd1 HI[369] insts\[369\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_277 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[271\] vssd1 vssd1 vccd1 vccd1 HI[271] insts\[271\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_72 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[117\] vssd1 vssd1 vccd1 vccd1 HI[117] insts\[117\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[234\] vssd1 vssd1 vccd1 vccd1 HI[234] insts\[234\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[401\] vssd1 vssd1 vccd1 vccd1 HI[401] insts\[401\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[351\] vssd1 vssd1 vccd1 vccd1 HI[351] insts\[351\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[449\] vssd1 vssd1 vccd1 vccd1 HI[449] insts\[449\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[184\] vssd1 vssd1 vccd1 vccd1 HI[184] insts\[184\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[64\] vssd1 vssd1 vccd1 vccd1 HI[64] insts\[64\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[399\] vssd1 vssd1 vccd1 vccd1 HI[399] insts\[399\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[147\] vssd1 vssd1 vccd1 vccd1 HI[147] insts\[147\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[314\] vssd1 vssd1 vccd1 vccd1 HI[314] insts\[314\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[27\] vssd1 vssd1 vccd1 vccd1 HI[27] insts\[27\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[431\] vssd1 vssd1 vccd1 vccd1 HI[431] insts\[431\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_289 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_245 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[264\] vssd1 vssd1 vccd1 vccd1 HI[264] insts\[264\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[381\] vssd1 vssd1 vccd1 vccd1 HI[381] insts\[381\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[94\] vssd1 vssd1 vccd1 vccd1 HI[94] insts\[94\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[227\] vssd1 vssd1 vccd1 vccd1 HI[227] insts\[227\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[344\] vssd1 vssd1 vccd1 vccd1 HI[344] insts\[344\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[177\] vssd1 vssd1 vccd1 vccd1 HI[177] insts\[177\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[57\] vssd1 vssd1 vccd1 vccd1 HI[57] insts\[57\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[461\] vssd1 vssd1 vccd1 vccd1 HI[461] insts\[461\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[294\] vssd1 vssd1 vccd1 vccd1 HI[294] insts\[294\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[307\] vssd1 vssd1 vccd1 vccd1 HI[307] insts\[307\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_471 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[424\] vssd1 vssd1 vccd1 vccd1 HI[424] insts\[424\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[257\] vssd1 vssd1 vccd1 vccd1 HI[257] insts\[257\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_85 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_511 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[374\] vssd1 vssd1 vccd1 vccd1 HI[374] insts\[374\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[87\] vssd1 vssd1 vccd1 vccd1 HI[87] insts\[87\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[122\] vssd1 vssd1 vccd1 vccd1 HI[122] insts\[122\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[337\] vssd1 vssd1 vccd1 vccd1 HI[337] insts\[337\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_108 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[8\] vssd1 vssd1 vccd1 vccd1 HI[8] insts\[8\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[454\] vssd1 vssd1 vccd1 vccd1 HI[454] insts\[454\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[287\] vssd1 vssd1 vccd1 vccd1 HI[287] insts\[287\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_653 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[202\] vssd1 vssd1 vccd1 vccd1 HI[202] insts\[202\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_461 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[417\] vssd1 vssd1 vccd1 vccd1 HI[417] insts\[417\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[152\] vssd1 vssd1 vccd1 vccd1 HI[152] insts\[152\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_97 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[32\] vssd1 vssd1 vccd1 vccd1 HI[32] insts\[32\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[367\] vssd1 vssd1 vccd1 vccd1 HI[367] insts\[367\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[115\] vssd1 vssd1 vccd1 vccd1 HI[115] insts\[115\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[232\] vssd1 vssd1 vccd1 vccd1 HI[232] insts\[232\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[447\] vssd1 vssd1 vccd1 vccd1 HI[447] insts\[447\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[182\] vssd1 vssd1 vccd1 vccd1 HI[182] insts\[182\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[62\] vssd1 vssd1 vccd1 vccd1 HI[62] insts\[62\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_665 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[397\] vssd1 vssd1 vccd1 vccd1 HI[397] insts\[397\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_484 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[145\] vssd1 vssd1 vccd1 vccd1 HI[145] insts\[145\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[312\] vssd1 vssd1 vccd1 vccd1 HI[312] insts\[312\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[25\] vssd1 vssd1 vccd1 vccd1 HI[25] insts\[25\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_281 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[262\] vssd1 vssd1 vccd1 vccd1 HI[262] insts\[262\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[108\] vssd1 vssd1 vccd1 vccd1 HI[108] insts\[108\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[92\] vssd1 vssd1 vccd1 vccd1 HI[92] insts\[92\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[225\] vssd1 vssd1 vccd1 vccd1 HI[225] insts\[225\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[342\] vssd1 vssd1 vccd1 vccd1 HI[342] insts\[342\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[175\] vssd1 vssd1 vccd1 vccd1 HI[175] insts\[175\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[55\] vssd1 vssd1 vccd1 vccd1 HI[55] insts\[55\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[292\] vssd1 vssd1 vccd1 vccd1 HI[292] insts\[292\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_441 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[138\] vssd1 vssd1 vccd1 vccd1 HI[138] insts\[138\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[305\] vssd1 vssd1 vccd1 vccd1 HI[305] insts\[305\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[18\] vssd1 vssd1 vccd1 vccd1 HI[18] insts\[18\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_293 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[422\] vssd1 vssd1 vccd1 vccd1 HI[422] insts\[422\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[255\] vssd1 vssd1 vccd1 vccd1 HI[255] insts\[255\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[372\] vssd1 vssd1 vccd1 vccd1 HI[372] insts\[372\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[85\] vssd1 vssd1 vccd1 vccd1 HI[85] insts\[85\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[120\] vssd1 vssd1 vccd1 vccd1 HI[120] insts\[120\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[218\] vssd1 vssd1 vccd1 vccd1 HI[218] insts\[218\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[335\] vssd1 vssd1 vccd1 vccd1 HI[335] insts\[335\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[168\] vssd1 vssd1 vccd1 vccd1 HI[168] insts\[168\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[48\] vssd1 vssd1 vccd1 vccd1 HI[48] insts\[48\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[6\] vssd1 vssd1 vccd1 vccd1 HI[6] insts\[6\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[452\] vssd1 vssd1 vccd1 vccd1 HI[452] insts\[452\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[285\] vssd1 vssd1 vccd1 vccd1 HI[285] insts\[285\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[200\] vssd1 vssd1 vccd1 vccd1 HI[200] insts\[200\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_261 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[415\] vssd1 vssd1 vccd1 vccd1 HI[415] insts\[415\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[150\] vssd1 vssd1 vccd1 vccd1 HI[150] insts\[150\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[248\] vssd1 vssd1 vccd1 vccd1 HI[248] insts\[248\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_581 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[30\] vssd1 vssd1 vccd1 vccd1 HI[30] insts\[30\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[365\] vssd1 vssd1 vccd1 vccd1 HI[365] insts\[365\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[198\] vssd1 vssd1 vccd1 vccd1 HI[198] insts\[198\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[78\] vssd1 vssd1 vccd1 vccd1 HI[78] insts\[78\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[113\] vssd1 vssd1 vccd1 vccd1 HI[113] insts\[113\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[230\] vssd1 vssd1 vccd1 vccd1 HI[230] insts\[230\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[328\] vssd1 vssd1 vccd1 vccd1 HI[328] insts\[328\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[445\] vssd1 vssd1 vccd1 vccd1 HI[445] insts\[445\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[278\] vssd1 vssd1 vccd1 vccd1 HI[278] insts\[278\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[180\] vssd1 vssd1 vccd1 vccd1 HI[180] insts\[180\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[60\] vssd1 vssd1 vccd1 vccd1 HI[60] insts\[60\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[395\] vssd1 vssd1 vccd1 vccd1 HI[395] insts\[395\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_273 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[408\] vssd1 vssd1 vccd1 vccd1 HI[408] insts\[408\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[143\] vssd1 vssd1 vccd1 vccd1 HI[143] insts\[143\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[310\] vssd1 vssd1 vccd1 vccd1 HI[310] insts\[310\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[23\] vssd1 vssd1 vccd1 vccd1 HI[23] insts\[23\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[358\] vssd1 vssd1 vccd1 vccd1 HI[358] insts\[358\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[260\] vssd1 vssd1 vccd1 vccd1 HI[260] insts\[260\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[106\] vssd1 vssd1 vccd1 vccd1 HI[106] insts\[106\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[90\] vssd1 vssd1 vccd1 vccd1 HI[90] insts\[90\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[223\] vssd1 vssd1 vccd1 vccd1 HI[223] insts\[223\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[438\] vssd1 vssd1 vccd1 vccd1 HI[438] insts\[438\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[340\] vssd1 vssd1 vccd1 vccd1 HI[340] insts\[340\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[173\] vssd1 vssd1 vccd1 vccd1 HI[173] insts\[173\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[53\] vssd1 vssd1 vccd1 vccd1 HI[53] insts\[53\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[388\] vssd1 vssd1 vccd1 vccd1 HI[388] insts\[388\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[290\] vssd1 vssd1 vccd1 vccd1 HI[290] insts\[290\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_230 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[136\] vssd1 vssd1 vccd1 vccd1 HI[136] insts\[136\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[303\] vssd1 vssd1 vccd1 vccd1 HI[303] insts\[303\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[16\] vssd1 vssd1 vccd1 vccd1 HI[16] insts\[16\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[420\] vssd1 vssd1 vccd1 vccd1 HI[420] insts\[420\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[253\] vssd1 vssd1 vccd1 vccd1 HI[253] insts\[253\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[370\] vssd1 vssd1 vccd1 vccd1 HI[370] insts\[370\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[83\] vssd1 vssd1 vccd1 vccd1 HI[83] insts\[83\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[216\] vssd1 vssd1 vccd1 vccd1 HI[216] insts\[216\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[166\] vssd1 vssd1 vccd1 vccd1 HI[166] insts\[166\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[333\] vssd1 vssd1 vccd1 vccd1 HI[333] insts\[333\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[46\] vssd1 vssd1 vccd1 vccd1 HI[46] insts\[46\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[450\] vssd1 vssd1 vccd1 vccd1 HI[450] insts\[450\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_209 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[283\] vssd1 vssd1 vccd1 vccd1 HI[283] insts\[283\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[4\] vssd1 vssd1 vccd1 vccd1 HI[4] insts\[4\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_710 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[129\] vssd1 vssd1 vccd1 vccd1 HI[129] insts\[129\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[413\] vssd1 vssd1 vccd1 vccd1 HI[413] insts\[413\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[246\] vssd1 vssd1 vccd1 vccd1 HI[246] insts\[246\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[196\] vssd1 vssd1 vccd1 vccd1 HI[196] insts\[196\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[363\] vssd1 vssd1 vccd1 vccd1 HI[363] insts\[363\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[76\] vssd1 vssd1 vccd1 vccd1 HI[76] insts\[76\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[209\] vssd1 vssd1 vccd1 vccd1 HI[209] insts\[209\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[111\] vssd1 vssd1 vccd1 vccd1 HI[111] insts\[111\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[326\] vssd1 vssd1 vccd1 vccd1 HI[326] insts\[326\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[159\] vssd1 vssd1 vccd1 vccd1 HI[159] insts\[159\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[39\] vssd1 vssd1 vccd1 vccd1 HI[39] insts\[39\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_722 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
Xinsts\[443\] vssd1 vssd1 vccd1 vccd1 HI[443] insts\[443\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_221 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_254 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xinsts\[276\] vssd1 vssd1 vccd1 vccd1 HI[276] insts\[276\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[393\] vssd1 vssd1 vccd1 vccd1 HI[393] insts\[393\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[406\] vssd1 vssd1 vccd1 vccd1 HI[406] insts\[406\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[141\] vssd1 vssd1 vccd1 vccd1 HI[141] insts\[141\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[239\] vssd1 vssd1 vccd1 vccd1 HI[239] insts\[239\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[21\] vssd1 vssd1 vccd1 vccd1 HI[21] insts\[21\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[356\] vssd1 vssd1 vccd1 vccd1 HI[356] insts\[356\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[189\] vssd1 vssd1 vccd1 vccd1 HI[189] insts\[189\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[69\] vssd1 vssd1 vccd1 vccd1 HI[69] insts\[69\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[104\] vssd1 vssd1 vccd1 vccd1 HI[104] insts\[104\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_617 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[221\] vssd1 vssd1 vccd1 vccd1 HI[221] insts\[221\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[319\] vssd1 vssd1 vccd1 vccd1 HI[319] insts\[319\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[436\] vssd1 vssd1 vccd1 vccd1 HI[436] insts\[436\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[171\] vssd1 vssd1 vccd1 vccd1 HI[171] insts\[171\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[269\] vssd1 vssd1 vccd1 vccd1 HI[269] insts\[269\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[51\] vssd1 vssd1 vccd1 vccd1 HI[51] insts\[51\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[386\] vssd1 vssd1 vccd1 vccd1 HI[386] insts\[386\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[99\] vssd1 vssd1 vccd1 vccd1 HI[99] insts\[99\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[134\] vssd1 vssd1 vccd1 vccd1 HI[134] insts\[134\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[301\] vssd1 vssd1 vccd1 vccd1 HI[301] insts\[301\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[14\] vssd1 vssd1 vccd1 vccd1 HI[14] insts\[14\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[349\] vssd1 vssd1 vccd1 vccd1 HI[349] insts\[349\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[251\] vssd1 vssd1 vccd1 vccd1 HI[251] insts\[251\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[299\] vssd1 vssd1 vccd1 vccd1 HI[299] insts\[299\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_629 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_673 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[81\] vssd1 vssd1 vccd1 vccd1 HI[81] insts\[81\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[214\] vssd1 vssd1 vccd1 vccd1 HI[214] insts\[214\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[429\] vssd1 vssd1 vccd1 vccd1 HI[429] insts\[429\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[164\] vssd1 vssd1 vccd1 vccd1 HI[164] insts\[164\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[331\] vssd1 vssd1 vccd1 vccd1 HI[331] insts\[331\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[44\] vssd1 vssd1 vccd1 vccd1 HI[44] insts\[44\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[379\] vssd1 vssd1 vccd1 vccd1 HI[379] insts\[379\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[2\] vssd1 vssd1 vccd1 vccd1 HI[2] insts\[2\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[281\] vssd1 vssd1 vccd1 vccd1 HI[281] insts\[281\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[127\] vssd1 vssd1 vccd1 vccd1 HI[127] insts\[127\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[411\] vssd1 vssd1 vccd1 vccd1 HI[411] insts\[411\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[244\] vssd1 vssd1 vccd1 vccd1 HI[244] insts\[244\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[459\] vssd1 vssd1 vccd1 vccd1 HI[459] insts\[459\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[361\] vssd1 vssd1 vccd1 vccd1 HI[361] insts\[361\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[194\] vssd1 vssd1 vccd1 vccd1 HI[194] insts\[194\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_641 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[74\] vssd1 vssd1 vccd1 vccd1 HI[74] insts\[74\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_405 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_449 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[207\] vssd1 vssd1 vccd1 vccd1 HI[207] insts\[207\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[157\] vssd1 vssd1 vccd1 vccd1 HI[157] insts\[157\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[324\] vssd1 vssd1 vccd1 vccd1 HI[324] insts\[324\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[37\] vssd1 vssd1 vccd1 vccd1 HI[37] insts\[37\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[441\] vssd1 vssd1 vccd1 vccd1 HI[441] insts\[441\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_533 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[274\] vssd1 vssd1 vccd1 vccd1 HI[274] insts\[274\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[391\] vssd1 vssd1 vccd1 vccd1 HI[391] insts\[391\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[404\] vssd1 vssd1 vccd1 vccd1 HI[404] insts\[404\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[237\] vssd1 vssd1 vccd1 vccd1 HI[237] insts\[237\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_609 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[354\] vssd1 vssd1 vccd1 vccd1 HI[354] insts\[354\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[187\] vssd1 vssd1 vccd1 vccd1 HI[187] insts\[187\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[67\] vssd1 vssd1 vccd1 vccd1 HI[67] insts\[67\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_697 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
Xinsts\[102\] vssd1 vssd1 vccd1 vccd1 HI[102] insts\[102\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_417 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[317\] vssd1 vssd1 vccd1 vccd1 HI[317] insts\[317\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[434\] vssd1 vssd1 vccd1 vccd1 HI[434] insts\[434\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_545 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[267\] vssd1 vssd1 vccd1 vccd1 HI[267] insts\[267\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_589 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[384\] vssd1 vssd1 vccd1 vccd1 HI[384] insts\[384\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_386 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[97\] vssd1 vssd1 vccd1 vccd1 HI[97] insts\[97\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[132\] vssd1 vssd1 vccd1 vccd1 HI[132] insts\[132\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[12\] vssd1 vssd1 vccd1 vccd1 HI[12] insts\[12\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[347\] vssd1 vssd1 vccd1 vccd1 HI[347] insts\[347\]/LO sky130_fd_sc_hd__conb_1
XFILLER_1_429 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[297\] vssd1 vssd1 vccd1 vccd1 HI[297] insts\[297\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[212\] vssd1 vssd1 vccd1 vccd1 HI[212] insts\[212\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[162\] vssd1 vssd1 vccd1 vccd1 HI[162] insts\[162\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[427\] vssd1 vssd1 vccd1 vccd1 HI[427] insts\[427\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_557 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_502 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[42\] vssd1 vssd1 vccd1 vccd1 HI[42] insts\[42\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[377\] vssd1 vssd1 vccd1 vccd1 HI[377] insts\[377\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_398 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_365 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[0\] vssd1 vssd1 vccd1 vccd1 HI[0] insts\[0\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[125\] vssd1 vssd1 vccd1 vccd1 HI[125] insts\[125\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[242\] vssd1 vssd1 vccd1 vccd1 HI[242] insts\[242\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[457\] vssd1 vssd1 vccd1 vccd1 HI[457] insts\[457\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[192\] vssd1 vssd1 vccd1 vccd1 HI[192] insts\[192\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[72\] vssd1 vssd1 vccd1 vccd1 HI[72] insts\[72\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[205\] vssd1 vssd1 vccd1 vccd1 HI[205] insts\[205\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_569 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_514 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[155\] vssd1 vssd1 vccd1 vccd1 HI[155] insts\[155\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[322\] vssd1 vssd1 vccd1 vccd1 HI[322] insts\[322\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[35\] vssd1 vssd1 vccd1 vccd1 HI[35] insts\[35\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[272\] vssd1 vssd1 vccd1 vccd1 HI[272] insts\[272\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_377 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_333 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[118\] vssd1 vssd1 vccd1 vccd1 HI[118] insts\[118\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_130 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_141 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[402\] vssd1 vssd1 vccd1 vccd1 HI[402] insts\[402\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[235\] vssd1 vssd1 vccd1 vccd1 HI[235] insts\[235\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_601 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_645 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[352\] vssd1 vssd1 vccd1 vccd1 HI[352] insts\[352\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[185\] vssd1 vssd1 vccd1 vccd1 HI[185] insts\[185\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[65\] vssd1 vssd1 vccd1 vccd1 HI[65] insts\[65\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[100\] vssd1 vssd1 vccd1 vccd1 HI[100] insts\[100\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[148\] vssd1 vssd1 vccd1 vccd1 HI[148] insts\[148\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_526 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
Xinsts\[315\] vssd1 vssd1 vccd1 vccd1 HI[315] insts\[315\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[28\] vssd1 vssd1 vccd1 vccd1 HI[28] insts\[28\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[265\] vssd1 vssd1 vccd1 vccd1 HI[265] insts\[265\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[432\] vssd1 vssd1 vccd1 vccd1 HI[432] insts\[432\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_345 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[382\] vssd1 vssd1 vccd1 vccd1 HI[382] insts\[382\]/LO sky130_fd_sc_hd__conb_1
XFILLER_2_197 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[95\] vssd1 vssd1 vccd1 vccd1 HI[95] insts\[95\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[130\] vssd1 vssd1 vccd1 vccd1 HI[130] insts\[130\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[228\] vssd1 vssd1 vccd1 vccd1 HI[228] insts\[228\]/LO sky130_fd_sc_hd__conb_1
XFILLER_0_613 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_657 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_12
Xinsts\[10\] vssd1 vssd1 vccd1 vccd1 HI[10] insts\[10\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[178\] vssd1 vssd1 vccd1 vccd1 HI[178] insts\[178\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[345\] vssd1 vssd1 vccd1 vccd1 HI[345] insts\[345\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[58\] vssd1 vssd1 vccd1 vccd1 HI[58] insts\[58\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[462\] vssd1 vssd1 vccd1 vccd1 HI[462] insts\[462\]/LO sky130_fd_sc_hd__conb_1
Xinsts\[295\] vssd1 vssd1 vccd1 vccd1 HI[295] insts\[295\]/LO sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_sc_hvl__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A VGND VPWR X VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt mgmt_protect_hv vccd vdda1 vdda2 mprj2_vdd_logic1 mprj_vdd_logic1 vssa1 vssd
+ vssa2
Xmprj2_logic_high_hvl vssa2 vssa2 vdda2 vdda2 mprj2_logic_high_lv/A mprj2_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_hvl vssa1 vssa1 vdda1 vdda1 mprj_logic_high_lv/A mprj_logic_high_hvl/LO
+ sky130_fd_sc_hvl__conb_1
Xmprj_logic_high_lv mprj_logic_high_lv/A vssd vdda1 mprj_vdd_logic1 vssd vdda1 vccd
+ sky130_fd_sc_hvl__lsbufhv2lv_1
Xmprj2_logic_high_lv mprj2_logic_high_lv/A vssd vdda2 mprj2_vdd_logic1 vssd vdda2
+ vccd sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd1 vccd2 vdda1 vdda2 vssa2 vssa1 vssd2 vssd vssd1
+ vccd
XFILLER_3_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1828_A wire1828/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3984 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4434 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3912 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3726 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1902 wire1903/X vssd vccd _615_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1913 wire1914/X vssd vccd wire1913/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1666 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1924 wire1924/A vssd vccd wire1924/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1935 wire1936/X vssd vccd wire1935/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1946 wire1947/X vssd vccd wire1946/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1957 wire1958/X vssd vccd _595_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1968 wire1968/A vssd vccd wire1968/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1979 wire1980/X vssd vccd _584_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input127_A la_data_out_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2044_A wire2044/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_501_ _501_/A _501_/B vssd vccd _501_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_202 _262_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_213 _230_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_224 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_235 _186_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_246 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_257 _480_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_432_ _560_/A _432_/B _432_/C vssd vccd _432_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_26_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_268 _544_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_279 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_363_ _363_/A _363_/B vssd vccd _363_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_35_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input92_A la_data_out_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_294_ _294_/A _294_/B vssd vccd _294_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_48_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[8\] mprj_dat_i_user[8] max_length1311/X vssd vccd _122_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4051 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1419 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4095 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2710 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output513_A wire1143/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1144_A _370_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1409_A wire1410/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] _188_/X vssd vccd _008_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1680_A wire1681/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1778_A wire1779/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1362 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__304__A _304_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1945_A wire1946/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput467 wire1063/X vssd vccd la_data_in_core[103] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput478 _482_/X vssd vccd la_data_in_core[113] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput489 _492_/X vssd vccd la_data_in_core[123] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2687 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1209 wire1210/X vssd vccd wire1209/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_792 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__A_N _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1126 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__214__A _214_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4382 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2161_A wire2161/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input244_A la_iena_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2186 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1710 wire1710/A vssd vccd _358_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1721 wire1722/X vssd vccd wire1721/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1732 wire1733/X vssd vccd _291_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1743 wire1743/A vssd vccd wire1743/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1754 wire1754/A vssd vccd wire1754/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input411_A mprj_adr_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1765 wire1766/X vssd vccd _276_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1776 wire1776/A vssd vccd wire1776/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1787 wire1788/X vssd vccd _264_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1798 wire1798/A vssd vccd _258_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_415_ _415_/A_N _415_/B _415_/C vssd vccd _415_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_32_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_346_ _346_/A _346_/B vssd vccd _346_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_30_957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1204 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_277_ _277_/A _277_/B vssd vccd _277_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_3972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output463_A wire1145/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4135 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_880 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1261_A _320_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1359_A wire1359/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1526_A wire1526/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1895_A wire1896/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__034__A _034_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1170 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1006 _550_/X vssd vccd wire1006/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1017 _539_/X vssd vccd wire1017/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1028 _521_/X vssd vccd wire1028/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1039 _510_/X vssd vccd wire1039/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1903 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__209__A _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_570 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_200_ _200_/A _200_/B vssd vccd _200_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_51_2837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2007_A wire2008/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_131_ _131_/A vssd vccd _131_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_36_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input194_A la_iena_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1092 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4411 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_062_ _062_/A vssd vccd _062_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_7_4505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__386__A_N _514_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4455 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input361_A la_oenb_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input459_A mprj_we_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input55_A la_data_out_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4010 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__598__B _598_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_512 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1540 wire1540/A vssd vccd _574_/A vssd vccd sky130_fd_sc_hd__buf_8
Xwire1551 wire1551/A vssd vccd _563_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1573 input31/X vssd vccd _493_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1584 wire1584/A vssd vccd _619_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1595 wire1595/A vssd vccd _608_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__119__A _119_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3146 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output580_A wire1076/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1107_A _406_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_329_ _329_/A _329_/B vssd vccd _329_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output845_A _596_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1476_A wire1476/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] wire1322/X vssd vccd wire965/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_45_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1643_A wire1644/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__301__B _301_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1908_A wire1909/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_710 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1210 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2338 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__211__B _211_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_810 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_526 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2124_A wire2125/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input207_A la_iena_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_114_ _114_/A vssd vccd _114_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_2331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_045_ _045_/A vssd vccd _045_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_49_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3391 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2060 wire2061/X vssd vccd _499_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2071 wire2072/X vssd vccd wire2071/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2082 wire2083/X vssd vccd _491_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2093 wire2093/A vssd vccd wire2093/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1057_A _478_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__401__A_N _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1370 wire1370/A vssd vccd _358_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_39_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1381 wire1382/X vssd vccd _351_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1392 wire1393/X vssd vccd wire1392/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1224_A wire1225/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output795_A wire1005/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[20\] mprj_dat_i_user[20] _294_/X vssd vccd _134_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_30_2729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1760_A wire1760/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1858_A wire1858/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__312__A _312_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__B _206_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3976 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3746 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2074_A wire2075/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input157_A la_iena_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput301 la_oenb_mprj[21] vssd vccd _518_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__424__A_N _552_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput312 la_oenb_mprj[31] vssd vccd _400_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput323 la_oenb_mprj[41] vssd vccd _538_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput334 la_oenb_mprj[51] vssd vccd _420_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput345 la_oenb_mprj[61] vssd vccd _558_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput356 la_oenb_mprj[71] vssd vccd wire1546/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput367 la_oenb_mprj[81] vssd vccd wire1536/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input324_A la_oenb_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1000 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput378 la_oenb_mprj[91] vssd vccd _588_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput389 mprj_adr_o_core[10] vssd vccd wire1521/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input18_A la_data_out_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_594_ _594_/A _594_/B vssd vccd _594_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_16_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2540 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1774 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_5 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput808 _562_/X vssd vccd la_oenb_core[65] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput819 _572_/X vssd vccd la_oenb_core[75] vssd vccd sky130_fd_sc_hd__buf_8
X_028_ _028_/A vssd vccd _028_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output543_A wire1084/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__132__A _132_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1174_A wire1175/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3234 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3328 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output808_A _562_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1439_A wire1440/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2599 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] _218_/X vssd vccd _038_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_48_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_610 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4362 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__307__A _307_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1975_A wire1975/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__447__A_N _575_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1815 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4491 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_142 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__217__A _217_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input274_A la_oenb_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2191_A wire2191/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input441_A mprj_dat_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput120 la_data_out_mprj[8] vssd vccd _377_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput131 la_data_out_mprj[9] vssd vccd _378_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput142 la_iena_mprj[109] vssd vccd _272_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput153 la_iena_mprj[119] vssd vccd _282_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput164 la_iena_mprj[13] vssd vccd _176_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput175 la_iena_mprj[23] vssd vccd wire1615/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput186 la_iena_mprj[33] vssd vccd _196_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput197 la_iena_mprj[43] vssd vccd _206_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3314 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_577_ _577_/A _577_/B vssd vccd _577_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2635 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output493_A _496_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__127__A _127_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output660_A _030_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output758_A wire1052/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1291_A wire1292/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4019 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput605 _095_/Y vssd vccd la_data_in_mprj[112] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1389_A wire1390/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput616 _105_/Y vssd vccd la_data_in_mprj[122] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput627 _000_/Y vssd vccd la_data_in_mprj[17] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput638 _010_/Y vssd vccd la_data_in_mprj[27] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output925_A wire1190/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput649 _020_/Y vssd vccd la_data_in_mprj[37] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3294 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1723_A wire1724/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4495 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4446 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__037__A _037_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_B _197_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1087 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1903 wire1904/X vssd vccd wire1903/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__500__A _500_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1914 wire1914/A vssd vccd wire1914/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1678 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1925 wire1926/X vssd vccd _608_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1936 wire1936/A vssd vccd wire1936/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_2081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1947 wire1947/A vssd vccd wire1947/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1958 wire1958/A vssd vccd wire1958/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1969 wire1970/X vssd vccd _591_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_500_ _500_/A _500_/B vssd vccd _500_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_19_3612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_203 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_214 _230_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_225 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2037_A wire2038/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_236 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_431_ _559_/A _431_/B _431_/C vssd vccd _431_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_14_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_247 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_258 _480_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_269 _197_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_362_ _362_/A _362_/B vssd vccd _362_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_9_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_293_ _293_/A _293_/B vssd vccd _293_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input391_A mprj_adr_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input85_A la_data_out_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2587 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_856 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4328 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output506_A wire1121/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1137_A _377_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1304_A wire1305/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output875_A _310_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] _181_/X vssd vccd _001_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_31_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1673_A wire1673/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[16\]_B _179_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[100\]_B _263_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__304__B _304_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2600 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1840_A wire1840/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput468 wire1062/X vssd vccd la_data_in_core[104] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1938_A wire1938/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput479 _483_/X vssd vccd la_data_in_core[114] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_1910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__320__A _320_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__214__B _214_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_826 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4394 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4236 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__230__A _230_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1700 wire1701/X vssd vccd _364_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1711 wire1711/A vssd vccd _357_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1722 wire1722/A vssd vccd wire1722/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2154_A wire2154/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input237_A la_iena_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1733 wire1734/X vssd vccd wire1733/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1744 wire1745/X vssd vccd _286_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1755 wire1756/X vssd vccd _281_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1766 wire1766/A vssd vccd wire1766/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1777 wire1777/A vssd vccd _270_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1788 wire1788/A vssd vccd wire1788/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1799 wire1799/A vssd vccd _257_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input404_A mprj_adr_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_414_ _542_/A _414_/B _414_/C vssd vccd _414_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_966 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_345_ _345_/A _345_/B vssd vccd _345_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2952 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_276_ _276_/A _276_/B vssd vccd _276_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_2351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1216 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4103 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4147 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1087_A wire1088/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__140__A _140_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1254_A wire1255/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2530 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2596 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1421_A wire1421/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1519_A wire1519/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1888_A wire1888/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__315__A _315_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1182 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3991 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__050__A _050_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1007 wire1008/X vssd vccd wire1007/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1604 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1018 _538_/X vssd vccd wire1018/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1029 _520_/X vssd vccd wire1029/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1915 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__209__B _209_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_582 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4084 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_130_ _130_/A vssd vccd _130_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_7_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__225__A _225_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_2682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_061_ _061_/A vssd vccd _061_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_27_4423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input187_A la_iena_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4467 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input354_A la_oenb_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3608 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4191 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input48_A la_data_out_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1530 wire1530/A vssd vccd _584_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1541 wire1541/A vssd vccd _573_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1552 wire1552/A vssd vccd _562_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1563 _415_/A_N vssd vccd _543_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1574 wire1574/A vssd vccd _526_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1585 wire1585/A vssd vccd _618_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1596 _479_/A_N vssd vccd _607_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_46_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1002_A wire1003/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_328_ _328_/A _328_/B vssd vccd _328_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_15_2479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output573_A _453_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__135__A _135_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_259_ _259_/A _259_/B vssd vccd _259_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output740_A _616_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output838_A _589_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1371_A wire1371/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1469_A wire1470/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1014 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__A_N _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] wire1329/X vssd vccd wire972/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_44_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3815 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1222 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__045__A _045_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4320 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4458 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_822 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_538 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input102_A la_data_out_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2117_A wire2118/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_113_ _113_/A vssd vccd _113_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_044_ _044_/A vssd vccd _044_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3416 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3140 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2050 wire2050/A vssd vccd wire2050/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2061 wire2061/A vssd vccd wire2061/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2072 wire2072/A vssd vccd wire2072/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2083 wire2084/X vssd vccd wire2083/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2094 wire2095/X vssd vccd _487_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1360 wire1361/X vssd vccd _339_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1371 wire1371/A vssd vccd _357_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1382 wire1382/A vssd vccd wire1382/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1393 wire1393/A vssd vccd wire1393/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1217_A wire1218/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output690_A _057_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output788_A _544_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output955_A wire1307/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[13\] mprj_dat_i_user[13] max_length1311/X vssd vccd _127_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_28_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1753_A wire1754/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__312__B _312_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_A mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1920_A wire1921/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] _274_/X vssd vccd wire988/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_1_3790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__A_N _504_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2696 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4415 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3703 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput302 la_oenb_mprj[22] vssd vccd _519_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput313 la_oenb_mprj[32] vssd vccd wire1570/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput324 la_oenb_mprj[42] vssd vccd _539_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput335 la_oenb_mprj[52] vssd vccd _549_/A vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_wire2067_A wire2068/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput346 la_oenb_mprj[62] vssd vccd wire1555/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput357 la_oenb_mprj[72] vssd vccd wire1545/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput368 la_oenb_mprj[82] vssd vccd wire1535/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput379 la_oenb_mprj[92] vssd vccd _589_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input317_A la_oenb_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_593_ _593_/A _593_/B vssd vccd _593_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2596 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_6 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput809 _563_/X vssd vccd la_oenb_core[66] vssd vccd sky130_fd_sc_hd__buf_8
X_027_ _027_/A vssd vccd _027_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_2924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output536_A wire1093/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1167_A wire1168/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_990 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__399__A_N _527_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1190 wire1191/X vssd vccd wire1190/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_39_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] _211_/X vssd vccd _031_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1501_A wire1502/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4374 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__307__B _307_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1870_A wire1870/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1968_A wire1968/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__A _323_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3791 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4230 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_154 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_894 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__A _233_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2184_A wire2185/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input267_A la_oenb_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_710 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input434_A mprj_dat_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput110 la_data_out_mprj[80] vssd vccd wire1624/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput121 la_data_out_mprj[90] vssd vccd _459_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input30_A la_data_out_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput132 la_iena_mprj[0] vssd vccd _625_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput143 la_iena_mprj[10] vssd vccd _173_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput154 la_iena_mprj[11] vssd vccd _174_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput165 la_iena_mprj[14] vssd vccd _177_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput176 la_iena_mprj[24] vssd vccd wire1614/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput187 la_iena_mprj[34] vssd vccd _197_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_2650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput198 la_iena_mprj[44] vssd vccd _207_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_576_ _576_/A _576_/B vssd vccd _576_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_16_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1236 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output486_A _489_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output653_A _023_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput606 _096_/Y vssd vccd la_data_in_mprj[113] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__143__A _143_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput617 _106_/Y vssd vccd la_data_in_mprj[123] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1284_A wire1285/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput628 _001_/Y vssd vccd la_data_in_mprj[18] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput639 _011_/Y vssd vccd la_data_in_mprj[28] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2776 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output820_A _573_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output918_A wire1211/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1451_A wire1451/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1716_A wire1716/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3860 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2026 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3003 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__A_N _542_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__053__A _053_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1099 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1904 wire1904/A vssd vccd wire1904/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__500__B _500_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1915 wire1916/X vssd vccd _611_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1926 wire1927/X vssd vccd wire1926/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1937 wire1938/X vssd vccd _604_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1948 wire1949/X vssd vccd _599_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1959 wire1960/X vssd vccd _297_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_204 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_215 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_226 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_237 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_430_ _558_/A _430_/B _430_/C vssd vccd _430_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_248 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_259 _480_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__228__A _228_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_361_ _361_/A _361_/B vssd vccd _361_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_14_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_292_ _292_/A _292_/B vssd vccd _292_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_42_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input384_A la_oenb_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2599 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input78_A la_data_out_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__B _410_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1032_A _517_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__437__A_N _565_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__138__A _138_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_2433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_559_ _559_/A _559_/B vssd vccd _559_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_14_2308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output868_A _333_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1499_A wire1500/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1666_A wire1667/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput469 wire1061/X vssd vccd la_data_in_core[105] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__601__A _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2415 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1833_A wire1834/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__320__B _320_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__048__A _048_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1231 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4362 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__511__A _511_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__230__B _230_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1701 wire1701/A vssd vccd wire1701/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1712 wire1712/A vssd vccd _356_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1723 wire1724/X vssd vccd wire1723/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1734 wire1734/A vssd vccd wire1734/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1745 wire1745/A vssd vccd wire1745/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input132_A la_iena_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1756 wire1756/A vssd vccd wire1756/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1767 wire1768/X vssd vccd _275_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2147_A wire2148/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1778 wire1779/X vssd vccd _269_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1789 wire1790/X vssd vccd _263_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_413_ _541_/A _413_/B _413_/C vssd vccd _413_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_37_1629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_344_ _344_/A _344_/B vssd vccd _344_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_53_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_275_ _275_/A _275_/B vssd vccd _275_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2964 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__405__B _405_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4159 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1207 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output616_A _105_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1247_A wire1248/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1414_A wire1415/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] _193_/X vssd vccd _013_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_33_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__315__B _315_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1950_A wire1951/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__331__A _331_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1008 _549_/X vssd vccd wire1008/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1019 _536_/X vssd vccd wire1019/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1616 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_4397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_A mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4096 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_594 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3362 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__A _506_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__225__B _225_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_060_ _060_/A vssd vccd _060_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_20_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2097_A wire2098/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__241__A _241_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input347_A la_oenb_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1520 wire1521/X vssd vccd _315_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1531 wire1531/A vssd vccd _583_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1542 wire1542/A vssd vccd _572_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_21_2643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1553 wire1553/A vssd vccd _561_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1564 _412_/A_N vssd vccd _540_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_24_1076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1575 wire1575/A vssd vccd _524_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1586 wire1586/A vssd vccd _617_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1597 _478_/A_N vssd vccd _606_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2583 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_327_ _327_/A _327_/B vssd vccd _327_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_258_ _258_/A _258_/B vssd vccd _258_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_3760 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output566_A _447_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_189_ _189_/A _189_/B vssd vccd _189_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_45_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output733_A _609_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1364_A wire1364/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1026 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2576 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] _241_/X vssd vccd wire978/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_6_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1531_A wire1531/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1629_A wire1629/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3950 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4372 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1998_A wire1999/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_594 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__A _326_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1234 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__061__A _061_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4103 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1779 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2012_A wire2013/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__236__A _236_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input297_A la_oenb_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_112_ _112_/A vssd vccd _112_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_043_ _043_/A vssd vccd _043_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2355 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input60_A la_data_out_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__402__C _402_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3428 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2040 wire2041/X vssd vccd _511_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2051 wire2051/A vssd vccd _505_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2062 wire2063/X vssd vccd _498_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2073 wire2074/X vssd vccd _494_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_300 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2670 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2084 wire2084/A vssd vccd wire2084/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1350 wire1351/X vssd vccd _343_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2095 wire2096/X vssd vccd wire2095/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1361 wire1361/A vssd vccd wire1361/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1372 wire1373/X vssd vccd _338_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1383 wire1384/X vssd vccd _350_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1394 wire1395/X vssd vccd _298_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_870 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_594 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output683_A _051_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output850_A wire1268/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output948_A wire1280/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1746_A wire1747/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[1\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1913_A wire1914/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] _267_/X vssd vccd _087_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_17_3700 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3608 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__056__A _056_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__503__B _503_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3715 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4140 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3759 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput303 la_oenb_mprj[23] vssd vccd _520_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput314 la_oenb_mprj[33] vssd vccd _530_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4184 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput325 la_oenb_mprj[43] vssd vccd _412_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput336 la_oenb_mprj[53] vssd vccd _550_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput347 la_oenb_mprj[63] vssd vccd wire1554/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput358 la_oenb_mprj[73] vssd vccd wire1544/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput369 la_oenb_mprj[83] vssd vccd wire1534/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input212_A la_iena_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_592_ _592_/A _592_/B vssd vccd _592_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__A_N _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_7 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4051 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_026_ _026_/A vssd vccd _026_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__413__B _413_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4095 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output529_A wire1100/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1062_A _473_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1180 wire1181/X vssd vccd wire1180/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1191 wire1192/X vssd vccd wire1191/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1327_A _250_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1696_A wire1697/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1362 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__A _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1395 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1863_A wire1864/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__323__B _323_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1806 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__493__A_N _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_4242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__514__A _514_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_2472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_4432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__233__B _233_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input162_A la_iena_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2177_A wire2178/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput100 la_data_out_mprj[71] vssd vccd wire1633/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput111 la_data_out_mprj[81] vssd vccd wire1623/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput122 la_data_out_mprj[91] vssd vccd _460_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput133 la_iena_mprj[100] vssd vccd _263_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput144 la_iena_mprj[110] vssd vccd _273_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input427_A mprj_dat_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput155 la_iena_mprj[120] vssd vccd _283_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput166 la_iena_mprj[15] vssd vccd _178_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input23_A la_data_out_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput177 la_iena_mprj[25] vssd vccd wire1613/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput188 la_iena_mprj[35] vssd vccd _198_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput199 la_iena_mprj[45] vssd vccd _208_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_29_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_575_ _575_/A _575_/B vssd vccd _575_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__408__B _408_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_2659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output479_A _483_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
Xoutput607 _097_/Y vssd vccd la_data_in_mprj[114] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3528 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput618 _107_/Y vssd vccd la_data_in_mprj[124] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput629 _002_/Y vssd vccd la_data_in_mprj[19] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output646_A _017_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_009_ _009_/A vssd vccd _009_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_46_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1277_A _312_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output813_A wire1047/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1444_A wire1445/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] _223_/X vssd vccd _043_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_2387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1709_A wire1709/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3872 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__318__B _318_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3015 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1980_A wire1980/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4194 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__334__A _334_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_max_length1311_A _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1905 wire1906/X vssd vccd _614_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1916 wire1917/X vssd vccd wire1916/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1927 wire1927/A vssd vccd wire1927/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1938 wire1938/A vssd vccd wire1938/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1949 wire1949/A vssd vccd wire1949/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_205 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_216 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_227 _204_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__509__A _509_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_238 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_249 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__228__B _228_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_360_ _360_/A _360_/B vssd vccd _360_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_17_3360 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_291_ _291_/A _291_/B vssd vccd _291_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_52_3295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__A _244_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__389__A_N _517_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input377_A la_oenb_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__410__C _410_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_558_ _558_/A _558_/B vssd vccd _558_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_wire1025_A _525_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output596_A _087_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_489_ _617_/A _489_/B _489_/C vssd vccd _489_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_20_618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output763_A wire1028/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1394_A wire1395/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output930_A wire1170/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_4059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3106 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1561_A wire1561/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3128 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1659_A wire1660/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__601__B _601_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2427 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1826_A wire1826/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__329__A _329_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1243 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1899 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__064__A _064_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3927 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput960 _295_/X vssd vccd user_reset vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__511__B _511_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2950 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1702 wire1703/X vssd vccd _363_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1713 wire1713/A vssd vccd _355_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1724 wire1725/X vssd vccd wire1724/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1735 wire1736/X vssd vccd _290_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1746 wire1747/X vssd vccd _285_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1757 wire1758/X vssd vccd _280_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1768 wire1768/A vssd vccd wire1768/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1779 wire1779/A vssd vccd wire1779/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2042_A wire2043/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input125_A la_data_out_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__239__A _239_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_412_ _412_/A_N _412_/B _412_/C vssd vccd _412_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_3319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3488 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_343_ _343_/A _343_/B vssd vccd _343_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_52_3070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input90_A la_data_out_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_274_ _274_/A _274_/B vssd vccd _274_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__C _405_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[6\] mprj_dat_i_user[6] max_length1311/X vssd vccd _120_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_10_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__421__B _421_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__A_N _532_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output511_A wire1116/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output609_A _099_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1142_A _372_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1407_A wire1408/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3820 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output880_A wire1306/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] _186_/X vssd vccd _006_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1776_A wire1776/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__612__A _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1943_A wire1944/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__331__B _331_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3802 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1009 wire1010/X vssd vccd wire1009/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__059__A _059_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_ack_gate_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__506__B _506_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_2640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__522__A _522_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__A_N _555_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__241__B _241_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2200 wire2200/A vssd vccd _306_/A vssd vccd sky130_fd_sc_hd__buf_6
Xoutput790 wire1011/X vssd vccd la_oenb_core[49] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_4118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input242_A la_iena_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3334 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1510 wire1511/X vssd vccd wire1510/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1521 wire1521/A vssd vccd wire1521/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1532 wire1532/A vssd vccd _582_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1543 wire1543/A vssd vccd _571_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1554 wire1554/A vssd vccd _560_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1565 _409_/A_N vssd vccd _537_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1576 wire1577/X vssd vccd _295_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1587 wire1587/A vssd vccd _616_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1598 input27/X vssd vccd _489_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_21_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_570 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2595 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_326_ _326_/A _326_/B vssd vccd _326_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_9_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__B _416_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_257_ _257_/A _257_/B vssd vccd _257_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_7_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_188_ _188_/A _188_/B vssd vccd _188_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_output559_A _440_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1092_A _420_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output726_A _603_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1038 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1357_A wire1357/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1524_A wire1525/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__A _607_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4384 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1893_A wire1894/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__326__B _326_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire977_A wire977/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[91\]_B wire1323/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__A _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2760 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__517__A _517_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__236__B _236_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2005_A wire2006/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_3182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_111_ _111_/A vssd vccd _111_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_14_2470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input192_A la_iena_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_042_ _042_/A vssd vccd _042_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_50_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__252__A _252_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input457_A mprj_sel_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4299 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input53_A la_data_out_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire2030 wire2030/A vssd vccd _520_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2041 wire2041/A vssd vccd wire2041/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2052 wire2052/A vssd vccd _504_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2063 wire2063/A vssd vccd wire2063/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2074 wire2075/X vssd vccd wire2074/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3175 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2502 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1340 input85/X vssd vccd _427_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire2085 wire2086/X vssd vccd _490_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1351 wire1351/A vssd vccd wire1351/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2096 wire2096/A vssd vccd wire2096/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1362 wire1362/A vssd vccd _366_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1373 wire1374/X vssd vccd wire1373/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1384 wire1384/A vssd vccd wire1384/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1395 wire1396/X vssd vccd wire1395/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2802 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_882 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1105_A _408_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_309_ _309_/A _309_/B vssd vccd _309_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_user_to_mprj_in_gates\[73\]_B _236_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3580 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output843_A _594_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3318 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__162__A _162_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1474_A wire1474/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] wire1324/X vssd vccd wire967/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_28_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1641_A wire1642/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1739_A wire1739/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1906_A wire1907/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3712 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__A _337_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_576 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3388 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__072__A _072_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput304 la_oenb_mprj[24] vssd vccd _521_/A vssd vccd sky130_fd_sc_hd__clkbuf_8
XFILLER_0_458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput315 la_oenb_mprj[34] vssd vccd _531_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_44_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput326 la_oenb_mprj[44] vssd vccd _541_/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput337 la_oenb_mprj[54] vssd vccd _551_/A vssd vccd sky130_fd_sc_hd__buf_8
Xinput348 la_oenb_mprj[64] vssd vccd wire1553/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput359 la_oenb_mprj[74] vssd vccd wire1543/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_591_ _591_/A _591_/B vssd vccd _591_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_21_1069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2122_A wire2122/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input205_A la_iena_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__247__A _247_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_025_ _025_/A vssd vccd _025_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_8 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__413__C _413_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4063 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1170 wire1171/X vssd vccd wire1170/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_19_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1181 _360_/X vssd vccd wire1181/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1192 wire1193/X vssd vccd wire1192/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__295__A_N _295_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1222_A _348_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output793_A _548_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1920 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1076 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1689_A wire1689/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1374 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__604__B _604_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1856_A wire1856/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2447 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__A _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__067__A _067_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[37\]_B _200_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_B _284_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__514__B _514_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__530__A _530_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3535 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input155_A la_iena_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput101 la_data_out_mprj[72] vssd vccd wire1632/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput112 la_data_out_mprj[82] vssd vccd wire1622/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput123 la_data_out_mprj[92] vssd vccd _461_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput134 la_iena_mprj[101] vssd vccd _264_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput145 la_iena_mprj[111] vssd vccd _274_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput156 la_iena_mprj[121] vssd vccd _284_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input322_A la_oenb_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput167 la_iena_mprj[16] vssd vccd _179_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput178 la_iena_mprj[26] vssd vccd wire1612/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput189 la_iena_mprj[36] vssd vccd _199_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input16_A la_data_out_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_574_ _574_/A _574_/B vssd vccd _574_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_user_wb_dat_gates\[30\]_A mprj_dat_i_user[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3940 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_184 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__424__B _424_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[112\]_B _275_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput608 _098_/Y vssd vccd la_data_in_mprj[115] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput619 _108_/Y vssd vccd la_data_in_mprj[125] vssd vccd sky130_fd_sc_hd__buf_8
X_008_ _008_/A vssd vccd _008_/Y vssd vccd sky130_fd_sc_hd__inv_4
XANTENNA_output541_A wire1087/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output639_A _011_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1172_A wire1173/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output806_A _560_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1437_A wire1438/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] _216_/X vssd vccd _036_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1604_A _472_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[21\]_A mprj_dat_i_user[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3027 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__A _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1973_A wire1974/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B _182_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__334__B _334_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_B wire1316/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4523 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__350__A _350_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2288 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4280 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__460__A_N _588_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input8_A la_data_out_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_1418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1906 wire1907/X vssd vccd wire1906/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1917 wire1918/X vssd vccd wire1917/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1928 wire1929/X vssd vccd _607_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1939 wire1940/X vssd vccd _603_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_206 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_217 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__509__B _509_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_228 _204_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_239 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[12\]_A mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3372 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_290_ _290_/A _290_/B vssd vccd _290_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__525__A _525_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__244__B _244_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input272_A la_oenb_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__260__A _260_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__B _419_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_557_ _557_/A _557_/B vssd vccd _557_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1018_A _538_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_488_ _616_/A _488_/B _488_/C vssd vccd _488_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output491_A _494_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output589_A wire1067/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3792 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output756_A wire1034/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4038 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3304 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1387_A wire1388/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__483__A_N _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output923_A wire1194/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__170__A _170_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2439 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4486 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1721_A wire1722/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__329__B _329_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1856 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__A _345_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3939 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__080__A _080_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput950 wire1299/X vssd vccd mprj_we_o_user vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_4375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1423 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1703 wire1703/A vssd vccd wire1703/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1714 wire1714/A vssd vccd _300_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1725 wire1725/A vssd vccd wire1725/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1736 wire1737/X vssd vccd wire1736/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4102 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1747 wire1748/X vssd vccd wire1747/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1758 wire1758/A vssd vccd wire1758/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_1000 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1769 wire1770/X vssd vccd _274_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_1011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__239__B _239_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2035_A wire2035/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input118_A la_data_out_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_411_ _539_/A _411_/B _411_/C vssd vccd _411_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_27_796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_446 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_342_ _342_/A _342_/B vssd vccd _342_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_30_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__255__A _255_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_273_ _273_/A _273_/B vssd vccd _273_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input83_A la_data_out_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__421__C _421_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2691 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output504_A wire1123/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1135_A _379_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_609_ _609_/A _609_/B vssd vccd _609_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_53_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3832 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1302_A _300_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output873_A _308_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_939 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__165__A _165_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] _179_/X vssd vccd _163_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
Xuser_wb_dat_gates\[29\] mprj_dat_i_user[29] max_length1310/X vssd vccd _143_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_31_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1671_A wire1671/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1769_A wire1770/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__612__B _612_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1936_A wire1936/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] _290_/X vssd vccd wire979/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_0_4355 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__379__A_N _507_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__075__A _075_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_950 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3703 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__522__B _522_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput780 wire1050/X vssd vccd la_oenb_core[3] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2201 wire2202/X vssd vccd _305_/A vssd vccd sky130_fd_sc_hd__buf_6
Xoutput791 wire1049/X vssd vccd la_oenb_core[4] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1500 wire1500/A vssd vccd wire1500/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3346 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1511 wire1511/A vssd vccd wire1511/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input235_A la_iena_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1522 wire1523/X vssd vccd _305_/B vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire2152_A wire2153/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1533 wire1533/A vssd vccd _581_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1544 wire1544/A vssd vccd _570_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1555 wire1555/A vssd vccd _559_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1566 input32/X vssd vccd _494_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1577 wire1578/X vssd vccd wire1577/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1588 wire1588/A vssd vccd _615_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1599 _477_/A_N vssd vccd _605_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_41_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input402_A mprj_adr_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_325_ _325_/A _325_/B vssd vccd _325_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_30_736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__416__C _416_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_256_ _256_/A _256_/B vssd vccd _256_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_7_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_187_ _187_/A _187_/B vssd vccd _187_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_48_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__B _432_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1085_A wire1086/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output719_A wire1053/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1252_A _337_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1517_A wire1517/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__607__B _607_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1886_A wire1887/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__A _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1583 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__342__B _342_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[4\]_A mprj_dat_i_user[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__517__B _517_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_110_ _110_/A vssd vccd _110_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__533__A _533_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_041_ _041_/A vssd vccd _041_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_50_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input185_A la_iena_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__252__B _252_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input352_A la_oenb_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input46_A la_data_out_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2020 wire2020/A vssd vccd _561_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2031 wire2031/A vssd vccd _519_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2042 wire2043/X vssd vccd _510_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2053 wire2054/X vssd vccd _503_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2064 wire2065/X vssd vccd _497_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1330 _247_/X vssd vccd wire1330/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire2075 wire2075/A vssd vccd wire2075/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1341 wire1341/A vssd vccd _300_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2086 wire2087/X vssd vccd wire2086/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1352 wire1353/X vssd vccd _342_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2097 wire2098/X vssd vccd _486_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1363 wire1363/A vssd vccd _365_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1374 wire1374/A vssd vccd wire1374/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2558 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1385 wire1386/X vssd vccd _349_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1396 wire1397/X vssd vccd wire1396/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__427__B _427_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2814 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_308_ _308_/A _308_/B vssd vccd _308_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1000_A wire1001/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output571_A _451_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_239_ _239_/A _239_/B vssd vccd _239_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_3592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output836_A wire994/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1467_A wire1468/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] wire1331/X vssd vccd wire974/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_26_3098 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1634_A wire1634/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__618__A _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4160 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__337__B _337_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__417__A_N _417_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_588 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__353__A _353_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1055 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput305 la_oenb_mprj[25] vssd vccd _522_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput316 la_oenb_mprj[35] vssd vccd wire1569/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput327 la_oenb_mprj[45] vssd vccd _542_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_22_3452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput338 la_oenb_mprj[55] vssd vccd _552_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput349 la_oenb_mprj[65] vssd vccd wire1552/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1026 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_590_ _590_/A _590_/B vssd vccd _590_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_2889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3292 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__A _528_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input100_A la_data_out_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2115_A wire2116/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__263__A _263_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_024_ _024_/A vssd vccd _024_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_9 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2938 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4075 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2651 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1160 wire1161/X vssd vccd wire1160/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1171 wire1172/X vssd vccd wire1171/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1182 wire1183/X vssd vccd wire1182/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_2344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1193 _357_/X vssd vccd wire1193/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1048_A _502_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1215_A wire1216/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output786_A wire1013/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output953_A wire2205/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__173__A _173_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[11\] mprj_dat_i_user[11] _294_/X vssd vccd _125_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_51_2991 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1751_A wire1752/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1849_A wire1849/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__620__B _620_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3888 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__348__A _348_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1186 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_363 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__083__A _083_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__530__B _530_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3547 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput102 la_data_out_mprj[73] vssd vccd wire1631/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput113 la_data_out_mprj[83] vssd vccd wire1621/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput124 la_data_out_mprj[93] vssd vccd _462_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire2065_A wire2065/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input148_A la_iena_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput135 la_iena_mprj[102] vssd vccd _265_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput146 la_iena_mprj[112] vssd vccd _275_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_22_3271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput157 la_iena_mprj[122] vssd vccd _285_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput168 la_iena_mprj[17] vssd vccd _180_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput179 la_iena_mprj[27] vssd vccd _190_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_29_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2592 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input315_A la_oenb_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__258__A _258_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_636 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_573_ _573_/A _573_/B vssd vccd _573_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[30\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3952 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__424__C _424_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput609 _099_/Y vssd vccd la_data_in_mprj[116] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_007_ _007_/A vssd vccd _007_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__B _440_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output534_A wire1095/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1165_A _364_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1332_A _243_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__168__A _168_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] _209_/X vssd vccd _029_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[21\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3039 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__615__B _615_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1003 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1183 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3906 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] _171_/X vssd vccd _155_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XANTENNA__350__B _350_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4292 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1907 wire1907/A vssd vccd wire1907/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1918 wire1918/A vssd vccd wire1918/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1929 wire1930/X vssd vccd wire1929/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__078__A _078_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_207 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_218 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_229 _204_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_978 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[12\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__525__B _525_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__541__A _541_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2182_A wire2183/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input265_A la_oenb_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__260__B _260_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4067 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input432_A mprj_dat_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2450 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_625_ _625_/A _625_/B vssd vccd _625_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_29_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__419__C _419_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_556_ _556_/A _556_/B vssd vccd _556_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_487_ _615_/A _487_/B _487_/C vssd vccd _487_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_32_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__435__B _435_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output484_A _488_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output651_A _022_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output749_A _624_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1282_A wire1283/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output916_A wire1217/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3742 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1714_A wire1714/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4258 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__345__B _345_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3907 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__361__A _361_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput940 wire1238/X vssd vccd mprj_dat_o_user[5] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput951 wire1723/X vssd vccd user1_vcc_powergood vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1435 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1704 wire1705/X vssd vccd _362_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1715 wire1715/A vssd vccd _354_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1726 wire1727/X vssd vccd _293_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1737 wire1737/A vssd vccd wire1737/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1748 wire1748/A vssd vccd wire1748/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1759 wire1760/X vssd vccd _279_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_410_ _538_/A _410_/B _410_/C vssd vccd _410_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_2_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_341_ _341_/A _341_/B vssd vccd _341_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_36_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_458 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__255__B _255_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_272_ _272_/A _272_/B vssd vccd _272_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input382_A la_oenb_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input76_A la_data_out_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__271__A _271_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_608_ _608_/A _608_/B vssd vccd _608_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1030_A _519_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1128_A _385_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_539_ _539_/A _539_/B vssd vccd _539_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3844 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__450__A_N _578_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output866_A _331_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1497_A wire1497/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__181__A _181_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1664_A wire1665/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1831_A wire1832/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1929_A wire1930/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__356__A _356_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_2653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__091__A _091_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1286 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3759 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput770 _527_/X vssd vccd la_oenb_core[30] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput781 _537_/X vssd vccd la_oenb_core[40] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2202 wire2202/A vssd vccd wire2202/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput792 wire1009/X vssd vccd la_oenb_core[50] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1501 wire1502/X vssd vccd _321_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1512 wire1513/X vssd vccd _318_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1523 wire1524/X vssd vccd wire1523/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1534 wire1534/A vssd vccd _580_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1545 wire1545/A vssd vccd _569_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input130_A la_data_out_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1556 wire1556/A vssd vccd _555_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2145_A wire2145/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1567 _406_/A_N vssd vccd _534_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1578 input3/X vssd vccd wire1578/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input228_A la_iena_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1589 wire1589/A vssd vccd _614_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_27_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__473__A_N _601_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__266__A _266_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_324_ _324_/A _324_/B vssd vccd _324_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_255_ _255_/A _255_/B vssd vccd _255_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_186_ _186_/A _186_/B vssd vccd _186_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_7_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__432__C _432_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3076 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1245_A _340_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1412_A wire1413/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__176__A _176_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1781_A wire1781/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1879_A wire1880/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__623__B _623_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4471 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[4\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_4379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1563 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__496__A_N _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1162 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__086__A _086_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_862 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_040_ _040_/A vssd vccd _040_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2095_A wire2096/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input178_A la_iena_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input345_A la_oenb_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2010 wire2011/X vssd vccd _569_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2021 wire2021/A vssd vccd _560_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2032 wire2032/A vssd vccd _518_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_out_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2043 wire2043/A vssd vccd wire2043/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2054 wire2054/A vssd vccd wire2054/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1320 _257_/X vssd vccd wire1320/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2065 wire2065/A vssd vccd wire2065/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2076 wire2077/X vssd vccd _493_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1331 _246_/X vssd vccd wire1331/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1342 wire1343/X vssd vccd _299_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2087 wire2087/A vssd vccd wire2087/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1353 wire1353/A vssd vccd wire1353/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2098 wire2098/A vssd vccd wire2098/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1364 wire1364/A vssd vccd _364_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1375 wire1375/A vssd vccd _356_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1386 wire1386/A vssd vccd wire1386/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1397 wire1397/A vssd vccd wire1397/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__427__C _427_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3972 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_307_ _307_/A _307_/B vssd vccd _307_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_238_ _238_/A _238_/B vssd vccd _238_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__443__B _443_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output564_A _445_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__369__A_N _497_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_169_ _169_/A _169_/B vssd vccd _169_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_7_796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1195_A wire1196/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output731_A _607_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output829_A _581_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3932 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] _239_/X vssd vccd _059_/A vssd vccd
+ sky130_fd_sc_hd__nand2_8
XFILLER_23_3976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1627_A wire1627/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__618__B _618_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1996_A wire1997/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__353__B _353_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1966 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput306 la_oenb_mprj[26] vssd vccd _523_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput317 la_oenb_mprj[36] vssd vccd _405_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput328 la_oenb_mprj[46] vssd vccd _415_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput339 la_oenb_mprj[56] vssd vccd _553_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_22_3464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1382 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3475 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2846 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1038 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__528__B _528_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2010_A wire2011/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2108_A wire2109/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__544__A _544_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input295_A la_oenb_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__263__B _263_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_023_ _023_/A vssd vccd _023_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_input462_A user_irq_ena[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_4087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2663 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3002 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1150 wire1151/X vssd vccd wire1150/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1161 _365_/X vssd vccd wire1161/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1172 wire1173/X vssd vccd wire1172/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1183 wire1184/X vssd vccd wire1183/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1194 wire1195/X vssd vccd wire1194/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__438__B _438_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1110_A _403_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1208_A wire1209/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3791 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output779_A wire1019/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_2678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output946_A wire1289/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1577_A wire1578/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1744_A wire1745/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1911_A wire1912/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] _265_/X vssd vccd _085_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XANTENNA__348__B _348_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__364__A _364_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3300 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput103 la_data_out_mprj[74] vssd vccd wire1630/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput114 la_data_out_mprj[84] vssd vccd wire1620/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_49_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput125 la_data_out_mprj[94] vssd vccd _463_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_27_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput136 la_iena_mprj[103] vssd vccd _266_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput147 la_iena_mprj[113] vssd vccd _276_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput158 la_iena_mprj[123] vssd vccd _286_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput169 la_iena_mprj[18] vssd vccd _181_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire2058_A wire2059/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__539__A _539_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input210_A la_iena_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_572_ _572_/A _572_/B vssd vccd _572_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_29_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_648 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input308_A la_oenb_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2342 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__274__A _274_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_186 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_006_ _006_/A vssd vccd _006_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_3459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__440__C _440_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__A_N _535_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2471 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3288 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output527_A wire1102/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1060_A _475_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1158_A wire1159/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1325_A _252_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output896_A _137_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_0 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] _202_/X vssd vccd _022_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__184__A _184_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4186 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1694_A wire1695/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1015 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1195 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1861_A wire1861/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1959_A wire1960/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1059 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1908 wire1909/X vssd vccd _613_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1919 wire1920/X vssd vccd _610_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2930 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__359__A _359_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_208 _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_219 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__094__A _094_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input160_A la_iena_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input258_A la_iena_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2175_A wire2176/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4079 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input425_A mprj_dat_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input21_A la_data_out_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__269__A _269_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_624_ _624_/A _624_/B vssd vccd _624_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_555_ _555_/A _555_/B vssd vccd _555_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_486_ _614_/A _486_/B _486_/C vssd vccd _486_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_18_2459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__435__C _435_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4007 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output477_A wire1054/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__451__B _451_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output644_A _015_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1275_A _314_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output811_A _565_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2290 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1442_A wire1443/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__179__A _179_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3776 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_702 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__361__B _361_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput930 wire1170/X vssd vccd mprj_dat_o_user[25] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput941 wire1235/X vssd vccd mprj_dat_o_user[6] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput952 output952/A vssd vccd user1_vdd_powergood vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1447 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1705 wire1705/A vssd vccd wire1705/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1716 wire1716/A vssd vccd _353_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1727 wire1728/X vssd vccd wire1727/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__089__A _089_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1738 wire1739/X vssd vccd _289_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1749 wire1750/X vssd vccd _284_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2771 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_340_ _340_/A _340_/B vssd vccd _340_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__536__B _536_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_271_ _271_/A _271_/B vssd vccd _271_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__552__A _552_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input375_A la_oenb_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__271__B _271_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_4040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input69_A la_data_out_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_607_ _607_/A _607_/B vssd vccd _607_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_45_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__B _446_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_538_ _538_/A _538_/B vssd vccd _538_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_50_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output594_A _085_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_469_ _597_/A _469_/B _469_/C vssd vccd _469_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_32_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output761_A wire1030/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output859_A _306_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1392_A wire1393/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__181__B _181_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3136 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1657_A wire1658/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2374 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__356__B _356_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_4056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[94\]_B wire1320/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3738 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1298 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput760 wire1031/X vssd vccd la_oenb_core[21] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3440 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput771 _528_/X vssd vccd la_oenb_core[31] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput782 wire1018/X vssd vccd la_oenb_core[41] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_1211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2203 wire2204/X vssd vccd _295_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput793 _548_/X vssd vccd la_oenb_core[51] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1502 wire1503/X vssd vccd wire1502/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1513 wire1514/X vssd vccd wire1513/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1524 wire1525/X vssd vccd wire1524/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1535 wire1535/A vssd vccd _579_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1546 wire1546/A vssd vccd _568_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1557 input34/X vssd vccd _496_/C vssd vccd sky130_fd_sc_hd__buf_4
Xwire1568 _405_/A_N vssd vccd _533_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1579 wire1579/A vssd vccd _624_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input123_A la_data_out_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2040_A wire2041/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2138_A wire2138/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__547__A _547_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__266__B _266_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_323_ _323_/A _323_/B vssd vccd _323_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_1132 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_B wire1329/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_254_ _254_/A _254_/B vssd vccd _254_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__282__A _282_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_185_ _185_/A _185_/B vssd vccd _185_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_45_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[4\] mprj_dat_i_user[4] max_length1311/X vssd vccd _118_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_6_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1140_A _374_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1238_A wire1239/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3907 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1405_A wire1406/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] _184_/X vssd vccd _004_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
XFILLER_15_3675 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_B _239_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3528 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__A _192_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1774_A wire1774/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1941_A wire1942/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4408 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1575 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3668 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4187 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__367__A _367_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3535 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2088_A wire2089/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2000 wire2000/A vssd vccd wire2000/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput590 wire1136/X vssd vccd la_data_in_core[9] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2011 wire2011/A vssd vccd wire2011/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire2022 wire2022/A vssd vccd _559_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input240_A la_iena_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2033 wire2033/A vssd vccd _517_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input338_A la_oenb_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2044 wire2044/A vssd vccd _509_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2400 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2055 wire2056/X vssd vccd _502_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__440__A_N _568_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1321 _256_/X vssd vccd wire1321/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2066 wire2067/X vssd vccd _496_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2077 wire2078/X vssd vccd wire2077/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1332 _243_/X vssd vccd wire1332/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1343 wire1343/A vssd vccd wire1343/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2088 wire2089/X vssd vccd _489_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2099 wire2100/X vssd vccd _485_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1354 wire1355/X vssd vccd _341_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1365 wire1365/A vssd vccd _363_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1376 wire1376/A vssd vccd _355_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1387 wire1388/X vssd vccd _348_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1398 wire1399/X vssd vccd _314_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__277__A _277_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_370 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_306_ _306_/A _306_/B vssd vccd _306_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_237_ _237_/A _237_/B vssd vccd _237_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__443__C _443_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_742 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_168_ _168_/A _168_/B vssd vccd _168_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_13_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output557_A wire1139/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_099_ _099_/A vssd vccd _099_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_wire1090_A _422_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1188_A wire1189/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output724_A _601_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2416 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3944 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1355_A wire1355/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3988 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] _232_/X vssd vccd _052_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1522_A wire1523/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__187__A _187_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1891_A wire1891/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1989_A wire1989/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3916 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__463__A_N _591_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput307 la_oenb_mprj[27] vssd vccd wire1575/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput318 la_oenb_mprj[37] vssd vccd _406_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput329 la_oenb_mprj[47] vssd vccd _416_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_3695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2803 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__097__A _097_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[124\]_B wire1312/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__544__B _544_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2003_A wire2004/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1758 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input190_A la_iena_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input288_A la_oenb_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_022_ _022_/A vssd vccd _022_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_6_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_712 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__A _560_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input455_A mprj_sel_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input51_A la_data_out_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2675 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_962 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1140 _374_/X vssd vccd wire1140/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1151 wire1152/X vssd vccd wire1151/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1162 wire1163/X vssd vccd wire1162/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1173 _362_/X vssd vccd wire1173/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1184 wire1185/X vssd vccd wire1184/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1195 wire1196/X vssd vccd wire1195/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__438__C _438_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__454__B _454_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[115\]_B _278_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1103_A _410_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3082 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__486__A_N _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output841_A _592_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output939_A wire1241/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1472_A wire1473/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3752 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1904_A wire1904/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[24\]_A mprj_dat_i_user[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_660 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[106\]_B _269_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__364__B _364_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2167 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput104 la_data_out_mprj[75] vssd vccd wire1629/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput115 la_data_out_mprj[85] vssd vccd wire1619/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput126 la_data_out_mprj[95] vssd vccd _464_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput137 la_iena_mprj[104] vssd vccd _267_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput148 la_iena_mprj[114] vssd vccd _277_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput159 la_iena_mprj[124] vssd vccd _287_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__539__B _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[15\]_A mprj_dat_i_user[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_571_ _571_/A _571_/B vssd vccd _571_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2120_A wire2120/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input203_A la_iena_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__555__A _555_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__274__B _274_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input99_A la_data_out_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_3976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__A _290_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_005_ _005_/A vssd vccd _005_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_21_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__B _449_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1053_A _497_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_958 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4408 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1220_A wire1221/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output791_A wire1049/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_1 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1318_A _259_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1687_A wire1687/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1854_A wire1855/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_2319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2258 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1909 wire1910/X vssd vccd wire1909/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_39_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__359__B _359_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_209 _232_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1864 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2070_A wire2071/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input153_A la_iena_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2168_A wire2168/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__269__B _269_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input320_A la_oenb_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input418_A mprj_adr_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_623_ _623_/A _623_/B vssd vccd _623_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_2391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input14_A la_data_out_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_554_ _554_/A _554_/B vssd vccd _554_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1795 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__285__A _285_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_485_ _613_/A _485_/B _485_/C vssd vccd _485_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2086 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4019 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__451__C _451_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2639 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output637_A _009_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1170_A wire1171/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1268_A wire1269/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output804_A wire996/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1435_A wire1436/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] _214_/X vssd vccd _034_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_714 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__195__A _195_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1214 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1971_A wire1971/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2000 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput920 wire1205/X vssd vccd mprj_dat_o_user[16] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput931 wire1166/X vssd vccd mprj_dat_o_user[26] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput942 wire1232/X vssd vccd mprj_dat_o_user[7] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_2116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput953 wire2205/X vssd vccd user2_vcc_powergood vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input6_A la_data_out_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1706 wire1707/X vssd vccd _361_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1717 wire1717/A vssd vccd _352_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1728 wire1728/A vssd vccd wire1728/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1739 wire1739/A vssd vccd wire1739/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_270_ _270_/A _270_/B vssd vccd _270_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_3902 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__552__B _552_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input270_A la_oenb_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input368_A la_oenb_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3290 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_606_ _606_/A _606_/B vssd vccd _606_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_37_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_91 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_537_ _537_/A _537_/B vssd vccd _537_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__446__C _446_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_468_ _596_/A _468_/B _468_/C vssd vccd _468_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_wire1016_A wire1017/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output587_A wire1069/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_399_ _527_/A _399_/B _399_/C vssd vccd _399_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_31_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1111 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__B _462_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output754_A wire1036/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1385_A wire1386/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3148 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output921_A wire1202/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] wire1317/X vssd vccd wire961/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_29_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3530 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1817_A wire1817/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_791 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__372__B _372_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2980 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[7\]_A mprj_dat_i_user[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_4131 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3502 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput750 wire1040/X vssd vccd la_oenb_core[12] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput761 wire1030/X vssd vccd la_oenb_core[22] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput772 _529_/X vssd vccd la_oenb_core[32] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput783 wire1016/X vssd vccd la_oenb_core[42] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2204 wire2204/A vssd vccd wire2204/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput794 wire1007/X vssd vccd la_oenb_core[52] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1223 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2030 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1503 wire1504/X vssd vccd wire1503/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1514 wire1514/A vssd vccd wire1514/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1525 wire1526/X vssd vccd wire1525/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1536 wire1536/A vssd vccd _578_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1547 wire1547/A vssd vccd _567_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1558 _420_/A_N vssd vccd _548_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1569 wire1569/A vssd vccd _532_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_27_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__547__B _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input116_A la_data_out_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2033_A wire2033/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_2511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_322_ _322_/A _322_/B vssd vccd _322_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire2200_A wire2200/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__563__A _563_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_253_ _253_/A _253_/B vssd vccd _253_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_975 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input81_A la_data_out_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_184_ _184_/A _184_/B vssd vccd _184_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3238 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output502_A wire1144/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__457__B _457_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1133_A wire1134/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_4491 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1300_A wire1301/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output871_A _335_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] _177_/X vssd vccd _161_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_2210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[27\] mprj_dat_i_user[27] _294_/X vssd vccd _141_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_33_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__192__B _192_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1767_A wire1768/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4440 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4495 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1934_A wire1935/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3636 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] _288_/X vssd vccd _108_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_9_1587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__367__B _367_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__A_N _520_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2608 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3547 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput580 wire1076/X vssd vccd la_data_in_core[90] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2001 wire2002/X vssd vccd _574_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_3271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput591 _147_/Y vssd vccd la_data_in_mprj[0] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2012 wire2013/X vssd vccd _568_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_27_2879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2023 wire2023/A vssd vccd _546_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_8_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2034 wire2034/A vssd vccd _516_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1300 wire1301/X vssd vccd wire1300/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2045 wire2046/X vssd vccd _508_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2056 wire2056/A vssd vccd wire2056/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1322 _255_/X vssd vccd wire1322/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire2067 wire2068/X vssd vccd wire2067/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2150_A wire2151/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input233_A la_iena_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2078 wire2078/A vssd vccd wire2078/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1333 _242_/X vssd vccd wire1333/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1344 wire1345/X vssd vccd _346_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2089 wire2090/X vssd vccd wire2089/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__558__A _558_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1355 wire1355/A vssd vccd wire1355/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1366 wire1366/A vssd vccd _362_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1377 wire1377/A vssd vccd _354_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1388 wire1388/A vssd vccd wire1388/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1399 wire1400/X vssd vccd wire1399/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input400_A mprj_adr_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__277__B _277_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__293__A _293_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_305_ _305_/A _305_/B vssd vccd _305_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4252 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_236_ _236_/A _236_/B vssd vccd _236_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_167_ _167_/A _167_/B vssd vccd _167_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_48_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_098_ _098_/A vssd vccd _098_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_26_3024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1083_A _427_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3956 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output717_A _082_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1250_A _338_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1348_A wire1349/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__187__B _187_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1515_A wire1516/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3304 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1884_A wire1885/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire968_A wire968/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3928 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput308 la_oenb_mprj[28] vssd vccd _525_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_9_2074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput319 la_oenb_mprj[38] vssd vccd _535_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1351 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1395 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2859 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3106 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_021_ _021_/A vssd vccd _021_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input183_A la_iena_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1423 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__560__B _560_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input350_A la_oenb_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input448_A mprj_dat_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3399 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input44_A la_data_out_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1130 _383_/X vssd vccd wire1130/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__288__A _288_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1141 _373_/X vssd vccd wire1141/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1152 wire1153/X vssd vccd wire1152/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1163 wire1164/X vssd vccd wire1163/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1174 wire1175/X vssd vccd wire1174/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1185 _359_/X vssd vccd wire1185/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1196 wire1197/X vssd vccd wire1196/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_628 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__454__C _454_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3094 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_219_ _219_/A _219_/B vssd vccd _219_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1298_A _301_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__470__B _470_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output834_A wire995/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2691 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1465_A wire1466/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] _244_/X vssd vccd wire975/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_3_3803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__198__A _198_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_606 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[24\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_672 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2747 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__430__A_N _558_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3178 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__380__B _380_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3471 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput105 la_data_out_mprj[76] vssd vccd wire1628/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput116 la_data_out_mprj[86] vssd vccd wire1618/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput127 la_data_out_mprj[96] vssd vccd _465_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput138 la_iena_mprj[105] vssd vccd _268_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput149 la_iena_mprj[115] vssd vccd _278_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_2551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[15\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_570_ _570_/A _570_/B vssd vccd _570_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1966 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__555__B _555_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2113_A wire2114/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input398_A mprj_adr_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3988 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__571__A _571_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_004_ _004_/A vssd vccd _004_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_46_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__290__B _290_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1800 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2495 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__C _449_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1046_A _504_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_2 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__465__B _465_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1213_A _351_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__453__A_N _581_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_4122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output784_A _540_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_4133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output951_A wire1723/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2791 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1847_A wire1848/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4356 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4378 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__375__B _375_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1810 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4015 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2063_A wire2063/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input146_A la_iena_mprj[112] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_622_ _622_/A _622_/B vssd vccd _622_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_2381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input313_A la_oenb_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__476__A_N _604_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__566__A _566_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_553_ _553_/A _553_/B vssd vccd _553_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_18_2406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4008 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__285__B _285_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_484_ _612_/A _484_/B _484_/C vssd vccd _484_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2098 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output532_A wire1097/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1163_A wire1164/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1330_A _247_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1428_A wire1429/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] _207_/X vssd vccd _027_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_4364 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1797_A wire1797/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1964_A wire1964/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput910 _121_/Y vssd vccd mprj_dat_i_core[7] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput921 wire1202/X vssd vccd mprj_dat_o_user[17] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput932 wire1162/X vssd vccd mprj_dat_o_user[27] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput943 wire1229/X vssd vccd mprj_dat_o_user[8] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3864 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] _169_/X vssd vccd _153_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_25_2900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput954 output954/A vssd vccd user2_vdd_powergood vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_3_4120 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1707 wire1707/A vssd vccd wire1707/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1718 wire1718/A vssd vccd _351_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1729 wire1730/X vssd vccd _292_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_767 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input263_A la_oenb_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2180_A wire2181/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3238 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input430_A mprj_dat_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__296__A _296_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4504 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_605_ _605_/A _605_/B vssd vccd _605_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_45_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_704 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_536_ _536_/A _536_/B vssd vccd _536_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_15_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_467_ _595_/A _467_/B _467_/C vssd vccd _467_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_14_962 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_398_ _526_/A _398_/B _398_/C vssd vccd _398_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output482_A _486_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1009_A wire1010/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__462__C _462_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output747_A _622_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1280_A wire1281/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1378_A wire1378/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output914_A wire1223/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3818 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1712_A wire1712/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4014 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[7\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2992 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput740 _616_/X vssd vccd la_oenb_core[119] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput751 wire1039/X vssd vccd la_oenb_core[13] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput762 wire1029/X vssd vccd la_oenb_core[23] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3514 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput773 wire1024/X vssd vccd la_oenb_core[33] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput784 _540_/X vssd vccd la_oenb_core[43] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2205 wire2206/X vssd vccd wire2205/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput795 wire1005/X vssd vccd la_oenb_core[53] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1504 wire1504/A vssd vccd wire1504/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2042 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1515 wire1516/X vssd vccd _317_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1526 wire1526/A vssd vccd wire1526/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1537 wire1537/A vssd vccd _577_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1279 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[7\]_B _170_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1548 wire1548/A vssd vccd _566_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1559 _417_/A_N vssd vccd _545_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_3224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2026_A wire2026/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input109_A la_data_out_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_321_ _321_/A _321_/B vssd vccd _321_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_252_ _252_/A _252_/B vssd vccd _252_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__563__B _563_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1156 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_183_ _183_/A _183_/B vssd vccd _183_/X vssd vccd sky130_fd_sc_hd__and2_1
XANTENNA_input380_A la_oenb_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input74_A la_data_out_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__C _457_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1126_A _387_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_360 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_519_ _519_/A _519_/B vssd vccd _519_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__473__B _473_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output864_A _329_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1495_A wire1496/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1662_A wire1662/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1927_A wire1927/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3648 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4084 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3580 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] _281_/X vssd vccd _101_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_3_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3488 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3290 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__383__B _383_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3559 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput570 _450_/X vssd vccd la_data_in_core[81] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput581 wire1075/X vssd vccd la_data_in_core[91] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2002 wire2002/A vssd vccd wire2002/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput592 _083_/Y vssd vccd la_data_in_mprj[100] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2013 wire2013/A vssd vccd wire2013/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2024 wire2024/A vssd vccd _539_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_43_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2035 wire2035/A vssd vccd _515_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1301 wire1302/X vssd vccd wire1301/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2046 wire2046/A vssd vccd wire2046/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1312 _287_/X vssd vccd wire1312/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire2057 wire2057/A vssd vccd _501_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2068 wire2068/A vssd vccd wire2068/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1323 _254_/X vssd vccd wire1323/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1334 input99/X vssd vccd _439_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire2079 wire2080/X vssd vccd _492_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1087 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1345 wire1345/A vssd vccd wire1345/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__558__B _558_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1356 wire1357/X vssd vccd _340_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2143_A wire2143/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input226_A la_iena_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1367 wire1367/A vssd vccd _361_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1378 wire1378/A vssd vccd _353_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1389 wire1390/X vssd vccd _347_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__574__A _574_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3855 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__293__B _293_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_4220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_304_ _304_/A _304_/B vssd vccd _304_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4264 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_235_ _235_/A _235_/B vssd vccd _235_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_166_ _166_/A _166_/B vssd vccd _166_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_097_ _097_/A vssd vccd _097_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1076_A _459_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__468__B _468_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1890 wire1891/X vssd vccd wire1890/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_106 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1410_A wire1411/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1508_A wire1508/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA_190 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3316 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1638 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1877_A wire1878/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4310 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4102 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput309 la_oenb_mprj[29] vssd vccd wire1574/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1363 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__B _378_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3118 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_16_2515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_150 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_020_ _020_/A vssd vccd _020_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_14_2283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1435 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2093_A wire2093/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input176_A la_iena_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input343_A la_oenb_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__569__A _569_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2699 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input37_A la_data_out_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1120 _393_/X vssd vccd wire1120/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1131 _382_/X vssd vccd wire1131/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__288__B _288_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1142 _372_/X vssd vccd wire1142/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1153 _367_/X vssd vccd wire1153/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1164 wire1165/X vssd vccd wire1164/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1175 wire1176/X vssd vccd wire1175/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1186 wire1187/X vssd vccd wire1186/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1197 _356_/X vssd vccd wire1197/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4495 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_218_ _218_/A _218_/B vssd vccd _218_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_45_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output562_A _443_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_149_ _149_/A vssd vccd _149_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__470__C _470_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output827_A _579_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__382__A_N _510_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1008 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1360_A wire1361/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1458_A wire1459/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] _237_/X vssd vccd _057_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_3848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1625_A wire1625/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3427 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1994_A wire1995/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_684 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1446 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__380__C _380_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3704 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3507 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3748 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput106 la_data_out_mprj[77] vssd vccd wire1627/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput117 la_data_out_mprj[87] vssd vccd wire1617/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput128 la_data_out_mprj[97] vssd vccd _466_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput139 la_iena_mprj[106] vssd vccd _269_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2635 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2106_A wire2107/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1546 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input293_A la_oenb_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__571__B _571_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3680 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_90 mprj_dat_i_user[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_003_ _003_/A vssd vccd _003_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input460_A user_irq_ena[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__299__A _299_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3916 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1039_A _510_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_3 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1206_A wire1207/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3422 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output777_A _534_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1608 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__481__B _481_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output944_A wire1226/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1742_A wire1743/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2900 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__002__A _002_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_938 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] _263_/X vssd vccd wire993/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_39_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4056 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_131 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__391__B _391_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_4027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2750 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input139_A la_iena_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2056_A wire2056/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_621_ _621_/A _621_/B vssd vccd _621_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1720 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1742 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_552_ _552_/A _552_/B vssd vccd _552_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__566__B _566_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input306_A la_oenb_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_483_ _611_/A _483_/B _483_/C vssd vccd _483_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_44_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__A _582_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_3077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output525_A wire1104/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1156_A wire1157/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__420__A_N _420_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__476__B _476_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1323_A _254_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4376 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output894_A _135_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] _200_/X vssd vccd _020_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1692_A wire1693/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1957_A wire1958/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput900 _141_/Y vssd vccd mprj_dat_i_core[27] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput911 _122_/Y vssd vccd mprj_dat_i_core[8] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput922 wire1198/X vssd vccd mprj_dat_o_user[18] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput933 wire1158/X vssd vccd mprj_dat_o_user[28] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput944 wire1226/X vssd vccd mprj_dat_o_user[9] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput955 wire1307/X vssd vccd user_clock vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3707 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[30\]_B _193_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_4176 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1708 wire1708/A vssd vccd _360_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1719 wire1719/A vssd vccd _350_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_45_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__386__B _386_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_B _260_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2630 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2173_A wire2174/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input256_A la_iena_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__443__A_N _571_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input423_A mprj_dat_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__577__A _577_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_604_ _604_/A _604_/B vssd vccd _604_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_15_4516 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3962 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_716 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_535_ _535_/A _535_/B vssd vccd _535_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[88\]_B wire1326/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_466_ _594_/A _466_/B _466_/C vssd vccd _466_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_53_1438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_397_ _525_/A _397_/B _397_/C vssd vccd _397_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output475_A wire1056/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3911 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output642_A _013_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3955 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1273_A _315_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1440_A wire1441/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1538_A wire1538/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2195 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_4075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B wire1333/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__466__A_N _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput730 wire1042/X vssd vccd la_oenb_core[10] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3651 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput741 wire1041/X vssd vccd la_oenb_core[11] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput752 wire1038/X vssd vccd la_oenb_core[14] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput763 wire1028/X vssd vccd la_oenb_core[24] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput774 wire1022/X vssd vccd la_oenb_core[34] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput785 wire1015/X vssd vccd la_oenb_core[44] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2206 wire2207/X vssd vccd wire2206/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput796 _551_/X vssd vccd la_oenb_core[54] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1505 wire1506/X vssd vccd _320_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1516 wire1517/X vssd vccd wire1516/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2054 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1527 wire1527/A vssd vccd _596_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1538 wire1538/A vssd vccd _576_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1549 wire1549/A vssd vccd _565_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_320_ _320_/A _320_/B vssd vccd _320_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_42_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2019_A wire2019/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_251_ _251_/A _251_/B vssd vccd _251_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_270 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3892 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_182_ _182_/A _182_/B vssd vccd _182_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_49_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input373_A la_oenb_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input67_A la_data_out_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__100__A _100_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_350 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_361 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_518_ _518_/A _518_/B vssd vccd _518_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_50_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output592_A _083_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1119_A _394_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_449_ _577_/A _449_/B _449_/C vssd vccd _449_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__489__A_N _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output857_A _323_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1488_A wire1489/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1655_A wire1656/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1534 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1359 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__383__C _383_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2590 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput560 _441_/X vssd vccd la_data_in_core[72] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput571 _451_/X vssd vccd la_data_in_core[82] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput582 wire1074/X vssd vccd la_data_in_core[92] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2003 wire2004/X vssd vccd _573_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput593 _084_/Y vssd vccd la_data_in_mprj[101] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_1011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire2014 wire2014/A vssd vccd _567_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_1573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2025 wire2025/A vssd vccd _535_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire2036 wire2036/A vssd vccd _514_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2047 wire2048/X vssd vccd _507_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1302 _300_/X vssd vccd wire1302/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1055 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2058 wire2059/X vssd vccd _500_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1313 _286_/X vssd vccd wire1313/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2069 wire2070/X vssd vccd _495_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1324 _253_/X vssd vccd wire1324/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_2583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1335 input97/X vssd vccd _438_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1099 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1346 wire1347/X vssd vccd _345_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1357 wire1357/A vssd vccd wire1357/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1368 wire1368/A vssd vccd _360_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1379 wire1380/X vssd vccd _352_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input121_A la_data_out_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input219_A la_iena_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2136_A wire2136/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__574__B _574_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[127\]_B _290_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_303_ _303_/A _303_/B vssd vccd _303_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_19_2398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_234_ _234_/A _234_/B vssd vccd _234_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_7_712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__A _590_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_165_ _165_/A _165_/B vssd vccd _165_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_767 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[2\] mprj_dat_i_user[2] max_length1310/X vssd vccd _116_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
X_096_ _096_/A vssd vccd _096_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_powergood_check_mprj_vdd_logic1 output952/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_940 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__468__C _468_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output605_A _095_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1880 wire1881/X vssd vccd wire1880/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1236_A wire1237/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1891 wire1891/A vssd vccd wire1891/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__484__B _484_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_B _281_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1403_A wire1404/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_180 _358_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_191 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1772_A wire1772/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4322 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__005__A _005_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1270 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[27\]_A mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__C _378_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__B _394_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[109\]_B _272_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1447 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2086_A wire2087/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input169_A la_iena_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__569__B _569_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input336_A la_oenb_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[18\]_A mprj_dat_i_user[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1110 _403_/X vssd vccd wire1110/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1121 _392_/X vssd vccd wire1121/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1132 _381_/X vssd vccd wire1132/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1143 _371_/X vssd vccd wire1143/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1154 wire1155/X vssd vccd wire1154/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_2316 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1165 _364_/X vssd vccd wire1165/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1176 wire1177/X vssd vccd wire1176/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1187 wire1188/X vssd vccd wire1187/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1198 wire1199/X vssd vccd wire1198/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_53_3907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__585__A _585_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4327 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_217_ _217_/A _217_/B vssd vccd _217_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_4084 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_148_ _148_/A vssd vccd _148_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_1071 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output555_A _437_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_079_ _079_/A vssd vccd _079_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1186_A wire1187/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output722_A _599_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__479__B _479_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1353_A wire1353/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4180 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] _230_/X vssd vccd _050_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1520_A wire1521/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1618_A wire1618/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1804 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_696 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1987_A wire1987/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire973_A wire973/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3294 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3519 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4091 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput107 la_data_out_mprj[78] vssd vccd wire1626/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput118 la_data_out_mprj[88] vssd vccd wire1616/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__389__B _389_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2750 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput129 la_data_out_mprj[98] vssd vccd _467_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1183 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_630 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2001_A wire2002/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1558 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input286_A la_oenb_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_80 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_002_ _002_/A vssd vccd _002_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_11_3692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_91 mprj_dat_i_user[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1391 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input453_A mprj_iena_wb vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__299__B _299_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3928 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_4 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1101_A _412_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__481__C _481_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output937_A wire1146/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1470_A wire1471/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1568_A _405_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1735_A wire1736/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3596 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1902_A wire1903/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4039 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3579 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_620_ _620_/A _620_/B vssd vccd _620_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_2361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2049_A wire2050/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_551_ _551_/A _551_/B vssd vccd _551_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_45_747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input201_A la_iena_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_482_ _610_/A _482_/B _482_/C vssd vccd _482_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_38_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__372__A_N _500_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__582__B _582_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input97_A la_data_out_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__103__A _103_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_570 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3758 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output518_A wire1110/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput460 user_irq_ena[0] vssd vccd _291_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1051_A _499_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3632 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__492__B _492_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3242 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1685_A wire1685/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3800 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput901 _142_/Y vssd vccd mprj_dat_i_core[28] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput912 _123_/Y vssd vccd mprj_dat_i_core[9] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1852_A wire1853/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput923 wire1194/X vssd vccd mprj_dat_o_user[19] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput934 wire1154/X vssd vccd mprj_dat_o_user[29] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput945 wire1294/X vssd vccd mprj_sel_o_user[0] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput956 _297_/X vssd vccd user_clock2 vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1709 wire1709/A vssd vccd _359_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_2979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2720 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__386__C _386_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__395__A_N _523_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2327 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2642 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input151_A la_iena_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2166_A wire2166/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input249_A la_iena_mprj[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__577__B _577_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input416_A mprj_adr_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_603_ _603_/A _603_/B vssd vccd _603_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input12_A la_data_out_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1551 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_534_ _534_/A _534_/B vssd vccd _534_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_15_4528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__593__A _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_465_ _593_/A _465_/B _465_/C vssd vccd _465_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_975 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_396_ _524_/A _396_/B _396_/C vssd vccd _396_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_3551 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1158 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output468_A wire1062/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1099_A _414_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3923 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2428 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3967 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output635_A _007_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1266_A wire1267/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output802_A wire1048/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__487__B _487_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1433_A wire1434/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput290 la_oenb_mprj[127] vssd vccd wire1579/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1003 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__008__A _008_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput720 _597_/X vssd vccd la_oenb_core[100] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput731 _607_/X vssd vccd la_oenb_core[110] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput742 _617_/X vssd vccd la_oenb_core[120] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3663 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4167 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput753 wire1037/X vssd vccd la_oenb_core[15] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput764 wire1027/X vssd vccd la_oenb_core[25] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput775 _532_/X vssd vccd la_oenb_core[35] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput786 wire1013/X vssd vccd la_oenb_core[45] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2207 wire2208/X vssd vccd wire2207/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput797 wire1004/X vssd vccd la_oenb_core[55] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input4_A la_data_out_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1506 wire1507/X vssd vccd wire1506/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2607 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1517 wire1517/A vssd vccd wire1517/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1528 wire1528/A vssd vccd _595_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1539 wire1539/A vssd vccd _575_/A vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__397__B _397_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3204 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_250_ _250_/A _250_/B vssd vccd _250_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_1125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2282 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_282 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_181_ _181_/A _181_/B vssd vccd _181_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_52_1450 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input199_A la_iena_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__410__A_N _538_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input366_A la_oenb_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_irq_gates\[1\] user_irq_core[1] _292_/X vssd vccd _112_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_43_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__588__A _588_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3864 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_340 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_351 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_517_ _517_/A _517_/B vssd vccd _517_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_362 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_448_ _576_/A _448_/B _448_/C vssd vccd _448_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output585_A wire1071/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3370 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_379_ _507_/A _379_/B _379_/C vssd vccd _379_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output752_A wire1038/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1383_A wire1384/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3731 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] _260_/X vssd vccd _080_/A vssd vccd
+ sky130_fd_sc_hd__nand2_8
XFILLER_6_3825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2247 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1648_A wire1649/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4103 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__A _498_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__A_N _561_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput550 _432_/X vssd vccd la_data_in_core[63] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput561 _442_/X vssd vccd la_data_in_core[73] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_27_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput572 _452_/X vssd vccd la_data_in_core[83] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput583 wire1073/X vssd vccd la_data_in_core[93] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2004 wire2004/A vssd vccd wire2004/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput594 _085_/Y vssd vccd la_data_in_mprj[102] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2015 wire2015/A vssd vccd _566_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2026 wire2026/A vssd vccd _531_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2037 wire2038/X vssd vccd _513_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2551 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1303 wire1304/X vssd vccd wire1303/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2048 wire2048/A vssd vccd wire2048/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1067 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__201__A _201_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2059 wire2059/A vssd vccd wire2059/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2415 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1314 _277_/X vssd vccd wire1314/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1325 _252_/X vssd vccd wire1325/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_2595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1336 input96/X vssd vccd _437_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1347 wire1347/A vssd vccd wire1347/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1358 wire1358/A vssd vccd _368_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1369 wire1369/A vssd vccd _359_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2031_A wire2031/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input114_A la_data_out_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2129_A wire2129/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_302_ _302_/A _302_/B vssd vccd _302_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_42_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_233_ _233_/A _233_/B vssd vccd _233_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__590__B _590_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_164_ _164_/A _164_/B vssd vccd _164_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_7_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_095_ _095_/A vssd vccd _095_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4362 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1870 wire1870/A vssd vccd wire1870/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_output500_A wire1126/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1881 wire1882/X vssd vccd wire1881/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1892 wire1893/X vssd vccd _618_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4100 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1131_A _382_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1229_A wire1230/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__456__A_N _584_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__C _484_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_170 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_181 _358_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_192 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] _175_/X vssd vccd _159_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[25\] mprj_dat_i_user[25] _294_/X vssd vccd _139_/A vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1006 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_2639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1765_A wire1766/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1932_A wire1933/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1282 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__021__A _021_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[27\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] wire1313/X vssd vccd wire981/A
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_2_2818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2079_A wire2080/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1100 _413_/X vssd vccd wire1100/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[18\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1111 _402_/X vssd vccd wire1111/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1122 _391_/X vssd vccd wire1122/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input231_A la_iena_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1133 wire1134/X vssd vccd wire1133/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input329_A la_oenb_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__479__A_N _479_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1144 _370_/X vssd vccd wire1144/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1155 wire1156/X vssd vccd wire1155/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1166 wire1167/X vssd vccd wire1166/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1177 _361_/X vssd vccd wire1177/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1188 wire1189/X vssd vccd wire1188/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1199 wire1200/X vssd vccd wire1199/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__585__B _585_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3638 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_216_ _216_/A _216_/B vssd vccd _216_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_11_594 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4096 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__106__A _106_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_147_ _147_/A vssd vccd _147_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_1050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1083 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_078_ _078_/A vssd vccd _078_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output548_A wire1079/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1081_A _428_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1179_A wire1180/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__479__C _479_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output715_A _080_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1346_A wire1347/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3596 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__B _495_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1513_A wire1514/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1816 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1882_A wire1882/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_2414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire966_A wire966/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__016__A _016_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput108 la_data_out_mprj[79] vssd vccd wire1625/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__389__C _389_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput119 la_data_out_mprj[89] vssd vccd _458_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1195 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_642 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_70 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_001_ _001_/A vssd vccd _001_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_81 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_92 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input181_A la_iena_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2196_A wire2196/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input279_A la_oenb_mprj[117] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1223 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3111 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input446_A mprj_dat_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input42_A la_data_out_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__596__A _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_5 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output498_A wire1128/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1296_A wire1297/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output832_A _584_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1463_A wire1464/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_4337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1630_A wire1630/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1728_A wire1728/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput90 la_data_out_mprj[62] vssd vccd _431_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_550_ _550_/A _550_/B vssd vccd _550_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_17_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_940 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_481_ _609_/A _481_/B _481_/C vssd vccd _481_/X vssd vccd sky130_fd_sc_hd__and3b_1
XFILLER_16_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2111_A wire2111/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2209_A wire2209/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input396_A mprj_adr_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput450 mprj_dat_o_core[7] vssd vccd wire1349/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput461 user_irq_ena[1] vssd vccd _292_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2091 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1044_A _506_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3644 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1211_A wire1212/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4091 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output782_A wire1018/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1309_A _296_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__492__C _492_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3254 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1678_A wire1679/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput902 _143_/Y vssd vccd mprj_dat_i_core[29] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput913 wire1251/X vssd vccd mprj_dat_o_user[0] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput924 wire1249/X vssd vccd mprj_dat_o_user[1] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput935 wire1246/X vssd vccd mprj_dat_o_user[2] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3615 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput946 wire1289/X vssd vccd mprj_sel_o_user[1] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput957 _111_/Y vssd vccd user_irq[0] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_7_4270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1845_A wire1845/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3372 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2732 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_442 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2339 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__204__A _204_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3388 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2518 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3090 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input144_A la_iena_mprj[110] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2061_A wire2061/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2159_A wire2160/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_602_ _602_/A _602_/B vssd vccd _602_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input311_A la_oenb_mprj[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input409_A mprj_adr_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_533_ _533_/A _533_/B vssd vccd _533_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_1563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1574 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__593__B _593_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_464_ _592_/A _464_/B _464_/C vssd vccd _464_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_395_ _523_/A _395_/B _395_/C vssd vccd _395_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3596 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3935 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3979 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output530_A wire1099/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1161_A _365_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1259_A _322_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__487__C _487_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3567 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput280 la_oenb_mprj[118] vssd vccd wire1588/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput291 la_oenb_mprj[12] vssd vccd _509_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] _205_/X vssd vccd _025_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1015 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1795_A wire1796/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2951 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1962_A wire1962/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput710 _075_/Y vssd vccd la_data_in_mprj[92] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput721 _598_/X vssd vccd la_oenb_core[101] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__024__A _024_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput732 _608_/X vssd vccd la_oenb_core[111] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput743 _618_/X vssd vccd la_oenb_core[121] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput754 wire1036/X vssd vccd la_oenb_core[16] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3675 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput765 wire1026/X vssd vccd la_oenb_core[26] vssd vccd sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] _167_/X vssd vccd _151_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xoutput776 _533_/X vssd vccd la_oenb_core[36] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput787 _543_/X vssd vccd la_oenb_core[46] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2208 wire2209/X vssd vccd wire2208/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput798 wire1002/X vssd vccd la_oenb_core[56] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1507 wire1508/X vssd vccd wire1507/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1518 wire1519/X vssd vccd _316_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2619 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1529 wire1529/A vssd vccd _585_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__397__C _397_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_751 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_180_ _180_/A _180_/B vssd vccd _180_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_3736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_294 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input261_A la_oenb_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_622 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input359_A la_oenb_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__588__B _588_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3876 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_330 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_341 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_352 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_516_ _516_/A _516_/B vssd vccd _516_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_363 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__109__A _109_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_447_ _575_/A _447_/B _447_/C vssd vccd _447_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_32_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1007_A wire1008/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_378_ _506_/A _378_/B _378_/C vssd vccd _378_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output480_A _484_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output578_A wire1077/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output745_A _620_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__385__A_N _513_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1376_A wire1376/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3743 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output912_A _123_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3787 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__498__B _498_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1543_A wire1543/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_4098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1710_A wire1710/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1808_A wire1808/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire996_A _558_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__019__A _019_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3507 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput540 wire1089/X vssd vccd la_data_in_core[54] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput551 _433_/X vssd vccd la_data_in_core[64] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3472 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput562 _443_/X vssd vccd la_data_in_core[74] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput573 _453_/X vssd vccd la_data_in_core[84] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput584 wire1072/X vssd vccd la_data_in_core[94] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2005 wire2006/X vssd vccd _572_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput595 _086_/Y vssd vccd la_data_in_mprj[103] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_21_3106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2016 wire2016/A vssd vccd _565_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2027 wire2027/A vssd vccd _525_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2038 wire2038/A vssd vccd wire2038/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1304 wire1305/X vssd vccd wire1304/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2049 wire2050/X vssd vccd _506_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1315 _270_/X vssd vccd wire1315/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1326 _251_/X vssd vccd wire1326/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1337 input95/X vssd vccd _436_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1348 wire1349/X vssd vccd _344_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1359 wire1359/A vssd vccd _367_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input107_A la_data_out_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_301_ _301_/A _301_/B vssd vccd _301_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_24_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_232_ _232_/A _232_/B vssd vccd _232_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_24_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_163_ _163_/A vssd vccd _163_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1254 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input72_A la_data_out_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_094_ _094_/A vssd vccd _094_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_13_1265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__599__A _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3640 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1860 wire1860/A vssd vccd wire1860/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1871 wire1871/A vssd vccd _625_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1882 wire1882/A vssd vccd wire1882/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1893 wire1894/X vssd vccd wire1893/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1124_A _389_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_160 _221_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_171 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_182 _358_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_193 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output862_A wire1254/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1018 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[18\] mprj_dat_i_user[18] max_length1311/X vssd vccd _132_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_28_3805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1660_A wire1660/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1758_A wire1758/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__302__A _302_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1925_A wire1926/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] _279_/X vssd vccd _099_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_28_128 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__400__A_N _400_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2460 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__A _212_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_934 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3094 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1101 _412_/X vssd vccd wire1101/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1112 _401_/X vssd vccd wire1112/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1123 _390_/X vssd vccd wire1123/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1134 _380_/X vssd vccd wire1134/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1145 _369_/X vssd vccd wire1145/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1156 wire1157/X vssd vccd wire1156/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1167 wire1168/X vssd vccd wire1167/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2141_A wire2141/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input224_A la_iena_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1178 wire1179/X vssd vccd wire1178/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1189 _358_/X vssd vccd wire1189/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_215_ _215_/A _215_/B vssd vccd _215_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_11_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_146_ _146_/A vssd vccd _146_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_1685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_077_ _077_/A vssd vccd _077_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__122__A _122_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1074_A _461_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__423__A_N _551_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3779 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output610_A _100_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1241_A wire1242/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1000 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__495__C _495_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1690 wire1691/X vssd vccd _368_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3528 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1828 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1506_A wire1507/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3252 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput109 la_data_out_mprj[7] vssd vccd _376_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2763 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2555 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_930 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_654 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_126 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2206 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_698 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__A _207_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_60 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_000_ _000_/A vssd vccd _000_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_71 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_82 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_93 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2091_A wire2092/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input174_A la_iena_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2189_A wire2190/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1279 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__446__A_N _574_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3167 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input341_A la_oenb_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input439_A mprj_dat_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input35_A la_data_out_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2262 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__596__B _596_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4120 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3739 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_6 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output560_A _441_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output658_A _028_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_129_ _129_/A vssd vccd _129_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_wire1191_A wire1192/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1289_A wire1290/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output825_A _577_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1456_A wire1456/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] _235_/X vssd vccd _055_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_2925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1623_A wire1623/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1992_A wire1993/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2846 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__A_N _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput80 la_data_out_mprj[53] vssd vccd _422_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput91 la_data_out_mprj[63] vssd vccd _432_/C vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_user_to_mprj_in_gates\[33\]_B _196_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_480_ _608_/A _480_/B _480_/C vssd vccd _480_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_26_974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1302 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3756 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input291_A la_oenb_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input389_A mprj_adr_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2506 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1087 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1838 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1415 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput440 mprj_dat_o_core[27] vssd vccd wire1364/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput451 mprj_dat_o_core[8] vssd vccd wire1347/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput462 user_irq_ena[2] vssd vccd _293_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_4215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1037_A _512_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1204_A _354_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output775_A _532_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output942_A wire1232/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput903 _116_/Y vssd vccd mprj_dat_i_core[2] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput914 wire1223/X vssd vccd mprj_dat_o_user[10] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[15\]_B _178_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput925 wire1190/X vssd vccd mprj_dat_o_user[20] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput936 wire1150/X vssd vccd mprj_dat_o_user[30] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3627 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput947 wire1284/X vssd vccd mprj_sel_o_user[2] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput958 _112_/Y vssd vccd user_irq[1] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1740_A wire1741/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_3401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1838_A wire1838/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2216 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__310__A _310_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_454 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_2487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2790 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__204__B _204_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3126 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2655 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input137_A la_iena_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_601_ _601_/A _601_/B vssd vccd _601_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_37_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_532_ _532_/A _532_/B vssd vccd _532_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input304_A la_oenb_mprj[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1586 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_463_ _591_/A _463_/B _463_/C vssd vccd _463_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_394_ _522_/A _394_/B _394_/C vssd vccd _394_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_41_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output523_A wire1105/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__130__A _130_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1154_A wire1155/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput270 la_oenb_mprj[109] vssd vccd _478_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_3579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput281 la_oenb_mprj[119] vssd vccd wire1587/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1256 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput292 la_oenb_mprj[13] vssd vccd _510_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_36_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1321_A _256_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_568 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1419_A wire1420/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] _198_/X vssd vccd _018_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1027 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1690_A wire1691/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1788_A wire1788/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__A _305_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1955_A wire1956/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput700 _066_/Y vssd vccd la_data_in_mprj[83] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput711 _076_/Y vssd vccd la_data_in_mprj[93] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput722 _599_/X vssd vccd la_oenb_core[102] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput733 _609_/X vssd vccd la_oenb_core[112] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput744 _619_/X vssd vccd la_oenb_core[122] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput755 wire1035/X vssd vccd la_oenb_core[17] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput766 _524_/X vssd vccd la_oenb_core[27] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput777 _534_/X vssd vccd la_oenb_core[37] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput788 _544_/X vssd vccd la_oenb_core[47] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput799 _554_/X vssd vccd la_oenb_core[57] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2209 wire2209/A vssd vccd wire2209/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_2734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3479 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1508 wire1508/A vssd vccd wire1508/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1519 wire1519/A vssd vccd wire1519/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_763 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3851 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3704 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3748 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__215__A _215_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1750 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3120 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2171_A wire2172/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input254_A la_iena_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_678 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input421_A mprj_dat_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3888 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_320 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_331 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_342 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_515_ _515_/A _515_/B vssd vccd _515_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_353 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_364 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_446_ _574_/A _446_/B _446_/C vssd vccd _446_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_3659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_377_ _505_/A _377_/B _377_/C vssd vccd _377_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_48_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output473_A wire1057/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output640_A _012_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output738_A _614_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3755 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1271_A wire1272/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1369_A wire1369/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3799 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3310 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1536_A wire1536/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__035__A _035_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3519 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4163 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput530 wire1099/X vssd vccd la_data_in_core[45] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput541 wire1087/X vssd vccd la_data_in_core[55] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput552 _434_/X vssd vccd la_data_in_core[65] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput563 _444_/X vssd vccd la_data_in_core[75] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput574 _454_/X vssd vccd la_data_in_core[85] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput585 wire1071/X vssd vccd la_data_in_core[95] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2006 wire2006/A vssd vccd wire2006/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput596 _087_/Y vssd vccd la_data_in_mprj[104] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2017 wire2017/A vssd vccd _564_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2028 wire2028/A vssd vccd _523_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_3287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2039 wire2039/A vssd vccd _512_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1305 _299_/X vssd vccd wire1305/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1316 _266_/X vssd vccd wire1316/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1327 _250_/X vssd vccd wire1327/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1338 input94/X vssd vccd _435_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1349 wire1349/A vssd vccd wire1349/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_39_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3924 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_858 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_300_ _300_/A _300_/B vssd vccd _300_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_42_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2017_A wire2017/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_571 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_231_ _231_/A _231_/B vssd vccd _231_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_162_ _162_/A vssd vccd _162_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3534 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input371_A la_oenb_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_093_ _093_/A vssd vccd _093_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_910 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input65_A la_data_out_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__599__B _599_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1850 wire1851/X vssd vccd _176_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1861 wire1861/A vssd vccd _169_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1872 wire1873/X vssd vccd _624_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1883 wire1884/X vssd vccd _621_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1894 wire1894/A vssd vccd wire1894/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_150 _210_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_161 _222_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_172 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_183 wire1459/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output590_A wire1136/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_194 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1117_A _396_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output688_A _055_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_429_ _557_/A _429_/B _429_/C vssd vccd _429_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1046 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output855_A wire1260/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1486_A wire1487/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4128 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1653_A wire1653/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__302__B _302_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_A mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput1 caravel_clk vssd vccd _296_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_37_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] _272_/X vssd vccd _092_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_0_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4039 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__212__B _212_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1102 _411_/X vssd vccd wire1102/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1113 _400_/X vssd vccd wire1113/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_3972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1124 _389_/X vssd vccd wire1124/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1135 _379_/X vssd vccd wire1135/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1146 wire1147/X vssd vccd wire1146/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1157 _366_/X vssd vccd wire1157/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1168 wire1169/X vssd vccd wire1168/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1179 wire1180/X vssd vccd wire1179/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_4400 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2134_A wire2134/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input217_A la_iena_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3754 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_214_ _214_/A _214_/B vssd vccd _214_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_7_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_145_ _145_/A vssd vccd _145_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[0\] mprj_dat_i_user[0] max_length1310/X vssd vccd _114_/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_32_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_076_ _076_/A vssd vccd _076_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_23_4404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1067_A _468_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output603_A _093_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1012 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1680 wire1681/X vssd vccd _373_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1691 wire1691/A vssd vccd wire1691/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1401_A wire1402/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[30\] mprj_dat_i_user[30] max_length1310/X vssd vccd _144_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_15_3264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1770_A wire1770/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1868_A wire1868/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__A _313_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__398__A_N _526_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3954 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2218 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__207__B _207_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_50 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_61 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_72 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_83 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_94 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2084_A wire2084/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input167_A la_iena_mprj[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_710 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input334_A la_oenb_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2274 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input28_A la_data_out_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4132 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_7 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_168 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_128_ _128_/A vssd vccd _128_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output553_A _435_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__133__A _133_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_059_ _059_/A vssd vccd _059_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1184_A wire1185/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output720_A _597_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output818_A _571_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3555 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1351_A wire1351/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1449_A wire1450/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] _228_/X vssd vccd _048_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1616_A wire1616/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3304 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__308__A _308_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1985_A wire1985/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire971_A wire971/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput70 la_data_out_mprj[44] vssd vccd _413_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_8_4239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput81 la_data_out_mprj[54] vssd vccd _423_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput92 la_data_out_mprj[64] vssd vccd _433_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_45_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__218__A _218_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1314 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__413__A_N _541_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input284_A la_oenb_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1011 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1055 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input451_A mprj_dat_o_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1099 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3936 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput430 mprj_dat_o_core[18] vssd vccd wire1376/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput441 mprj_dat_o_core[28] vssd vccd wire1363/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput452 mprj_dat_o_core[9] vssd vccd wire1345/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_4314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output768_A _526_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4504 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1399_A wire1400/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output935_A wire1246/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput904 _144_/Y vssd vccd mprj_dat_i_core[30] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput915 wire1220/X vssd vccd mprj_dat_o_user[11] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput926 wire1186/X vssd vccd mprj_dat_o_user[21] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput937 wire1146/X vssd vccd mprj_dat_o_user[31] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput948 wire1280/X vssd vccd mprj_sel_o_user[3] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput959 _113_/Y vssd vccd user_irq[2] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_4169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1733_A wire1734/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__310__B _310_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1062 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1900_A wire1901/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2302 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__A_N _564_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__038__A _038_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_967 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__A _501_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2667 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_600_ _600_/A _600_/B vssd vccd _600_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire2047_A wire2048/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_531_ _531_/A _531_/B vssd vccd _531_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_17_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_462_ _590_/A _462_/B _462_/C vssd vccd _462_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3808 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_393_ _521_/A _393_/B _393_/C vssd vccd _393_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_25_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input95_A la_data_out_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1707 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_820 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output516_A wire1112/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput260 la_oenb_mprj[0] vssd vccd _497_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput271 la_oenb_mprj[10] vssd vccd _507_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput282 la_oenb_mprj[11] vssd vccd _508_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput293 la_oenb_mprj[14] vssd vccd _511_/A vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_wire1147_A wire1148/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__459__A_N _587_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1314_A _277_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_3307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] _191_/X vssd vccd _011_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1039 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1683_A wire1683/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__305__B _305_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3600 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput701 _067_/Y vssd vccd la_data_in_mprj[84] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput712 _077_/Y vssd vccd la_data_in_mprj[94] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1850_A wire1851/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput723 _600_/X vssd vccd la_oenb_core[103] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1948_A wire1949/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput734 _610_/X vssd vccd la_oenb_core[113] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput745 _620_/X vssd vccd la_oenb_core[123] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput756 wire1034/X vssd vccd la_oenb_core[18] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput767 wire1025/X vssd vccd la_oenb_core[28] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput778 wire1020/X vssd vccd la_oenb_core[38] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput789 _545_/X vssd vccd la_oenb_core[48] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__321__A _321_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_powergood_check_mprj2_vdd_logic1 output954/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3160 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1509 wire1510/X vssd vccd _319_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1106 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3863 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3716 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__215__B _215_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3132 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1183 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3176 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__A _231_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input247_A la_iena_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3834 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input414_A mprj_adr_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input10_A la_data_out_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4306 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_310 _437_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_321 wire1985/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_332 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_514_ _514_/A _514_/B vssd vccd _514_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_33_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_343 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_354 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3616 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1916 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_365 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_445_ _573_/A _445_/B _445_/C vssd vccd _445_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_32_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_376_ _504_/A _376_/B _376_/C vssd vccd _376_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_2216 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output466_A wire1064/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1097_A _416_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output633_A _005_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3767 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__141__A _141_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4034 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1264_A wire1265/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3491 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output800_A wire1000/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1529_A wire1529/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4130 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1898_A wire1899/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__A _316_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4175 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput520 wire1108/X vssd vccd la_data_in_core[36] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput531 wire1098/X vssd vccd la_data_in_core[46] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput542 wire1085/X vssd vccd la_data_in_core[56] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput553 _435_/X vssd vccd la_data_in_core[66] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput564 _445_/X vssd vccd la_data_in_core[76] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput575 _455_/X vssd vccd la_data_in_core[86] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__051__A _051_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput586 wire1070/X vssd vccd la_data_in_core[96] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2007 wire2008/X vssd vccd _571_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput597 _088_/Y vssd vccd la_data_in_mprj[105] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2018 wire2018/A vssd vccd _563_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2029 wire2029/A vssd vccd _521_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1306 _298_/X vssd vccd wire1306/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input2_A caravel_clk2 vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1317 _262_/X vssd vccd wire1317/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1328 _249_/X vssd vccd wire1328/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_41_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1339 input93/X vssd vccd _434_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_230_ _230_/A _230_/B vssd vccd _230_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_23_583 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__226__A _226_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_161_ _161_/A vssd vccd _161_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input197_A la_iena_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3568 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_092_ _092_/A vssd vccd _092_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input364_A la_oenb_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input58_A la_data_out_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_966 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_454 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1571 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1840 wire1840/A vssd vccd _184_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1851 wire1851/A vssd vccd wire1851/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1862 wire1862/A vssd vccd _168_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1873 wire1874/X vssd vccd wire1873/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1884 wire1885/X vssd vccd wire1884/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1895 wire1896/X vssd vccd _617_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_140 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_151 _210_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_162 _222_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_173 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_184 wire1461/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_195 _524_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_428_ _556_/A _428_/B _428_/C vssd vccd _428_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_18_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output583_A wire1073/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__136__A _136_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_359_ _359_/A _359_/B vssd vccd _359_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output750_A wire1040/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1381_A wire1382/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1479_A wire1480/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3531 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] wire1319/X vssd vccd wire962/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_44_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1646_A wire1647/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[0\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput2 caravel_clk2 vssd vccd _297_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_2509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__046__A _046_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4007 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1103 _410_/X vssd vccd wire1103/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1114 _399_/X vssd vccd wire1114/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1125 _388_/X vssd vccd wire1125/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1136 _378_/X vssd vccd wire1136/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1147 wire1148/X vssd vccd wire1147/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1158 wire1159/X vssd vccd wire1158/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_0_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1169 _363_/X vssd vccd wire1169/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4412 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input112_A la_data_out_mprj[82] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_196 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_213_ _213_/A _213_/B vssd vccd _213_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_3332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_144_ _144_/A vssd vccd _144_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_075_ _075_/A vssd vccd _075_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__B _403_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3895 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3472 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1670 wire1671/X vssd vccd _377_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1681 wire1681/A vssd vccd wire1681/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1692 wire1693/X vssd vccd _367_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1227_A wire1228/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output798_A wire1002/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] _173_/X vssd vccd _157_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xuser_wb_dat_gates\[23\] mprj_dat_i_user[23] max_length1310/X vssd vccd _137_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1596_A _479_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1763_A wire1764/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__313__B _313_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1930_A wire1930/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3247 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] _284_/X vssd vccd _104_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_29_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_40 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_51 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_62 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_73 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_84 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_95 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__504__A _504_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_46_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2077_A wire2078/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input327_A la_oenb_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_954 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__492__A_N _620_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_8 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1126 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_49_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_127_ _127_/A vssd vccd _127_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_058_ _058_/A vssd vccd _058_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output546_A wire1140/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output713_A _078_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1344_A wire1345/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2190 wire2190/A vssd vccd wire2190/X vssd vccd sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] _221_/X vssd vccd _041_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_19_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1511_A wire1511/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3316 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__308__B _308_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1880_A wire1881/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2372 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1978_A wire1978/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3972 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire964_A wire964/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2247 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__324__A _324_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
Xinput60 la_data_out_mprj[35] vssd vccd _404_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1546 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput71 la_data_out_mprj[45] vssd vccd _414_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput82 la_data_out_mprj[55] vssd vccd _424_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput93 la_data_out_mprj[65] vssd vccd input93/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_4431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1326 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__234__A _234_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2194_A wire2194/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input277_A la_oenb_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1067 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4555 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input444_A mprj_dat_o_core[30] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3843 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input40_A la_data_out_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput420 mprj_cyc_o_core vssd vccd wire1397/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput431 mprj_dat_o_core[19] vssd vccd wire1375/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput442 mprj_dat_o_core[29] vssd vccd wire1362/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__400__C _400_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput453 mprj_iena_wb vssd vccd _294_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1502 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output496_A wire1130/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1579 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4516 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__144__A _144_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__388__A_N _516_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1294_A wire1295/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput905 _145_/Y vssd vccd mprj_dat_i_core[31] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput916 wire1217/X vssd vccd mprj_dat_o_user[12] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output830_A _582_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput927 wire1182/X vssd vccd mprj_dat_o_user[22] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput938 wire1244/X vssd vccd mprj_dat_o_user[3] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output928_A wire1178/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput949 wire1303/X vssd vccd mprj_stb_o_user vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1461_A wire1461/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1559_A _417_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1726_A wire1727/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__054__A _054_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__501__B _501_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2679 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_530_ _530_/A _530_/B vssd vccd _530_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__229__A _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_461_ _589_/A _461_/B _461_/C vssd vccd _461_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_392_ _520_/A _392_/B _392_/C vssd vccd _392_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_17_3680 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2207_A wire2208/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input394_A mprj_adr_o_core[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input88_A la_data_out_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__411__B _411_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3892 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput250 la_iena_mprj[91] vssd vccd _254_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput261 la_oenb_mprj[100] vssd vccd wire1607/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput272 la_oenb_mprj[110] vssd vccd _479_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput283 la_oenb_mprj[120] vssd vccd wire1586/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_23_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output509_A wire1118/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput294 la_oenb_mprj[15] vssd vccd _512_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_53_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1042_A wire1043/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_4047 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__139__A _139_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output780_A wire1050/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1307_A wire1308/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output878_A wire1276/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2342 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1676_A wire1677/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput702 _068_/Y vssd vccd la_data_in_mprj[85] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput713 _078_/Y vssd vccd la_data_in_mprj[95] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput724 _601_/X vssd vccd la_oenb_core[104] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput735 _611_/X vssd vccd la_oenb_core[114] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__602__A _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput746 _621_/X vssd vccd la_oenb_core[124] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput757 wire1033/X vssd vccd la_oenb_core[19] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1843_A wire1843/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput768 _526_/X vssd vccd la_oenb_core[29] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput779 wire1019/X vssd vccd la_oenb_core[39] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__321__B _321_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_4496 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__A_N _531_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__049__A _049_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__512__A _512_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4503 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__231__B _231_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3846 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input142_A la_iena_mprj[109] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2157_A wire2158/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input407_A mprj_adr_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_300 wire1907/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_311 _341_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_322 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_513_ _513_/A _513_/B vssd vccd _513_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_333 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_344 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_355 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_366 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_444_ _572_/A _444_/B _444_/C vssd vccd _444_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_375_ _503_/A _375_/B _375_/C vssd vccd _375_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__406__B _406_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2651 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__426__A_N _554_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1257_A _324_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1424_A wire1425/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] _203_/X vssd vccd _023_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_24_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1793_A wire1794/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__316__B _316_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_1774 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1960_A wire1961/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[90\]_B wire1324/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput510 wire1117/X vssd vccd la_data_in_core[27] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__332__A _332_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput521 wire1107/X vssd vccd la_data_in_core[37] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_4187 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput532 wire1097/X vssd vccd la_data_in_core[47] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput543 wire1084/X vssd vccd la_data_in_core[57] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput554 _436_/X vssd vccd la_data_in_core[67] vssd vccd sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] _165_/X vssd vccd _149_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xoutput565 _446_/X vssd vccd la_data_in_core[77] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput576 _456_/X vssd vccd la_data_in_core[87] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput587 wire1069/X vssd vccd la_data_in_core[97] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2008 wire2008/A vssd vccd wire2008/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput598 _089_/Y vssd vccd la_data_in_mprj[106] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2019 wire2019/A vssd vccd _562_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_3278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1307 wire1308/X vssd vccd wire1307/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1318 _259_/X vssd vccd wire1318/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1329 _248_/X vssd vccd wire1329/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__507__A _507_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3650 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_595 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_160_ _160_/A vssd vccd _160_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__226__B _226_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_091_ _091_/A vssd vccd _091_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_B _244_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__449__A_N _577_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__242__A _242_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input357_A la_oenb_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1830 wire1830/A vssd vccd _190_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1841 wire1841/A vssd vccd _183_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1852 wire1853/X vssd vccd _175_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1863 wire1864/X vssd vccd _167_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1874 wire1875/X vssd vccd wire1874/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1885 wire1885/A vssd vccd wire1885/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1896 wire1897/X vssd vccd wire1896/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_130 _527_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_141 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4148 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_152 _212_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_163 _228_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3594 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_174 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_185 _559_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_196 _618_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_427_ _555_/A _427_/B _427_/C vssd vccd _427_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_42_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_358_ _358_/A _358_/B vssd vccd _358_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_50_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1005_A wire1006/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output576_A _456_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_289_ _289_/A _289_/B vssd vccd _289_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[72\]_B _235_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output743_A _618_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1374_A wire1374/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] wire1326/X vssd vccd wire969/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_26_3587 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1541_A wire1541/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1639_A wire1640/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput3 caravel_rstn vssd vccd input3/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire994_A _587_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__327__A _327_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_510 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4019 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__062__A _062_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2639 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3272 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1104 _409_/X vssd vccd wire1104/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1115 _398_/X vssd vccd wire1115/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1126 _387_/X vssd vccd wire1126/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1137 _377_/X vssd vccd wire1137/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1148 wire1149/X vssd vccd wire1148/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1159 wire1160/X vssd vccd wire1159/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input105_A la_data_out_mprj[76] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2022_A wire2022/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__237__A _237_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_690 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_212_ _212_/A _212_/B vssd vccd _212_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_3300 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_143_ _143_/A vssd vccd _143_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_52_1081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3388 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input70_A la_data_out_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_074_ _074_/A vssd vccd _074_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__403__C _403_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_230 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1391 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1660 wire1660/A vssd vccd wire1660/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1671 wire1671/A vssd vccd wire1671/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2844 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1682 wire1683/X vssd vccd _372_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1693 wire1693/A vssd vccd wire1693/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1122_A _391_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output860_A wire1256/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[16\] mprj_dat_i_user[16] max_length1311/X vssd vccd _130_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_31_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1491_A wire1492/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire990 wire990/A vssd vccd _091_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1756_A wire1756/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3204 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__610__A _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_2503 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1923_A wire1924/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3259 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] wire1314/X vssd vccd wire985/A
+ vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_39_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_602 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__057__A _057_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_30 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_41 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_52 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_63 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_74 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_85 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_B _199_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_96 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__504__B _504_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[120\]_B _283_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__520__A _520_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input222_A la_iena_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_9 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3174 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_126_ _126_/A vssd vccd _126_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__414__B _414_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[111\]_B _274_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_057_ _057_/A vssd vccd _057_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_3721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4236 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3671 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output539_A wire1090/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1072_A _463_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_4190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2180 wire2181/X vssd vccd _444_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2191 wire2191/A vssd vccd _438_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1337_A input95/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3386 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1490 wire1491/X vssd vccd _324_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3328 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1504_A wire1504/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[20\]_A mprj_dat_i_user[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__605__A _605_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3984 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1873_A wire1874/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__324__B _324_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[102\]_B _265_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3402 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput50 la_data_out_mprj[26] vssd vccd _395_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput61 la_data_out_mprj[36] vssd vccd _405_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput72 la_data_out_mprj[46] vssd vccd _415_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput83 la_data_out_mprj[56] vssd vccd _425_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_28_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput94 la_data_out_mprj[66] vssd vccd input94/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3242 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[11\]_A mprj_dat_i_user[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3895 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__515__A _515_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__234__B _234_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input172_A la_iena_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__250__A _250_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3855 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2266 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input437_A mprj_dat_o_core[24] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput410 mprj_adr_o_core[2] vssd vccd wire1441/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput421 mprj_dat_o_core[0] vssd vccd wire1393/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_3899 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input33_A la_data_out_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput432 mprj_dat_o_core[1] vssd vccd wire1374/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput443 mprj_dat_o_core[2] vssd vccd wire1361/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput454 mprj_sel_o_core[0] vssd vccd _301_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1383 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__409__B _409_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1514 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output489_A _492_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_4456 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output656_A _026_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_109_ _109_/A vssd vccd _109_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
Xoutput906 _117_/Y vssd vccd mprj_dat_i_core[3] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput917 wire1214/X vssd vccd mprj_dat_o_user[13] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput928 wire1178/X vssd vccd mprj_dat_o_user[23] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_7_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4000 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1287_A wire1288/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput939 wire1241/X vssd vccd mprj_dat_o_user[4] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output823_A _576_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1454_A wire1455/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] _233_/X vssd vccd _053_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XANTENNA_wire1621_A wire1621/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__319__B _319_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1990_A wire1991/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2760 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__335__A _335_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__A_N _610_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__070__A _070_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_460_ _588_/A _460_/B _460_/C vssd vccd _460_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__229__B _229_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_4360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_391_ _519_/A _391_/B _391_/C vssd vccd _391_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_53_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2102_A wire2103/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__A _245_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input387_A la_oenb_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3860 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4386 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_4160 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput240 la_iena_mprj[82] vssd vccd _245_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput251 la_iena_mprj[92] vssd vccd _255_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput262 la_oenb_mprj[101] vssd vccd wire1606/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput273 la_oenb_mprj[111] vssd vccd wire1595/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput284 la_oenb_mprj[121] vssd vccd wire1585/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput295 la_oenb_mprj[16] vssd vccd _513_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_18_3412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1035_A _514_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_589_ _589_/A _589_/B vssd vccd _589_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_18_3489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_766 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1202_A wire1203/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output773_A wire1024/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__155__A _155_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2354 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output940_A wire1238/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2387 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4336 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput703 _069_/Y vssd vccd la_data_in_mprj[86] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1571_A _400_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput714 _079_/Y vssd vccd la_data_in_mprj[96] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1669_A wire1669/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput725 _602_/X vssd vccd la_oenb_core[105] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput736 _612_/X vssd vccd la_oenb_core[115] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__602__B _602_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput747 _622_/X vssd vccd la_oenb_core[125] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput758 wire1052/X vssd vccd la_oenb_core[1] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput769 wire1051/X vssd vccd la_oenb_core[2] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1836_A wire1836/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__065__A _065_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__512__B _512_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_2411 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2455 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3814 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3983 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2052_A wire2052/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input135_A la_iena_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_4411 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__378__A_N _506_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_301 wire1951/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_512_ _512_/A _512_/B vssd vccd _512_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_312 _351_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_323 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input302_A la_oenb_mprj[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_334 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_345 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_356 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_443_ _571_/A _443_/B _443_/C vssd vccd _443_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4032 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_374_ _502_/A _374_/B _374_/C vssd vccd _374_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3808 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output521_A wire1107/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1152_A wire1153/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2623 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_814 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1417_A wire1418/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] _196_/X vssd vccd _016_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_51_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__613__A _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1953_A wire1954/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput500 wire1126/X vssd vccd la_data_in_core[18] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput511 wire1116/X vssd vccd la_data_in_core[28] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput522 wire1106/X vssd vccd la_data_in_core[38] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__332__B _332_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput533 wire1096/X vssd vccd la_data_in_core[48] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput544 wire1082/X vssd vccd la_data_in_core[58] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput555 _437_/X vssd vccd la_data_in_core[68] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput566 _447_/X vssd vccd la_data_in_core[78] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_A mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput577 _457_/X vssd vccd la_data_in_core[88] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput588 wire1068/X vssd vccd la_data_in_core[98] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2009 wire2009/A vssd vccd _570_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput599 _090_/Y vssd vccd la_data_in_mprj[107] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1308 wire1309/X vssd vccd wire1308/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1319 _258_/X vssd vccd wire1319/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__507__B _507_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_090_ _090_/A vssd vccd _090_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_30_2240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__523__A _523_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input252_A la_iena_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1820 wire1820/A vssd vccd _206_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1831 wire1832/X vssd vccd _189_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1842 wire1842/A vssd vccd _329_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1853 wire1853/A vssd vccd wire1853/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1864 wire1864/A vssd vccd wire1864/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_836 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1875 wire1875/A vssd vccd wire1875/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1886 wire1887/X vssd vccd _620_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1897 wire1897/A vssd vccd wire1897/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_120 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_131 _527_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_142 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_153 _212_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_164 _228_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_175 _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_186 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_426_ _554_/A _426_/B _426_/C vssd vccd _426_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__417__B _417_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_197 _303_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_357_ _357_/A _357_/B vssd vccd _357_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_32_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_288_ _288_/A _288_/B vssd vccd _288_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output471_A wire1059/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output569_A _449_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_740 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output736_A _612_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1367_A wire1367/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3599 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1534_A wire1534/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput4 la_data_out_mprj[0] vssd vccd _369_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_20_3176 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1701_A wire1701/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__608__A _608_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__327__B _327_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_2360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire987_A wire987/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__343__A _343_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2607 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1105 _408_/X vssd vccd wire1105/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1116 _397_/X vssd vccd wire1116/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1127 _386_/X vssd vccd wire1127/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1138 _376_/X vssd vccd wire1138/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1149 _368_/X vssd vccd wire1149/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__518__A _518_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__237__B _237_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2015_A wire2015/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__416__A_N _416_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_211_ _211_/A _211_/B vssd vccd _211_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_142_ _142_/A vssd vccd _142_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__A _253_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_073_ _073_/A vssd vccd _073_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_2655 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input63_A la_data_out_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4131 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_286 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_600 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1650 wire1651/X vssd vccd _386_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1661 wire1662/X vssd vccd _381_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1672 wire1673/X vssd vccd _376_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1683 wire1683/A vssd vccd wire1683/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1694 wire1695/X vssd vccd _366_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4071 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1115_A _398_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output686_A _053_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_409_ _409_/A_N _409_/B _409_/C vssd vccd _409_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_50_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output853_A wire1262/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__163__A _163_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1484_A wire1484/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire980 wire980/A vssd vccd _109_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_31_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire991 wire991/A vssd vccd _090_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1749_A wire1750/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__610__B _610_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1916_A wire1917/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] wire1315/X vssd vccd wire991/A
+ vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA__439__A_N _567_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__A _338_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1011 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_20 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_31 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_42 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_53 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_64 mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_75 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__073__A _073_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_86 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_97 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2415 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__520__B _520_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3750 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input215_A la_iena_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2132_A wire2132/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__248__A _248_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_125_ _125_/A vssd vccd _125_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__414__C _414_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3186 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_056_ _056_/A vssd vccd _056_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__430__B _430_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3490 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1065_A _470_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2170 wire2170/A vssd vccd wire2170/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2181 wire2181/A vssd vccd wire2181/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2192 wire2192/A vssd vccd _437_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1480 wire1481/X vssd vccd wire1480/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1491 wire1492/X vssd vccd wire1491/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1232_A wire1233/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[20\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2639 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1699_A wire1699/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__605__B _605_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput40 la_data_out_mprj[17] vssd vccd _386_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1866_A wire1866/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput51 la_data_out_mprj[27] vssd vccd _396_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4159 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput62 la_data_out_mprj[37] vssd vccd _406_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput73 la_data_out_mprj[47] vssd vccd _416_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_3436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput84 la_data_out_mprj[57] vssd vccd _426_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_890 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput95 la_data_out_mprj[67] vssd vccd input95/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__621__A _621_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__340__B _340_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_912 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__068__A _068_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[11\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__515__B _515_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__531__A _531_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input165_A la_iena_mprj[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2082_A wire2083/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2278 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput400 mprj_adr_o_core[20] vssd vccd wire1484/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput411 mprj_adr_o_core[30] vssd vccd wire1436/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput422 mprj_dat_o_core[10] vssd vccd wire1390/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input332_A la_oenb_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput433 mprj_dat_o_core[20] vssd vccd wire1371/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput444 mprj_dat_o_core[30] vssd vccd wire1359/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput455 mprj_sel_o_core[1] vssd vccd _302_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input26_A la_data_out_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__409__C _409_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3362 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1526 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__425__B _425_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_108_ _108_/A vssd vccd _108_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_29_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput907 _118_/Y vssd vccd mprj_dat_i_core[4] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_49_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output551_A _433_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput918 wire1211/X vssd vccd mprj_dat_o_user[14] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput929 wire1174/X vssd vccd mprj_dat_o_user[24] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output649_A _020_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_4012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_039_ _039_/A vssd vccd _039_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_wire1182_A wire1183/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output816_A _569_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1447_A wire1448/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] _226_/X vssd vccd _046_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_36_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3159 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__616__A _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1983_A wire1983/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__335__B _335_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4028 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1356 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__351__A _351_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_318 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_390_ _518_/A _390_/B _390_/C vssd vccd _390_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_0_1270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__526__A _526_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__245__B _245_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3871 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input282_A la_oenb_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2318 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__A _261_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4354 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3631 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3872 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3675 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput230 la_iena_mprj[73] vssd vccd _236_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput241 la_iena_mprj[83] vssd vccd _246_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput252 la_iena_mprj[93] vssd vccd _256_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput263 la_oenb_mprj[102] vssd vccd wire1605/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput274 la_oenb_mprj[112] vssd vccd wire1594/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_49_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput285 la_oenb_mprj[122] vssd vccd wire1584/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput296 la_oenb_mprj[17] vssd vccd _514_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_35_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_712 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_588_ _588_/A _588_/B vssd vccd _588_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_34_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_970 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3094 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output766_A _524_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1397_A wire1397/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4107 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4348 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1080 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output933_A wire1158/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput704 _070_/Y vssd vccd la_data_in_mprj[87] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput715 _080_/Y vssd vccd la_data_in_mprj[97] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__171__A _171_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput726 _603_/X vssd vccd la_oenb_core[106] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3406 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput737 _613_/X vssd vccd la_oenb_core[116] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1564_A _412_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3428 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput748 _623_/X vssd vccd la_oenb_core[126] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_7_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput759 wire1032/X vssd vccd la_oenb_core[20] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2006 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1731_A wire1731/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1829_A wire1829/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__346__A _346_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1407 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__081__A _081_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_616 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3951 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2467 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3995 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2191 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_506 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input128_A la_data_out_mprj[97] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2045_A wire2046/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_302 wire1954/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_511_ _511_/A _511_/B vssd vccd _511_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_313 wire1885/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_324 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_335 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_346 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4000 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_357 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_442_ _570_/A _442_/B _442_/C vssd vccd _442_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_19_3788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__256__A _256_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4044 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_373_ _501_/A _373_/B _373_/C vssd vccd _373_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input93_A la_data_out_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[9\] mprj_dat_i_user[9] _294_/X vssd vccd _123_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_26_3715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__422__C _422_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4004 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3680 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output514_A wire1114/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2635 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1145_A _369_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3232 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1312_A _287_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3276 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__A_N _472_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__166__A _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] _189_/X vssd vccd _009_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_14_2417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1681_A wire1681/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1779_A wire1779/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__613__B _613_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput501 wire1125/X vssd vccd la_data_in_core[19] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput512 wire1115/X vssd vccd la_data_in_core[29] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput523 wire1105/X vssd vccd la_data_in_core[39] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput534 wire1095/X vssd vccd la_data_in_core[49] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1946_A wire1947/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput545 wire1081/X vssd vccd la_data_in_core[59] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput556 _438_/X vssd vccd la_data_in_core[69] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_wb_dat_gates\[3\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput567 _448_/X vssd vccd la_data_in_core[79] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput578 wire1077/X vssd vccd la_data_in_core[89] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput589 wire1067/X vssd vccd la_data_in_core[99] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_3_3021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1309 _296_/X vssd vccd wire1309/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3892 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_358 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__076__A _076_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2252 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__523__B _523_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2231 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2162_A wire2163/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_2275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input245_A la_iena_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1810 wire1810/A vssd vccd _233_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1821 wire1821/A vssd vccd _205_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1832 wire1832/A vssd vccd wire1832/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1843 wire1843/A vssd vccd _182_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1854 wire1855/X vssd vccd _174_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1865 wire1866/X vssd vccd _166_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input412_A mprj_adr_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1876 wire1877/X vssd vccd _623_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1887 wire1888/X vssd vccd wire1887/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__495__A_N _623_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1898 wire1899/X vssd vccd _616_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_110 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_121 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_132 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_143 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_154 _213_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_165 _228_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_176 _342_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_187 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_425_ _553_/A _425_/B _425_/C vssd vccd _425_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_35_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_198 _303_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__417__C _417_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_356_ _356_/A _356_/B vssd vccd _356_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_31_2027 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_287_ _287_/A _287_/B vssd vccd _287_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_31_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__433__B _433_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output464_A wire1066/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1095_A _418_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output729_A _606_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1262_A wire1263/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput5 la_data_out_mprj[100] vssd vccd _469_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_42_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3188 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__B _608_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1896_A wire1897/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__624__A _624_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__343__B _343_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2619 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_906 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1106 _407_/X vssd vccd wire1106/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1117 _396_/X vssd vccd wire1117/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1128 _385_/X vssd vccd wire1128/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1139 _375_/X vssd vccd wire1139/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4426 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__518__B _518_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_210_ _210_/A _210_/B vssd vccd _210_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_51_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__534__A _534_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
X_141_ _141_/A vssd vccd _141_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_49_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input195_A la_iena_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__253__B _253_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_072_ _072_/A vssd vccd _072_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_2645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2667 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4555 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input362_A la_oenb_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input56_A la_data_out_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1640 wire1640/A vssd vccd wire1640/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1651 wire1651/A vssd vccd wire1651/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1662 wire1662/A vssd vccd wire1662/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1673 wire1673/A vssd vccd wire1673/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1684 wire1685/X vssd vccd _371_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1695 wire1695/A vssd vccd wire1695/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__428__B _428_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_372 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_408_ _536_/A _408_/B _408_/C vssd vccd _408_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output581_A wire1075/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1108_A _405_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_32_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_339_ _339_/A _339_/B vssd vccd _339_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_35_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire970 wire970/A vssd vccd _070_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_output846_A wire1044/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire981 wire981/A vssd vccd _106_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire992 wire992/A vssd vccd _086_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1477_A wire1478/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] wire1321/X vssd vccd wire964/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_6_4159 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3364 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1644_A wire1644/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1811_A wire1811/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_2312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1909_A wire1910/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__619__A _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__338__B _338_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1023 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_692 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_10 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_21 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_32 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__354__A _354_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_43 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_54 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_65 mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_76 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_87 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_98 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2427 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4463 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3762 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__529__A _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__248__B _248_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input110_A la_data_out_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2125_A wire2125/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input208_A la_iena_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1243 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__264__A _264_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_124_ _124_/A vssd vccd _124_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_32_2188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3198 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_055_ _055_/A vssd vccd _055_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__430__C _430_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1550 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2160 wire2161/X vssd vccd wire2160/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2171 wire2172/X vssd vccd _448_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2182 wire2183/X vssd vccd _443_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2193 wire2193/A vssd vccd _436_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1058_A _477_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_2560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1470 wire1471/X vssd vccd wire1470/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1481 wire1481/A vssd vccd wire1481/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1492 wire1493/X vssd vccd wire1492/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1225_A _347_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output796_A _551_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__174__A _174_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2807 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[21\] mprj_dat_i_user[21] max_length1310/X vssd vccd _135_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput30 la_data_out_mprj[123] vssd vccd _492_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_50_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput41 la_data_out_mprj[18] vssd vccd _387_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput52 la_data_out_mprj[28] vssd vccd _397_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput63 la_data_out_mprj[38] vssd vccd _407_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput74 la_data_out_mprj[48] vssd vccd _417_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1761_A wire1762/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput85 la_data_out_mprj[58] vssd vccd input85/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput96 la_data_out_mprj[68] vssd vccd input96/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1859_A wire1860/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__621__B _621_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2769 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__406__A_N _406_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__349__A _349_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3875 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__531__B _531_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2075_A wire2075/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input158_A la_iena_mprj[123] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_4332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput401 mprj_adr_o_core[21] vssd vccd wire1481/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput412 mprj_adr_o_core[31] vssd vccd wire1431/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput423 mprj_dat_o_core[11] vssd vccd wire1388/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput434 mprj_dat_o_core[21] vssd vccd wire1370/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput445 mprj_dat_o_core[31] vssd vccd wire1358/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput456 mprj_sel_o_core[2] vssd vccd _303_/B vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input325_A la_oenb_mprj[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__259__A _259_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input19_A la_data_out_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_2651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__425__C _425_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_107_ _107_/A vssd vccd _107_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput908 _119_/Y vssd vccd mprj_dat_i_core[5] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput919 wire1208/X vssd vccd mprj_dat_o_user[15] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__429__A_N _557_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_038_ _038_/A vssd vccd _038_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__441__B _441_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output544_A wire1082/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1175_A wire1176/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output809_A _563_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1342_A wire1343/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__169__A _169_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] _219_/X vssd vccd _039_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_35_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__616__B _616_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1976_A wire1976/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__351__B _351_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3030 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__079__A _079_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_776 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3514 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__526__B _526_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__A _542_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2192_A wire2192/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input275_A la_oenb_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__261__B _261_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input442_A mprj_dat_o_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3518 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3687 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput220 la_iena_mprj[64] vssd vccd _227_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput231 la_iena_mprj[74] vssd vccd _237_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_0_374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput242 la_iena_mprj[84] vssd vccd _247_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput253 la_iena_mprj[94] vssd vccd _257_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput264 la_oenb_mprj[103] vssd vccd _472_/A_N vssd vccd sky130_fd_sc_hd__buf_6
Xinput275 la_oenb_mprj[113] vssd vccd wire1593/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput286 la_oenb_mprj[123] vssd vccd wire1583/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput297 la_oenb_mprj[18] vssd vccd _515_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_587_ _587_/A _587_/B vssd vccd _587_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__436__B _436_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output494_A wire1132/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_779 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_982 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output661_A _031_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output759_A wire1032/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1292_A wire1293/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4119 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput705 _071_/Y vssd vccd la_data_in_mprj[88] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput716 _081_/Y vssd vccd la_data_in_mprj[98] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput727 _604_/X vssd vccd la_oenb_core[107] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput738 _614_/X vssd vccd la_oenb_core[117] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput749 _624_/X vssd vccd la_oenb_core[127] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output926_A wire1186/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2430 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1724_A wire1725/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_890 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__346__B _346_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[93\]_B wire1321/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__362__A _362_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1799 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3963 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_518 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_510_ _510_/A _510_/B vssd vccd _510_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_303 wire1956/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_314 wire2109/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_325 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_336 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__537__A _537_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_347 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3767 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_441_ _569_/A _441_/B _441_/C vssd vccd _441_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_52_4061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_358 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4012 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__256__B _256_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_372_ _500_/A _372_/B _372_/C vssd vccd _372_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_4056 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2205_A wire2206/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input392_A mprj_adr_o_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[84\]_B wire1330/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2692 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input86_A la_data_out_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__272__A _272_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4428 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3692 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3462 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_827 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output507_A wire1120/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1040_A _509_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1138_A _376_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3244 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1305_A _299_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output876_A wire1278/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] _182_/X vssd vccd _002_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[75\]_B _238_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__182__A _182_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1674_A wire1675/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_4157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput502 wire1144/X vssd vccd la_data_in_core[1] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput513 wire1143/X vssd vccd la_data_in_core[2] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput524 wire1142/X vssd vccd la_data_in_core[3] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput535 wire1141/X vssd vccd la_data_in_core[4] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput546 wire1140/X vssd vccd la_data_in_core[5] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2650 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput557 wire1139/X vssd vccd la_data_in_core[6] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1841_A wire1841/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput568 wire1138/X vssd vccd la_data_in_core[7] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1939_A wire1940/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3259 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput579 wire1137/X vssd vccd la_data_in_core[8] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3860 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_3998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__357__A _357_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1964 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1243 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__092__A _092_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2243 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3771 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1800 wire1800/A vssd vccd _256_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input140_A la_iena_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1811 wire1811/A vssd vccd _298_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2155_A wire2155/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1822 wire1822/A vssd vccd _204_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input238_A la_iena_mprj[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1833 wire1834/X vssd vccd _188_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1844 wire1844/A vssd vccd _181_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1855 wire1855/A vssd vccd wire1855/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1866 wire1866/A vssd vccd wire1866/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1877 wire1878/X vssd vccd wire1877/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1888 wire1888/A vssd vccd wire1888/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1899 wire1900/X vssd vccd wire1899/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input405_A mprj_adr_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_100 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_111 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__267__A _267_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_122 mprj_dat_i_user[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_133 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_144 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1706 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_155 _219_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_166 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_424_ _552_/A _424_/B _424_/C vssd vccd _424_/X vssd vccd sky130_fd_sc_hd__and3b_1
XFILLER_37_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_177 _380_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_188 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_199 _303_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_355_ _355_/A _355_/B vssd vccd _355_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_50_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_286_ _286_/A _286_/B vssd vccd _286_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_2451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__433__C _433_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4203 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1339 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1255_A _327_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2674 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput6 la_data_out_mprj[101] vssd vccd _470_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1422_A wire1423/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__177__A _177_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1791_A wire1792/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1889_A wire1890/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__624__B _624_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_568 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] _625_/X vssd vccd _147_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_40_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1107 _406_/X vssd vccd wire1107/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1118 _395_/X vssd vccd wire1118/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1129 _384_/X vssd vccd wire1129/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__087__A _087_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4438 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_660 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[39\]_B _202_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_140_ _140_/A vssd vccd _140_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_user_to_mprj_in_gates\[123\]_B wire1313/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_071_ _071_/A vssd vccd _071_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4523 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input188_A la_iena_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1360 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2679 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4567 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__550__A _550_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input355_A la_oenb_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4100 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_767 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__462__A_N _590_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input49_A la_data_out_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1630 wire1630/A vssd vccd _443_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1641 wire1642/X vssd vccd _391_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1652 wire1653/X vssd vccd _385_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1663 wire1664/X vssd vccd _380_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1674 wire1675/X vssd vccd _375_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4040 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1685 wire1685/A vssd vccd wire1685/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1696 wire1697/X vssd vccd _365_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__428__C _428_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_407_ _535_/A _407_/B _407_/C vssd vccd _407_/X vssd vccd sky130_fd_sc_hd__and3b_4
XPHY_90 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_384 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__444__B _444_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[114\]_B wire1314/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_338_ _338_/A _338_/B vssd vccd _338_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output574_A _454_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_269_ _269_/A _269_/B vssd vccd _269_/X vssd vccd sky130_fd_sc_hd__and2_4
Xwire971 wire971/A vssd vccd _069_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_31_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_4011 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire982 wire982/A vssd vccd _105_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire993 wire993/A vssd vccd _083_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_output741_A wire1041/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output839_A _590_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1372_A wire1373/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3376 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] wire1328/X vssd vccd wire971/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_39_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1637_A wire1638/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__619__B _619_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[23\]_A mprj_dat_i_user[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_11 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_22 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_B _268_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__354__B _354_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_33 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_44 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_55 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_66 mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_77 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_88 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_99 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__485__A_N _613_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2382 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_A mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2020_A wire2020/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input103_A la_data_out_mprj[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2118_A wire2118/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__545__A _545_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__264__B _264_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_123_ _123_/A vssd vccd _123_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_054_ _054_/A vssd vccd _054_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__280__A _280_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire2150 wire2151/X vssd vccd wire2150/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_4068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2161 wire2161/A vssd vccd wire2161/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2172 wire2172/A vssd vccd wire2172/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2183 wire2183/A vssd vccd wire2183/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2194 wire2194/A vssd vccd _435_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1460 wire1461/X vssd vccd wire1460/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1471 wire1471/A vssd vccd wire1471/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__439__B _439_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1482 wire1483/X vssd vccd _325_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2583 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1493 wire1493/A vssd vccd wire1493/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1120_A _393_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1218_A wire1219/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output691_A _058_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output789_A _545_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[14\] mprj_dat_i_user[14] _294_/X vssd vccd _128_/A vssd vccd sky130_fd_sc_hd__nand2_2
Xinput20 la_data_out_mprj[114] vssd vccd _483_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_28_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput31 la_data_out_mprj[124] vssd vccd input31/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_50_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput42 la_data_out_mprj[19] vssd vccd _388_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_out_mprj[29] vssd vccd _398_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput64 la_data_out_mprj[39] vssd vccd _408_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput75 la_data_out_mprj[49] vssd vccd _418_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput86 la_data_out_mprj[59] vssd vccd _428_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__A _190_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput97 la_data_out_mprj[69] vssd vccd input97/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1921_A wire1921/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] _275_/X vssd vccd wire987/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XANTENNA__349__B _349_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4408 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__365__A _365_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput402 mprj_adr_o_core[22] vssd vccd wire1476/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput413 mprj_adr_o_core[3] vssd vccd wire1426/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_2190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput424 mprj_dat_o_core[12] vssd vccd wire1386/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_3790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2068_A wire2068/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput435 mprj_dat_o_core[22] vssd vccd wire1369/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput446 mprj_dat_o_core[3] vssd vccd wire1357/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput457 mprj_sel_o_core[3] vssd vccd _304_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_22_3582 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input220_A la_iena_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input318_A la_oenb_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__A _275_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2554 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2674 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_106_ _106_/A vssd vccd _106_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput909 _120_/Y vssd vccd mprj_dat_i_core[6] vssd vccd sky130_fd_sc_hd__buf_8
X_037_ _037_/A vssd vccd _037_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__441__C _441_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4036 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output537_A wire1092/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1070_A _465_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1168_A wire1169/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1056 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1290 wire1291/X vssd vccd wire1290/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_39_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] _212_/X vssd vccd _032_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_34_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1502_A wire1503/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__A _185_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_991 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1871_A wire1871/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1969_A wire1970/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1888 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4210 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4243 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3640 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3531 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_788 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__095__A _095_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3294 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__542__B _542_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input170_A la_iena_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input268_A la_oenb_mprj[107] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input435_A mprj_dat_o_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_814 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput210 la_iena_mprj[55] vssd vccd _218_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_4_3749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input31_A la_data_out_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput221 la_iena_mprj[65] vssd vccd _228_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_23_1207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput232 la_iena_mprj[75] vssd vccd _238_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput243 la_iena_mprj[85] vssd vccd _248_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput254 la_iena_mprj[95] vssd vccd _258_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput265 la_oenb_mprj[104] vssd vccd wire1603/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput276 la_oenb_mprj[114] vssd vccd wire1592/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput287 la_oenb_mprj[124] vssd vccd wire1582/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput298 la_oenb_mprj[19] vssd vccd _516_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_586_ _586_/A _586_/B vssd vccd _586_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_16_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__436__C _436_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output487_A _490_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__452__B _452_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output654_A _024_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput706 _072_/Y vssd vccd la_data_in_mprj[89] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput717 _082_/Y vssd vccd la_data_in_mprj[99] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput728 _605_/X vssd vccd la_oenb_core[108] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1285_A wire1286/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput739 _615_/X vssd vccd la_oenb_core[118] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output821_A _574_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output919_A wire1208/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3290 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1452_A wire1453/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_2453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3851 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__362__B _362_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[6\]_A mprj_dat_i_user[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_304 _582_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_315 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_326 wire2078/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_337 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_440_ _568_/A _440_/B _440_/C vssd vccd _440_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_52_4051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_348 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_359 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__419__A_N _547_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_371_ _499_/A _371_/B _371_/C vssd vccd _371_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4068 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2100_A wire2101/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__553__A _553_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input385_A la_oenb_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_975 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__272__B _272_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input79_A la_data_out_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_2659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__447__B _447_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1033_A _516_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_569_ _569_/A _569_/B vssd vccd _569_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1200_A wire1201/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output771_A _528_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output869_A _334_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput503 wire1124/X vssd vccd la_data_in_core[20] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput514 wire1114/X vssd vccd la_data_in_core[30] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1667_A wire1667/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput525 wire1104/X vssd vccd la_data_in_core[40] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_48_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3446 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput536 wire1093/X vssd vccd la_data_in_core[50] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput547 wire1080/X vssd vccd la_data_in_core[60] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2662 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput558 _439_/X vssd vccd la_data_in_core[70] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput569 _449_/X vssd vccd la_data_in_core[80] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1834_A wire1834/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3872 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4300 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__357__B _357_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_216 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3698 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4326 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3783 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1801 wire1801/A vssd vccd _255_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_1_3708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2299 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1812 wire1812/A vssd vccd _334_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1823 wire1823/A vssd vccd _331_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1834 wire1834/A vssd vccd wire1834/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1845 wire1845/A vssd vccd _180_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input133_A la_iena_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2050_A wire2050/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1856 wire1856/A vssd vccd _173_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1867 wire1868/X vssd vccd _165_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1878 wire1878/A vssd vccd wire1878/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__548__A _548_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1889 wire1890/X vssd vccd _619_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1070 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_101 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_112 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input300_A la_oenb_mprj[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__267__B _267_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_123 mprj_dat_i_user[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_134 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_145 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_156 _219_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_423_ _551_/A _423_/B _423_/C vssd vccd _423_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_167 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_178 _400_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_189 _529_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__391__A_N _519_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_354_ _354_/A _354_/B vssd vccd _354_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_41_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__283__A _283_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_285_ _285_/A _285_/B vssd vccd _285_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1307 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1246 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2846 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1150_A wire1151/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput7 la_data_out_mprj[102] vssd vccd _471_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2686 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__177__B _177_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1415_A wire1416/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] _194_/X vssd vccd _014_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_51_138 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__193__A _193_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1784_A wire1784/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1951_A wire1952/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2542 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1108 _405_/X vssd vccd wire1108/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1119 _394_/X vssd vccd wire1119/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__368__A _368_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4196 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1150 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_070_ _070_/A vssd vccd _070_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_17_1194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2051 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2098_A wire2098/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__550__B _550_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_4112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input250_A la_iena_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input348_A la_oenb_mprj[64] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4156 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1620 wire1620/A vssd vccd _453_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1631 wire1631/A vssd vccd _442_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1642 wire1642/A vssd vccd wire1642/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1653 wire1653/A vssd vccd wire1653/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__278__A _278_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1664 wire1665/X vssd vccd wire1664/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1675 wire1675/A vssd vccd wire1675/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1686 wire1687/X vssd vccd _370_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1697 wire1697/A vssd vccd wire1697/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2650 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_406_ _406_/A_N _406_/B _406_/C vssd vccd _406_/X vssd vccd sky130_fd_sc_hd__and3b_4
XPHY_80 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_91 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_337_ _337_/A _337_/B vssd vccd _337_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__444__C _444_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_268_ _268_/A _268_/B vssd vccd _268_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output567_A _448_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire961 wire961/A vssd vccd _082_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_3609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire972 wire972/A vssd vccd _068_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire983 wire983/A vssd vccd _100_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_31_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4023 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire994 _587_/X vssd vccd wire994/X vssd vccd sky130_fd_sc_hd__buf_6
X_199_ _199_/A _199_/B vssd vccd _199_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1198_A wire1199/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__460__B _460_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4067 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output734_A _610_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1365_A wire1365/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output901_A _142_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] wire1333/X vssd vccd wire977/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_39_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1532_A wire1532/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__A _188_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[23\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1999_A wire2000/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire985_A wire985/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3602 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_12 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_23 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_34 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_867 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_45 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_56 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3668 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_67 mprj_dat_i_user[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_78 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_89 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__370__B _370_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__098__A _098_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[14\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__545__B _545_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input298_A la_oenb_mprj[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_122_ _122_/A vssd vccd _122_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_11_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__561__A _561_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_053_ _053_/A vssd vccd _053_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_27_4343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__280__B _280_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input61_A la_data_out_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4387 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3528 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2952 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4014 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2140 wire2140/A vssd vccd _464_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2151 wire2151/A vssd vccd wire2151/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2162 wire2163/X vssd vccd _452_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2173 wire2174/X vssd vccd _447_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2184 wire2185/X vssd vccd _442_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1450 wire1451/X vssd vccd wire1450/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2195 wire2195/A vssd vccd _308_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1461 wire1461/A vssd vccd wire1461/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1472 wire1473/X vssd vccd _328_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__439__C _439_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1483 wire1484/X vssd vccd wire1483/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1494 wire1495/X vssd vccd _323_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2595 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__455__B _455_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output684_A _052_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput10 la_data_out_mprj[105] vssd vccd _474_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_output851_A wire1266/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput21 la_data_out_mprj[115] vssd vccd _484_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_28_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput32 la_data_out_mprj[125] vssd vccd input32/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_11_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output949_A wire1303/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput43 la_data_out_mprj[1] vssd vccd _370_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput54 la_data_out_mprj[2] vssd vccd _371_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_50_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput65 la_data_out_mprj[3] vssd vccd _372_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1482_A wire1483/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput76 la_data_out_mprj[4] vssd vccd _373_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput87 la_data_out_mprj[5] vssd vccd _374_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__190__B _190_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput98 la_data_out_mprj[6] vssd vccd _375_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1747_A wire1748/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] _268_/X vssd vccd _088_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_0_2144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3702 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xmprj2_logic_high_inst wire2209/A vccd2 vssd2 mprj2_logic_high
XFILLER_11_4100 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__365__B _365_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_992 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__452__A_N _580_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3826 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput403 mprj_adr_o_core[23] vssd vccd wire1474/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput414 mprj_adr_o_core[4] vssd vccd wire1421/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput425 mprj_dat_o_core[13] vssd vccd wire1384/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_3550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput436 mprj_dat_o_core[23] vssd vccd wire1368/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput447 mprj_dat_o_core[4] vssd vccd wire1355/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput458 mprj_stb_o_core vssd vccd wire1343/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_1260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2130_A wire2131/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input213_A la_iena_mprj[58] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_959 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__556__A _556_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__275__B _275_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2090 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__291__A _291_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_105_ _105_/A vssd vccd _105_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4151 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_036_ _036_/A vssd vccd _036_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4048 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3483 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1063_A _472_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1280 wire1281/X vssd vccd wire1280/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1291 wire1292/X vssd vccd wire1291/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1230_A wire1231/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__475__A_N _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1328_A _249_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_406 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__185__B _185_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_4420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_491 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1697_A wire1697/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1864_A wire1864/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1906 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xmprj_logic_high_inst wire2204/A _395_/B _396_/B _397_/B _398_/B _399_/B _400_/B _401_/B
+ _402_/B _403_/B _404_/B wire2202/A _405_/B _406_/B _407_/B _408_/B _409_/B _410_/B
+ _411_/B _412_/B _413_/B _414_/B wire2200/A _415_/B _416_/B _417_/B _418_/B _419_/B
+ _420_/B _421_/B _422_/B _423_/B _424_/B wire2199/A _425_/B _426_/B _427_/B _428_/B
+ _429_/B _430_/B _431_/B wire2198/A wire2197/A wire2196/A wire2195/A wire2194/A wire2193/A
+ wire2192/A wire2191/A wire2190/A wire2188/A wire2187/A wire2185/A wire2183/A wire2181/A
+ wire2179/A wire2178/A wire2176/A wire2174/A wire2172/A wire2170/A wire2168/A wire2166/A
+ wire2164/A wire2161/A wire2158/A wire2155/A wire2154/A wire2151/A wire2148/A wire2145/A
+ wire2144/A wire2143/A wire2142/A _462_/B wire2141/A wire2140/A _311_/A wire2139/A
+ wire2138/A wire2136/A wire2135/A wire2134/A wire2132/A wire2131/A wire2129/A wire2127/A
+ wire2125/A _312_/A wire2123/A wire2122/A wire2120/A wire2118/A wire2116/A wire2114/A
+ wire2111/A wire2109/A wire2107/A wire2104/A _313_/A wire2101/A wire2098/A wire2096/A
+ wire2093/A wire2090/A wire2087/A wire2084/A wire2081/A wire2078/A wire2075/A _314_/A
+ _296_/A wire2072/A wire2068/A wire2065/A wire2063/A wire2061/A wire2059/A wire2057/A
+ wire2056/A wire2054/A wire2052/A _315_/A wire2051/A wire2050/A wire2048/A wire2046/A
+ wire2044/A wire2043/A wire2041/A wire2039/A wire2038/A wire2036/A _316_/A wire2035/A
+ wire2034/A wire2033/A wire2032/A wire2031/A wire2030/A wire2029/A _522_/B wire2028/A
+ _524_/B _317_/A wire2027/A _526_/B _527_/B _528_/B _529_/B _530_/B wire2026/A _532_/B
+ _533_/B _534_/B _318_/A wire2025/A _536_/B _537_/B _538_/B wire2024/A _540_/B _541_/B
+ _542_/B _543_/B _544_/B _319_/A _545_/B wire2023/A _547_/B _548_/B _549_/B _550_/B
+ _551_/B _552_/B _553_/B _554_/B _320_/A _555_/B _556_/B _557_/B _558_/B wire2022/A
+ wire2021/A wire2020/A wire2019/A wire2018/A wire2017/A _321_/A wire2016/A wire2015/A
+ wire2014/A wire2013/A wire2011/A wire2009/A wire2008/A wire2006/A wire2004/A wire2002/A
+ _322_/A wire2000/A wire1997/A wire1995/A wire1993/A wire1991/A wire1989/A wire1987/A
+ wire1985/A wire1983/A wire1980/A _323_/A wire1978/A wire1976/A wire1975/A wire1974/A
+ wire1972/A wire1971/A wire1970/A wire1968/A wire1966/A wire1964/A _324_/A wire1962/A
+ wire1958/A wire1956/A wire1954/A wire1952/A wire1949/A wire1947/A wire1944/A wire1942/A
+ wire1940/A wire1938/A _325_/A wire1936/A wire1933/A wire1930/A wire1927/A wire1924/A
+ wire1921/A wire1918/A wire1914/A wire1910/A wire1907/A _326_/A wire1904/A wire1901/A
+ wire1897/A wire1894/A wire1891/A wire1888/A wire1885/A wire1882/A wire1878/A wire1875/A
+ _327_/A wire1871/A wire1870/A wire1868/A wire1866/A wire1864/A wire1862/A wire1861/A
+ wire1860/A wire1858/A wire1857/A _328_/A wire1856/A wire1855/A wire1853/A wire1851/A
+ wire1849/A wire1848/A wire1846/A wire1845/A wire1844/A wire1843/A wire1842/A wire1841/A
+ wire1840/A wire1839/A wire1838/A wire1836/A wire1834/A wire1832/A wire1830/A wire1829/A
+ wire1828/A wire1827/A wire1826/A wire1825/A wire1824/A _196_/A _197_/A _198_/A _199_/A
+ _200_/A _201_/A _202_/A wire1823/A _203_/A wire1822/A wire1821/A wire1820/A wire1819/A
+ wire1818/A _209_/A _210_/A _211_/A _212_/A wire1817/A _213_/A _214_/A _215_/A _216_/A
+ _217_/A _218_/A _219_/A _220_/A _221_/A _222_/A wire1816/A _223_/A _224_/A _225_/A
+ _226_/A _227_/A _228_/A _229_/A wire1815/A wire1814/A wire1813/A wire1812/A wire1811/A
+ wire1810/A _234_/A _235_/A _236_/A _237_/A _238_/A _239_/A _240_/A _241_/A _242_/A
+ wire1809/A _243_/A wire1808/A wire1807/A _246_/A _247_/A _248_/A wire1806/A wire1805/A
+ wire1804/A _252_/A wire1803/A _253_/A wire1802/A wire1801/A wire1800/A wire1799/A
+ wire1798/A wire1797/A wire1796/A wire1794/A wire1792/A _337_/A wire1790/A wire1788/A
+ wire1786/A wire1784/A wire1783/A wire1781/A wire1779/A wire1777/A wire1776/A wire1774/A
+ _338_/A wire1772/A wire1770/A wire1768/A wire1766/A wire1764/A wire1762/A wire1760/A
+ wire1758/A wire1756/A wire1754/A _339_/A wire1752/A wire1750/A wire1748/A wire1745/A
+ wire1743/A wire1741/A wire1739/A wire1737/A wire1734/A wire1731/A _340_/A wire1728/A
+ wire1725/A wire1722/A _341_/A _342_/A _343_/A _344_/A _299_/A _345_/A _346_/A _347_/A
+ _348_/A _349_/A wire1719/A wire1718/A wire1717/A wire1716/A wire1715/A wire1714/A
+ wire1713/A wire1712/A wire1711/A wire1710/A wire1709/A wire1708/A wire1707/A wire1705/A
+ wire1703/A wire1701/A wire1699/A wire1697/A wire1695/A wire1693/A wire1691/A wire1689/A
+ wire1687/A wire1685/A wire1683/A wire1681/A wire1679/A wire1677/A wire1675/A wire1673/A
+ wire1671/A wire1669/A wire1667/A wire1665/A wire1662/A wire1660/A wire1658/A wire1656/A
+ wire1654/A wire1653/A wire1651/A wire1649/A wire1647/A wire1645/A wire1644/A wire1642/A
+ wire1640/A wire1638/A wire1636/A wire1634/A vccd1 vssd1 mprj_logic_high
XFILLER_2_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1215 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_995 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2583 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2080_A wire2081/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input163_A la_iena_mprj[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2178_A wire2178/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput200 la_iena_mprj[46] vssd vccd _209_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput211 la_iena_mprj[56] vssd vccd _219_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_44_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput222 la_iena_mprj[66] vssd vccd _229_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_0_365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput233 la_iena_mprj[76] vssd vccd _239_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input330_A la_oenb_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput244 la_iena_mprj[86] vssd vccd _249_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input428_A mprj_dat_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput255 la_iena_mprj[96] vssd vccd _259_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput266 la_oenb_mprj[105] vssd vccd wire1602/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input24_A la_data_out_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput277 la_oenb_mprj[115] vssd vccd wire1591/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput288 la_oenb_mprj[125] vssd vccd wire1581/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput299 la_oenb_mprj[1] vssd vccd _498_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_29_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2762 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__286__A _286_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_585_ _585_/A _585_/B vssd vccd _585_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3151 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__452__C _452_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput707 _155_/Y vssd vccd la_data_in_mprj[8] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput718 _156_/Y vssd vccd la_data_in_mprj[9] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput729 _606_/X vssd vccd la_oenb_core[109] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output647_A _018_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_019_ _019_/A vssd vccd _019_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1180_A wire1181/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1278_A wire1279/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output814_A _567_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1445_A wire1446/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] _224_/X vssd vccd _044_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_23_2498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__196__A _196_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_715 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3972 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1981_A wire1982/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[6\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_3077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1703 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_305 _579_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_316 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_327 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_338 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_349 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_370_ _498_/A _370_/B _370_/C vssd vccd _370_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2623 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__553__B _553_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input280_A la_oenb_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input378_A la_oenb_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_542 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__447__C _447_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_568_ _568_/A _568_/B vssd vccd _568_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1026_A _523_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1702 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output597_A _088_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2578 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_499_ _499_/A _499_/B vssd vccd _499_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__B _463_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output764_A wire1027/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1395_A wire1396/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput504 wire1123/X vssd vccd la_data_in_core[21] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output931_A wire1166/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput515 wire1113/X vssd vccd la_data_in_core[31] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput526 wire1103/X vssd vccd la_data_in_core[41] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput537 wire1092/X vssd vccd la_data_in_core[51] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput548 wire1079/X vssd vccd la_data_in_core[61] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput559 _440_/X vssd vccd la_data_in_core[71] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2674 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1827_A wire1827/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1911 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1944 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__B _373_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1207 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_928 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4338 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3795 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1802 wire1802/A vssd vccd _254_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1813 wire1813/A vssd vccd _232_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1824 wire1824/A vssd vccd _195_/A vssd vccd sky130_fd_sc_hd__buf_4
Xwire1835 wire1836/X vssd vccd _187_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1846 wire1846/A vssd vccd _179_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3580 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1857 wire1857/A vssd vccd _172_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1868 wire1868/A vssd vccd wire1868/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1879 wire1880/X vssd vccd _622_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__548__B _548_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2043_A wire2043/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input126_A la_data_out_mprj[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_102 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_113 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_124 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_135 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_146 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_157 _220_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_422_ _550_/A _422_/B _422_/C vssd vccd _422_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_168 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_179 _550_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__564__A _564_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
X_353_ _353_/A _353_/B vssd vccd _353_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_14_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3154 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input91_A la_data_out_mprj[63] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_284_ _284_/A _284_/B vssd vccd _284_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_48_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[7\] mprj_dat_i_user[7] max_length1311/X vssd vccd _121_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1258 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3283 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output512_A wire1115/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput8 la_data_out_mprj[103] vssd vccd _472_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__458__B _458_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2698 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1143_A _371_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1408_A wire1408/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2222 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] _187_/X vssd vccd _007_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XANTENNA__193__B _193_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1777_A wire1777/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1944_A wire1944/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__409__A_N _409_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2554 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2482 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1109 _404_/X vssd vccd wire1109/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_4476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__368__B _368_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_136 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1474 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_51_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4028 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1026 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2626 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1059 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3802 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput890 _132_/Y vssd vccd mprj_dat_i_core[18] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2160_A wire2161/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input243_A la_iena_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4168 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3434 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1610 wire1610/A vssd vccd _230_/B vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__559__A _559_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1621 wire1621/A vssd vccd _452_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1632 wire1632/A vssd vccd _441_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1643 wire1644/X vssd vccd _390_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1654 wire1654/A vssd vccd _303_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input410_A mprj_adr_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__278__B _278_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1665 wire1665/A vssd vccd wire1665/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1676 wire1677/X vssd vccd _302_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1687 wire1687/A vssd vccd wire1687/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1698 wire1699/X vssd vccd _301_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__294__A _294_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_405_ _405_/A_N _405_/B _405_/C vssd vccd _405_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_19_2662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_70 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_92 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_336_ _336_/A _336_/B vssd vccd _336_/X vssd vccd sky130_fd_sc_hd__and2_4
X_267_ _267_/A _267_/B vssd vccd _267_/X vssd vccd sky130_fd_sc_hd__and2_4
Xwire962 wire962/A vssd vccd _078_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire973 wire973/A vssd vccd _067_/A vssd vccd sky130_fd_sc_hd__buf_6
X_198_ _198_/A _198_/B vssd vccd _198_/X vssd vccd sky130_fd_sc_hd__and2_2
Xwire984 wire984/A vssd vccd _098_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire995 _586_/X vssd vccd wire995/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_26_4035 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__460__C _460_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1093_A wire1094/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4079 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output727_A _604_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1358_A wire1358/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__188__B _188_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1525_A wire1526/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_651 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2615 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1894_A wire1894/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_13 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_846 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_24 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_35 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_46 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1947 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_57 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_68 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_79 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__C _370_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__381__A_N _509_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2215 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1803 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2006_A wire2006/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_3124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_121_ _121_/A vssd vccd _121_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input193_A la_iena_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_052_ _052_/A vssd vccd _052_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__561__B _561_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2456 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4355 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input360_A la_oenb_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input458_A mprj_stb_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4399 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input54_A la_data_out_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3687 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2130 wire2131/X vssd vccd _471_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2141 wire2141/A vssd vccd _463_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__289__A _289_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2152 wire2153/X vssd vccd _455_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2760 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2163 wire2164/X vssd vccd wire2163/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2174 wire2174/A vssd vccd wire2174/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1440 wire1441/X vssd vccd wire1440/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2185 wire2185/A vssd vccd wire2185/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1451 wire1451/A vssd vccd wire1451/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2196 wire2196/A vssd vccd _434_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1462 wire1463/X vssd vccd _330_/B vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_21_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1473 wire1474/X vssd vccd wire1473/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1484 wire1484/A vssd vccd wire1484/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1495 wire1496/X vssd vccd wire1495/X vssd vccd sky130_fd_sc_hd__buf_6
Xpowergood_check vccd vdda1 vdda2 output954/A output952/A vssa1 vssd vssa2 mgmt_protect_hv
XFILLER_19_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__455__C _455_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1106_A _407_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_319_ _319_/A _319_/B vssd vccd _319_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput11 la_data_out_mprj[106] vssd vccd _475_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput22 la_data_out_mprj[116] vssd vccd input22/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput33 la_data_out_mprj[126] vssd vccd input33/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__471__B _471_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput44 la_data_out_mprj[20] vssd vccd _389_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_out_mprj[30] vssd vccd _399_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3680 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output844_A _595_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput66 la_data_out_mprj[40] vssd vccd _409_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput77 la_data_out_mprj[50] vssd vccd _419_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput88 la_data_out_mprj[60] vssd vccd _429_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput99 la_data_out_mprj[70] vssd vccd input99/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_2717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1475_A wire1476/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] wire1323/X vssd vccd wire966/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_48_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3236 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3258 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1642_A wire1642/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__199__A _199_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1907_A wire1907/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1466 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4292 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4156 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3488 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__B _381_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_514 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4252 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput404 mprj_adr_o_core[24] vssd vccd wire1471/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput415 mprj_adr_o_core[5] vssd vccd wire1416/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput426 mprj_dat_o_core[14] vssd vccd wire1382/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_3781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput437 mprj_dat_o_core[24] vssd vccd wire1367/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput448 mprj_dat_o_core[5] vssd vccd wire1353/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput459 mprj_we_o_core vssd vccd wire1341/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_798 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2123_A wire2123/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input206_A la_iena_mprj[51] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1032 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2687 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__572__A _572_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_104_ _104_/A vssd vccd _104_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_8_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__291__B _291_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_035_ _035_/A vssd vccd _035_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4163 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3495 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1056_A _479_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1270 _316_/X vssd vccd wire1270/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1281 wire1282/X vssd vccd wire1281/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1292 wire1293/X vssd vccd wire1292/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__466__B _466_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1223_A wire1224/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output794_A wire1007/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_971 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2754 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1857_A wire1857/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__376__B _376_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_B wire1318/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_985 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2073_A wire2074/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input156_A la_iena_mprj[121] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput201 la_iena_mprj[47] vssd vccd _210_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_2_4143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput212 la_iena_mprj[57] vssd vccd _220_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput223 la_iena_mprj[67] vssd vccd wire1610/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput234 la_iena_mprj[77] vssd vccd _240_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput245 la_iena_mprj[87] vssd vccd _250_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput256 la_iena_mprj[97] vssd vccd _260_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_2_3453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput267 la_oenb_mprj[106] vssd vccd wire1601/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input323_A la_oenb_mprj[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput278 la_oenb_mprj[116] vssd vccd wire1590/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput289 la_oenb_mprj[126] vssd vccd wire1580/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__567__A _567_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input17_A la_data_out_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__286__B _286_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_584_ _584_/A _584_/B vssd vccd _584_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_16_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[87\]_B wire1327/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2927 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2495 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput708 _073_/Y vssd vccd la_data_in_mprj[90] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput719 wire1053/X vssd vccd la_oenb_core[0] vssd vccd sky130_fd_sc_hd__buf_8
X_018_ _018_/A vssd vccd _018_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA_output542_A wire1085/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2867 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1173_A _362_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[11\]_B _174_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__442__A_N _570_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output807_A _561_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1438_A wire1439/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] _217_/X vssd vccd _037_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_1550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_4565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3984 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[78\]_B _241_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1974_A wire1974/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input9_A la_data_out_mprj[104] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_306 _565_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_317 wire1985/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_328 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_339 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3450 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1972 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_999 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input273_A la_oenb_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_2381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__465__A_N _593_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input440_A mprj_dat_o_core[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3272 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__297__A _297_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3203 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_567_ _567_/A _567_/B vssd vccd _567_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_18_2568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_498_ _498_/A _498_/B vssd vccd _498_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output492_A _495_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1019_A _536_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__463__C _463_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2194 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2779 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output757_A wire1033/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1290_A wire1291/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput505 wire1122/X vssd vccd la_data_in_core[22] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput516 wire1112/X vssd vccd la_data_in_core[32] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput527 wire1102/X vssd vccd la_data_in_core[42] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput538 wire1091/X vssd vccd la_data_in_core[52] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output924_A wire1249/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput549 wire1078/X vssd vccd la_data_in_core[62] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1722_A wire1722/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__000__A _000_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2092 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__488__A_N _616_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1803 wire1803/A vssd vccd _336_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1814 wire1814/A vssd vccd _231_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1825 wire1825/A vssd vccd _194_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1836 wire1836/A vssd vccd wire1836/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3570 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1847 wire1848/X vssd vccd _178_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1858 wire1858/A vssd vccd _171_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1869 wire1870/X vssd vccd _164_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_318 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_103 mprj_dat_i_user[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_114 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2036_A wire2036/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_125 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input119_A la_data_out_mprj[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_421_ _549_/A _421_/B _421_/C vssd vccd _421_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_136 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_147 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_158 _220_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_169 _229_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__564__B _564_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_352_ _352_/A _352_/B vssd vccd _352_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_user_to_mprj_in_gates\[126\]_B _289_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2203_A wire2204/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_3193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_283_ _283_/A _283_/B vssd vccd _283_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input390_A mprj_adr_o_core[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input84_A la_data_out_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__580__A _580_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3470 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3295 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput9 la_data_out_mprj[104] vssd vccd _473_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2508 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__458__C _458_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output505_A wire1122/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1136_A _378_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_619_ _619_/A _619_/B vssd vccd _619_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__B _474_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_2354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[117\]_B _280_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1303_A wire1304/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] _180_/X vssd vccd _000_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_31_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1672_A wire1673/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3223 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1937_A wire1938/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2494 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1094 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_A mprj_dat_i_user[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_148 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3008 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__B _384_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[108\]_B _271_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1038 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput880 wire1306/X vssd vccd mprj_cyc_o_user vssd vccd sky130_fd_sc_hd__buf_8
Xoutput891 _133_/Y vssd vccd mprj_dat_i_core[19] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1600 wire1600/A vssd vccd _604_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1611 input22/X vssd vccd _485_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_21_3446 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__559__B _559_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1622 wire1622/A vssd vccd _451_/C vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input236_A la_iena_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2153_A wire2154/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[17\]_A mprj_dat_i_user[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1633 wire1633/A vssd vccd _440_/C vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_4_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1644 wire1644/A vssd vccd wire1644/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1655 wire1656/X vssd vccd _384_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1167 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1666 wire1667/X vssd vccd _379_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4032 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1677 wire1677/A vssd vccd wire1677/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1688 wire1689/X vssd vccd _369_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1699 wire1699/A vssd vccd wire1699/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input403_A mprj_adr_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__575__A _575_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_170 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__294__B _294_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_404_ _532_/A _404_/B _404_/C vssd vccd _404_/X vssd vccd sky130_fd_sc_hd__and3b_4
XPHY_60 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_71 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_82 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_335_ _335_/A _335_/B vssd vccd _335_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_30_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_266_ _266_/A _266_/B vssd vccd _266_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_3840 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire963 wire963/A vssd vccd _077_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_26_4003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_197_ _197_/A _197_/B vssd vccd _197_/X vssd vccd sky130_fd_sc_hd__and2_2
Xwire974 wire974/A vssd vccd _066_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire985 wire985/A vssd vccd _097_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire996 _558_/X vssd vccd wire996/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_26_4047 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2623 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__469__B _469_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1253_A _328_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_936 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1420_A wire1421/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1518_A wire1519/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_14 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3784 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_25 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1887_A wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_36 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_47 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_58 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_69 mprj_dat_i_user[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1694 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3891 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__379__B _379_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_696 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_120_ _120_/A vssd vccd _120_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_051_ _051_/A vssd vccd _051_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input186_A la_iena_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input353_A la_oenb_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input47_A la_data_out_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2120 wire2120/A vssd vccd wire2120/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_4027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2131 wire2131/A vssd vccd wire2131/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__289__B _289_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2142 wire2142/A vssd vccd _461_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2153 wire2154/X vssd vccd wire2153/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2164 wire2164/A vssd vccd wire2164/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1430 wire1431/X vssd vccd wire1430/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2175 wire2176/X vssd vccd _446_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1441 wire1441/A vssd vccd wire1441/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_2614 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2186 wire2187/X vssd vccd _441_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1452 wire1453/X vssd vccd _332_/B vssd vccd sky130_fd_sc_hd__buf_8
Xwire2197 wire2197/A vssd vccd _433_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1463 wire1464/X vssd vccd wire1463/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1474 wire1474/A vssd vccd wire1474/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1485 wire1486/X vssd vccd _306_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1496 wire1497/X vssd vccd wire1496/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_318_ _318_/A _318_/B vssd vccd _318_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1001_A _555_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output572_A _452_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput12 la_data_out_mprj[107] vssd vccd _476_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_35_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput23 la_data_out_mprj[117] vssd vccd _486_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput34 la_data_out_mprj[127] vssd vccd input34/X vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput45 la_data_out_mprj[21] vssd vccd _390_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__471__C _471_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_249_ _249_/A _249_/B vssd vccd _249_/X vssd vccd sky130_fd_sc_hd__and2_4
Xinput56 la_data_out_mprj[31] vssd vccd _400_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput67 la_data_out_mprj[41] vssd vccd _410_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3692 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput78 la_data_out_mprj[51] vssd vccd _420_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput89 la_data_out_mprj[61] vssd vccd _430_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output837_A _588_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1370_A wire1370/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1468_A wire1469/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] wire1330/X vssd vccd wire973/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_44_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__199__B _199_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1635_A wire1636/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3846 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_600 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3570 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3478 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__C _381_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4264 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput405 mprj_adr_o_core[25] vssd vccd wire1466/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput416 mprj_adr_o_core[6] vssd vccd wire1411/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput427 mprj_dat_o_core[15] vssd vccd wire1380/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput438 mprj_dat_o_core[25] vssd vccd wire1366/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput449 mprj_dat_o_core[6] vssd vccd wire1351/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input101_A la_data_out_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1055 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__572__B _572_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_103_ _103_/A vssd vccd _103_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4131 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_034_ _034_/A vssd vccd _034_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_7_4225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4175 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2762 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1260 _321_/X vssd vccd wire1260/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1271 wire1272/X vssd vccd wire1271/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1282 wire1283/X vssd vccd wire1282/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_2394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1293 _302_/X vssd vccd wire1293/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1049_A _501_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1743 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__466__C _466_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1100 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1216_A _350_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output787_A _543_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__A_N _499_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__B _482_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output954_A output954/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[12\] mprj_dat_i_user[12] max_length1311/X vssd vccd _126_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_12_3787 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1752_A wire1752/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3966 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] _273_/X vssd vccd wire989/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_27_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1108 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_1239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__392__B _392_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_A mprj_dat_i_user[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput202 la_iena_mprj[48] vssd vccd _211_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput213 la_iena_mprj[58] vssd vccd _221_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput224 la_iena_mprj[68] vssd vccd wire1609/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input149_A la_iena_mprj[115] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2066_A wire2067/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput235 la_iena_mprj[78] vssd vccd _241_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput246 la_iena_mprj[88] vssd vccd _251_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_24_2979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput257 la_iena_mprj[98] vssd vccd _261_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput268 la_oenb_mprj[107] vssd vccd wire1600/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput279 la_oenb_mprj[117] vssd vccd wire1589/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_4108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__567__B _567_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input316_A la_oenb_mprj[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1039 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_583_ _583_/A _583_/B vssd vccd _583_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__394__A_N _522_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2619 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__A _583_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1306 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_3175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2939 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput709 _074_/Y vssd vccd la_data_in_mprj[91] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_7_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_017_ _017_/A vssd vccd _017_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_46_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output535_A wire1141/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1166_A wire1167/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__477__B _477_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1090 _422_/X vssd vccd wire1090/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] _210_/X vssd vccd _030_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_1540 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1228 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1967_A wire1968/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1147 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] _172_/X vssd vccd _156_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_41_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__387__B _387_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1232 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_307 wire2116/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_318 wire1985/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_329 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_4174 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3462 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3326 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1003 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4320 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4364 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2183_A wire2183/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input266_A la_oenb_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input433_A mprj_dat_o_core[20] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__578__A _578_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2503 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_566_ _566_/A _566_/B vssd vccd _566_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_497_ _497_/A _497_/B vssd vccd _497_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2140 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output485_A wire1133/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1423 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput506 wire1121/X vssd vccd la_data_in_core[23] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3427 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput517 wire1111/X vssd vccd la_data_in_core[33] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput528 wire1101/X vssd vccd la_data_in_core[43] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1283_A _304_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput539 wire1090/X vssd vccd la_data_in_core[53] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_10_1191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output917_A wire1214/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1450_A wire1451/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1715_A wire1715/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1535 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1804 wire1804/A vssd vccd _251_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1815 wire1815/A vssd vccd _230_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1826 wire1826/A vssd vccd _193_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1837 wire1838/X vssd vccd _186_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1848 wire1848/A vssd vccd wire1848/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1859 wire1860/X vssd vccd _170_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2870 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_104 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_115 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_126 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_420_ _420_/A_N _420_/B _420_/C vssd vccd _420_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_137 _547_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_148 _209_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3568 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_159 _221_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2029_A wire2029/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_351_ _351_/A _351_/B vssd vccd _351_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_36_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4160 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_282_ _282_/A _282_/B vssd vccd _282_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__432__A_N _560_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input383_A la_oenb_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__580__B _580_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input77_A la_data_out_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4036 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3482 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__101__A _101_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_618_ _618_/A _618_/B vssd vccd _618_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1031_A _518_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1129_A _384_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_549_ _549_/A _549_/B vssd vccd _549_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2366 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3988 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output867_A _332_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1498_A wire1499/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__B _490_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1832_A wire1832/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4412 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2359 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[26\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__455__A_N _583_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__384__C _384_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1000 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1938 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput870 _307_/X vssd vccd mprj_adr_o_user[2] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput881 _114_/Y vssd vccd mprj_dat_i_core[0] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput892 _115_/Y vssd vccd mprj_dat_i_core[1] vssd vccd sky130_fd_sc_hd__buf_8
Xwire1601 wire1601/A vssd vccd _603_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1612 wire1612/A vssd vccd _189_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3458 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1623 wire1623/A vssd vccd _450_/C vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_user_wb_dat_gates\[17\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1634 wire1634/A vssd vccd _304_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1645 wire1645/A vssd vccd _389_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input131_A la_data_out_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1656 wire1656/A vssd vccd wire1656/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2146_A wire2147/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1667 wire1667/A vssd vccd wire1667/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input229_A la_iena_mprj[72] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1678 wire1679/X vssd vccd _374_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1689 wire1689/A vssd vccd wire1689/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__575__B _575_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_403_ _531_/A _403_/B _403_/C vssd vccd _403_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_26_182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_50 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_3229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_61 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_83 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_94 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_334_ _334_/A _334_/B vssd vccd _334_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__A _591_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_265_ _265_/A _265_/B vssd vccd _265_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire964 wire964/A vssd vccd _076_/A vssd vccd sky130_fd_sc_hd__buf_6
X_196_ _196_/A _196_/B vssd vccd _196_/X vssd vccd sky130_fd_sc_hd__and2_4
Xwire975 wire975/A vssd vccd _064_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire986 wire986/A vssd vccd _096_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire997 wire998/X vssd vccd wire997/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1079_A _430_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__469__C _469_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1246_A wire1247/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__478__A_N _478_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__B _485_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1413_A wire1414/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3763 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_15 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_26 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_37 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_48 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1782_A wire1783/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_59 mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1348 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__006__A _006_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2320 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__379__C _379_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__395__B _395_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3295 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_050_ _050_/A vssd vccd _050_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_49_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2096_A wire2096/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input179_A la_iena_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input346_A la_oenb_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2110 wire2111/X vssd vccd _481_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2121 wire2122/X vssd vccd _476_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2132 wire2132/A vssd vccd _470_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2143 wire2143/A vssd vccd _460_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3316 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2154 wire2154/A vssd vccd wire2154/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1420 wire1421/X vssd vccd wire1420/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2165 wire2166/X vssd vccd _451_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1431 wire1431/A vssd vccd wire1431/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2176 wire2176/A vssd vccd wire2176/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1442 wire1443/X vssd vccd _334_/B vssd vccd sky130_fd_sc_hd__buf_8
Xwire2187 wire2187/A vssd vccd wire2187/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1453 wire1454/X vssd vccd wire1453/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2198 wire2198/A vssd vccd _432_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__586__A _586_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1464 wire1465/X vssd vccd wire1464/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1475 wire1476/X vssd vccd _327_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1486 wire1487/X vssd vccd wire1486/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1497 wire1497/A vssd vccd wire1497/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_317_ _317_/A _317_/B vssd vccd _317_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_50_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput13 la_data_out_mprj[108] vssd vccd _477_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput24 la_data_out_mprj[118] vssd vccd _487_/C vssd vccd sky130_fd_sc_hd__buf_4
X_248_ _248_/A _248_/B vssd vccd _248_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_7_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput35 la_data_out_mprj[12] vssd vccd _381_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput46 la_data_out_mprj[22] vssd vccd _391_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_output565_A _446_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput57 la_data_out_mprj[32] vssd vccd _401_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput68 la_data_out_mprj[42] vssd vccd _411_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput79 la_data_out_mprj[52] vssd vccd _421_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
X_179_ _179_/A _179_/B vssd vccd _179_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1196_A wire1197/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output732_A _608_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1803 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] _240_/X vssd vccd _060_/A vssd vccd
+ sky130_fd_sc_hd__nand2_8
XFILLER_38_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1530_A wire1530/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1628_A wire1628/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4504 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1997_A wire1997/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire983_A wire983/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput406 mprj_adr_o_core[26] vssd vccd wire1461/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput417 mprj_adr_o_core[7] vssd vccd wire1408/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput428 mprj_dat_o_core[16] vssd vccd wire1378/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput439 mprj_dat_o_core[26] vssd vccd wire1365/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4047 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2109_A wire2109/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input296_A la_oenb_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_102_ _102_/A vssd vccd _102_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_2211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_033_ _033_/A vssd vccd _033_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_27_4143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2299 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4187 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3475 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2846 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1250 _338_/X vssd vccd wire1250/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1261 _320_/X vssd vccd wire1261/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1272 wire1273/X vssd vccd wire1272/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1283 _304_/X vssd vccd wire1283/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1294 wire1295/X vssd vccd wire1294/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1209_A wire1210/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output682_A _050_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__482__C _482_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output947_A wire1284/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1480_A wire1481/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1912_A wire1913/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_3989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] wire1316/X vssd vccd wire992/A
+ vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_26_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3508 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1999 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__392__C _392_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3232 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[9\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3276 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2564 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput203 la_iena_mprj[49] vssd vccd _212_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_user_to_mprj_in_gates\[9\]_B _172_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput214 la_iena_mprj[59] vssd vccd _222_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3422 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput225 la_iena_mprj[69] vssd vccd _232_/B vssd vccd sky130_fd_sc_hd__buf_4
Xinput236 la_iena_mprj[79] vssd vccd _242_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput247 la_iena_mprj[89] vssd vccd _252_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput258 la_iena_mprj[99] vssd vccd _262_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_5_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput269 la_oenb_mprj[108] vssd vccd _477_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_2721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2059_A wire2059/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input211_A la_iena_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_582_ _582_/A _582_/B vssd vccd _582_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_29_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input309_A la_oenb_mprj[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__583__B _583_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_016_ _016_/A vssd vccd _016_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__104__A _104_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output528_A wire1101/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1061_A _474_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1159_A wire1160/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1080 _429_/X vssd vccd wire1080/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_4523 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1091 _421_/X vssd vccd wire1091/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1326_A _251_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1596 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__493__B _493_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_740 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1695_A wire1695/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1115 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1738 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1862_A wire1862/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3108 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_512 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_308 wire2209/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_4131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_319 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_length1562_A _416_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_4186 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_239 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3316 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1015 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4376 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input161_A la_iena_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3434 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2176_A wire2176/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input259_A la_iena_mprj[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2755 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2023 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__578__B _578_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input426_A mprj_dat_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input22_A la_data_out_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__594__A _594_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_565_ _565_/A _565_/B vssd vccd _565_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_1883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_496_ _624_/A _496_/B _496_/C vssd vccd _496_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2152 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_2283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output478_A _482_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput507 wire1120/X vssd vccd la_data_in_core[24] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3356 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput518 wire1110/X vssd vccd la_data_in_core[34] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput529 wire1100/X vssd vccd la_data_in_core[44] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output645_A _016_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1276_A _313_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output812_A _566_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__B _488_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1443_A wire1444/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1708_A wire1708/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3940 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_max_length1310_A _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__384__A_N _512_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4455 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1547 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1306 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__398__B _398_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1805 wire1805/A vssd vccd _250_/A vssd vccd sky130_fd_sc_hd__buf_4
Xwire1816 wire1816/A vssd vccd _333_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1827 wire1827/A vssd vccd _330_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1838 wire1838/A vssd vccd wire1838/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1849 wire1849/A vssd vccd _177_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_1052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_105 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_116 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_127 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_138 _556_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_149 _210_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_350_ _350_/A _350_/B vssd vccd _350_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_281_ _281_/A _281_/B vssd vccd _281_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_14_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_2445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input376_A la_oenb_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3507 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4048 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__589__A _589_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_617_ _617_/A _617_/B vssd vccd _617_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_45_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_548_ _548_/A _548_/B vssd vccd _548_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1024_A _530_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output595_A _086_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_479_ _479_/A_N _479_/B _479_/C vssd vccd _479_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_31_2501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output762_A wire1029/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__490__C _490_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1393_A wire1393/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2430 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1658_A wire1658/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__499__A _499_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3916 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3444 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_17_1143 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3488 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput860 wire1256/X vssd vccd mprj_adr_o_user[20] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput871 _335_/X vssd vccd mprj_adr_o_user[30] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2034 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput882 _124_/Y vssd vccd mprj_dat_i_core[10] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput893 _134_/Y vssd vccd mprj_dat_i_core[20] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__202__A _202_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1602 wire1602/A vssd vccd _602_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_2089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1613 wire1613/A vssd vccd _188_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1624 wire1624/A vssd vccd _449_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1635 wire1636/X vssd vccd _394_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1646 wire1647/X vssd vccd _388_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1657 wire1658/X vssd vccd _383_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1668 wire1669/X vssd vccd _378_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1679 wire1679/A vssd vccd wire1679/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2041_A wire2041/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input124_A la_data_out_mprj[93] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2139_A wire2139/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_402_ _530_/A _402_/B _402_/C vssd vccd _402_/X vssd vccd sky130_fd_sc_hd__and3b_2
XPHY_40 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_3388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_73 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_333_ _333_/A _333_/B vssd vccd _333_/X vssd vccd sky130_fd_sc_hd__and2_4
XPHY_84 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_95 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__591__B _591_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_264_ _264_/A _264_/B vssd vccd _264_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_195_ _195_/A _195_/B vssd vccd _195_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_6_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire965 wire965/A vssd vccd _075_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire976 wire976/A vssd vccd _063_/A vssd vccd sky130_fd_sc_hd__buf_6
Xuser_wb_dat_gates\[5\] mprj_dat_i_user[5] max_length1311/X vssd vccd _119_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
Xwire987 wire987/A vssd vccd _095_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire998 _557_/X vssd vccd wire998/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2658 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output510_A wire1117/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output608_A _098_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1141_A _373_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1239_A wire1240/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4410 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__485__C _485_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1406_A wire1407/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] _185_/X vssd vccd _005_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_32_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_3775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_16 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_27 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_38 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_49 mprj_dat_i_user[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_371 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1775_A wire1776/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1942_A wire1942/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__422__A_N _550_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1686 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1274 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__395__C _395_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_2426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1714 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2089_A wire2090/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_4154 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2100 wire2101/X vssd vccd wire2100/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput690 _057_/Y vssd vccd la_data_in_mprj[74] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2111 wire2111/A vssd vccd wire2111/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input241_A la_iena_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2122 wire2122/A vssd vccd wire2122/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2133 wire2134/X vssd vccd _469_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input339_A la_oenb_mprj[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2144 wire2144/A vssd vccd _459_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1410 wire1411/X vssd vccd wire1410/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2155 wire2155/A vssd vccd _310_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1421 wire1421/A vssd vccd wire1421/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2166 wire2166/A vssd vccd wire2166/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1432 wire1433/X vssd vccd _335_/B vssd vccd sky130_fd_sc_hd__buf_8
Xwire2177 wire2178/X vssd vccd _445_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1443 wire1444/X vssd vccd wire1443/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire2188 wire2188/A vssd vccd _440_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1454 wire1455/X vssd vccd wire1454/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2199 wire2199/A vssd vccd _307_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1465 wire1466/X vssd vccd wire1465/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1476 wire1476/A vssd vccd wire1476/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__586__B _586_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1487 wire1488/X vssd vccd wire1487/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1498 wire1499/X vssd vccd _322_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_316_ _316_/A _316_/B vssd vccd _316_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3948 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__107__A _107_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput14 la_data_out_mprj[109] vssd vccd _478_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
X_247_ _247_/A _247_/B vssd vccd _247_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput25 la_data_out_mprj[119] vssd vccd input25/X vssd vccd sky130_fd_sc_hd__buf_6
Xinput36 la_data_out_mprj[13] vssd vccd _382_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput47 la_data_out_mprj[23] vssd vccd _392_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput58 la_data_out_mprj[33] vssd vccd _402_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput69 la_data_out_mprj[43] vssd vccd _412_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_13_1360 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_178_ _178_/A _178_/B vssd vccd _178_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output558_A _439_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1091_A _421_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__445__A_N _573_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output725_A _602_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1356_A wire1357/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4491 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__B _496_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1523_A wire1524/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4516 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1892_A wire1893/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_646 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire976_A wire976/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[32\]_B _195_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput407 mprj_adr_o_core[27] vssd vccd wire1456/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput418 mprj_adr_o_core[8] vssd vccd wire1404/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput429 mprj_dat_o_core[17] vssd vccd wire1377/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[99\]_B wire1317/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2004_A wire2004/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_101_ _101_/A vssd vccd _101_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_36_1393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input191_A la_iena_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input289_A la_oenb_mprj[126] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2223 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_032_ _032_/A vssd vccd _032_/Y vssd vccd sky130_fd_sc_hd__inv_2
XANTENNA__468__A_N _596_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input456_A mprj_sel_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_4199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input52_A la_data_out_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__597__A _597_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1240 _342_/X vssd vccd wire1240/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1251 wire1252/X vssd vccd wire1251/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1262 wire1263/X vssd vccd wire1262/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1273 _315_/X vssd vccd wire1273/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1284 wire1285/X vssd vccd wire1284/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_2446 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1295 wire1296/X vssd vccd wire1295/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1104_A _409_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output842_A _593_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1473_A wire1474/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[14\]_B _177_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1640_A wire1640/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3852 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1738_A wire1739/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_3957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__300__A _300_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1905_A wire1906/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_900 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3288 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3802 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput204 la_iena_mprj[4] vssd vccd _167_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput215 la_iena_mprj[5] vssd vccd _168_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_6_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput226 la_iena_mprj[6] vssd vccd _169_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4096 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput237 la_iena_mprj[7] vssd vccd _170_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput248 la_iena_mprj[8] vssd vccd _171_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2711 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput259 la_iena_mprj[9] vssd vccd _172_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__210__A _210_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3180 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_581_ _581_/A _581_/B vssd vccd _581_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input204_A la_iena_mprj[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2121_A wire2122/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1600 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_015_ _015_/A vssd vccd _015_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__120__A _120_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1070 _465_/X vssd vccd wire1070/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1081 _428_/X vssd vccd wire1081/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1092 _420_/X vssd vccd wire1092/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_14_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1221_A wire1222/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output792_A wire1009/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1319_A _258_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__493__C _493_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3586 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1688_A wire1689/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1127 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1855_A wire1855/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_3765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1328 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_309 _380_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__205__A _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4158 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input154_A la_iena_mprj[11] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2071_A wire2072/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2169_A wire2170/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3479 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input321_A la_oenb_mprj[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input419_A mprj_adr_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input15_A la_data_out_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__594__B _594_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1873 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_564_ _564_/A _564_/B vssd vccd _564_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4118 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_495_ _623_/A _495_/B _495_/C vssd vccd _495_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2874 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4108 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput508 wire1119/X vssd vccd la_data_in_core[25] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput519 wire1109/X vssd vccd la_data_in_core[35] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output540_A wire1089/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output638_A _010_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1171_A wire1172/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_ack_gate mprj_ack_i_user max_length1310/X vssd vccd _146_/A vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_wire1269_A wire1270/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3800 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__488__C _488_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output805_A _559_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1436_A wire1436/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] _215_/X vssd vccd _035_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_48_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_888 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3784 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1227 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4084 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1972_A wire1972/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__025__A _025_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3952 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4467 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_A mprj_dat_i_user[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1806 wire1806/A vssd vccd _249_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_41_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input7_A la_data_out_mprj[102] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1559 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__398__C _398_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1817 wire1817/A vssd vccd _332_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1828 wire1828/A vssd vccd _192_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1839 wire1839/A vssd vccd _185_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_106 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_117 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_128 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_139 _556_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_280_ _280_/A _280_/B vssd vccd _280_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input271_A la_oenb_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3519 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input369_A la_oenb_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1491 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__589__B _589_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_616_ _616_/A _616_/B vssd vccd _616_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_40_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_547_ _547_/A _547_/B vssd vccd _547_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_35_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_478_ _478_/A_N _478_/B _478_/C vssd vccd _478_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output490_A _493_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output588_A wire1068/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3692 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output755_A wire1035/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2442 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output922_A wire1198/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__499__B _499_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_3928 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4364 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1720_A wire1721/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3746 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3456 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput850 wire1268/X vssd vccd mprj_adr_o_user[11] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_4275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput861 _326_/X vssd vccd mprj_adr_o_user[21] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput872 _336_/X vssd vccd mprj_adr_o_user[31] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput883 _125_/Y vssd vccd mprj_dat_i_core[11] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput894 _135_/Y vssd vccd mprj_dat_i_core[21] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1603 wire1603/A vssd vccd _601_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_4071 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1614 wire1614/A vssd vccd _187_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1625 wire1625/A vssd vccd _448_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1636 wire1636/A vssd vccd wire1636/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1647 wire1647/A vssd vccd wire1647/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1658 wire1658/A vssd vccd wire1658/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1669 wire1669/A vssd vccd wire1669/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4046 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input117_A la_data_out_mprj[87] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2034_A wire2034/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3356 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_30 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_401_ _529_/A _401_/B _401_/C vssd vccd _401_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_15_3209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_41 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_63 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_74 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_332_ _332_/A _332_/B vssd vccd _332_/X vssd vccd sky130_fd_sc_hd__and2_4
XPHY_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_4500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2201_A wire2202/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_96 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_263_ _263_/A _263_/B vssd vccd _263_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_6_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input82_A la_data_out_mprj[55] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_194_ _194_/A _194_/B vssd vccd _194_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire966 wire966/A vssd vccd _074_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire977 wire977/A vssd vccd _062_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire988 wire988/A vssd vccd _094_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire999 _556_/X vssd vccd wire999/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output503_A wire1124/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__374__A_N _502_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1301_A wire1302/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output872_A _336_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_17 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[28\] mprj_dat_i_user[28] max_length1310/X vssd vccd _142_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XANTENNA_28 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] _178_/X vssd vccd _162_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XANTENNA_39 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1670_A wire1671/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1768_A wire1768/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4551 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__A _303_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1935_A wire1936/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3999 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] _289_/X vssd vccd wire980/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_0_4244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1698 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2596 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3603 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3647 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4280 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__213__A _213_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4166 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput680 _048_/Y vssd vccd la_data_in_mprj[65] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2101 wire2101/A vssd vccd wire2101/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_27_2979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2112 wire2113/X vssd vccd _480_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput691 _058_/Y vssd vccd la_data_in_mprj[75] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2123 wire2123/A vssd vccd _475_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2134 wire2134/A vssd vccd wire2134/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1400 wire1400/A vssd vccd wire1400/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2145 wire2145/A vssd vccd _458_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1411 wire1411/A vssd vccd wire1411/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2156 wire2157/X vssd vccd _454_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1422 wire1423/X vssd vccd _308_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2167 wire2168/X vssd vccd _450_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input234_A la_iena_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1433 wire1434/X vssd vccd wire1433/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2178 wire2178/A vssd vccd wire2178/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1444 wire1445/X vssd vccd wire1444/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2189 wire2190/X vssd vccd _439_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1455 wire1456/X vssd vccd wire1455/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1466 wire1466/A vssd vccd wire1466/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1477 wire1478/X vssd vccd _326_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__397__A_N _525_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1488 wire1489/X vssd vccd wire1488/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1499 wire1500/X vssd vccd wire1499/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input401_A mprj_adr_o_core[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_315_ _315_/A _315_/B vssd vccd _315_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_246_ _246_/A _246_/B vssd vccd _246_/X vssd vccd sky130_fd_sc_hd__and2_4
Xinput15 la_data_out_mprj[10] vssd vccd _379_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput26 la_data_out_mprj[11] vssd vccd _380_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_4396 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput37 la_data_out_mprj[14] vssd vccd _383_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_32_1951 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput48 la_data_out_mprj[24] vssd vccd _393_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_out_mprj[34] vssd vccd _403_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_45_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_177_ _177_/A _177_/B vssd vccd _177_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_1372 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1084_A _426_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2478 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1251_A wire1252/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1349_A wire1349/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__496__C _496_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_4528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1516_A wire1517/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_482 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1885_A wire1885/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_1283 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire969_A wire969/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__033__A _033_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput408 mprj_adr_o_core[28] vssd vccd wire1451/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_44_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput419 mprj_adr_o_core[9] vssd vccd wire1400/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1451 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__208__A _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_100_ _100_/A vssd vccd _100_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_51_1837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_031_ _031_/A vssd vccd _031_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input184_A la_iena_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2199_A wire2199/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input351_A la_oenb_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input449_A mprj_dat_o_core[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input45_A la_data_out_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__597__B _597_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1230 wire1231/X vssd vccd wire1230/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1241 wire1242/X vssd vccd wire1241/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1252 _337_/X vssd vccd wire1252/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1263 _319_/X vssd vccd wire1263/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1274 wire1275/X vssd vccd wire1274/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1285 wire1286/X vssd vccd wire1285/X vssd vccd sky130_fd_sc_hd__buf_8
Xwire1296 wire1297/X vssd vccd wire1296/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3860 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__118__A _118_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3735 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__A_N _412_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output570_A _450_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_229_ _229_/A _229_/B vssd vccd _229_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_wire1299_A wire1300/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output835_A wire1045/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1466_A wire1466/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] _245_/X vssd vccd _065_/A vssd vccd
+ sky130_fd_sc_hd__nand2_8
XFILLER_44_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3864 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_3875 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__300__B _300_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_3515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1935 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2803 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3668 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1091 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2599 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_3814 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput205 la_iena_mprj[50] vssd vccd _213_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput216 la_iena_mprj[60] vssd vccd _223_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput227 la_iena_mprj[70] vssd vccd _233_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_6_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput238 la_iena_mprj[80] vssd vccd _243_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3363 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput249 la_iena_mprj[90] vssd vccd _253_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__210__B _210_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_580_ _580_/A _580_/B vssd vccd _580_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3003 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_2411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__435__A_N _563_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input399_A mprj_adr_o_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_786 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_014_ _014_/A vssd vccd _014_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_2805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3230 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_687 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1060 _475_/X vssd vccd wire1060/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1071 _464_/X vssd vccd wire1071/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1082 wire1083/X vssd vccd wire1082/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1093 wire1094/X vssd vccd wire1093/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1047_A _503_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2288 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3808 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1214_A wire1215/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output785_A wire1015/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output952_A output952/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[10\] mprj_dat_i_user[10] _294_/X vssd vccd _124_/A vssd vccd sky130_fd_sc_hd__nand2_2
XFILLER_12_3598 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1750_A wire1750/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4384 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3708 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4100 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__458__A_N _586_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_4024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2639 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__205__B _205_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1695 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2064_A wire2065/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input147_A la_iena_mprj[113] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input314_A la_oenb_mprj[33] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_563_ _563_/A _563_/B vssd vccd _563_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_494_ _622_/A _494_/B _494_/C vssd vccd _494_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_38_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2110 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2886 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput509 wire1118/X vssd vccd la_data_in_core[26] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output533_A wire1096/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__131__A _131_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1164_A wire1165/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1331_A _246_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1429_A wire1430/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] _208_/X vssd vccd _028_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_4355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_804 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4486 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1798_A wire1798/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_4096 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__306__A _306_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2650 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1965_A wire1966/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1094 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] _170_/X vssd vccd _154_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_28_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[29\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1807 wire1807/A vssd vccd _245_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1818 wire1818/A vssd vccd _208_/A vssd vccd sky130_fd_sc_hd__buf_4
Xwire1829 wire1829/A vssd vccd _191_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_107 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_118 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_129 _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3262 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_572 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__216__A _216_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2181_A wire2181/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input264_A la_oenb_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input431_A mprj_dat_o_core[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2598 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_300 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_615_ _615_/A _615_/B vssd vccd _615_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_29_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_546_ _546_/A _546_/B vssd vccd _546_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_45_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_477_ _477_/A_N _477_/B _477_/C vssd vccd _477_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_50_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output483_A _487_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__126__A _126_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1223 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output650_A _021_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output748_A _623_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1281_A wire1282/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2454 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1379_A wire1380/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2307 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output915_A wire1220/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_4376 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1713_A wire1713/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire999_A _556_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_678 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_1156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__036__A _036_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_2480 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput840 _591_/X vssd vccd la_oenb_core[94] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput851 wire1266/X vssd vccd mprj_adr_o_user[12] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_2014 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput862 wire1254/X vssd vccd mprj_adr_o_user[22] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput873 _308_/X vssd vccd mprj_adr_o_user[3] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput884 _126_/Y vssd vccd mprj_dat_i_core[12] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_21_3406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput895 _136_/Y vssd vccd mprj_dat_i_core[22] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1335 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1604 _472_/A_N vssd vccd _600_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1615 wire1615/A vssd vccd _186_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1626 wire1626/A vssd vccd _447_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1637 wire1638/X vssd vccd _393_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_24_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1648 wire1649/X vssd vccd _387_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1659 wire1660/X vssd vccd _382_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_400_ _400_/A_N _400_/B _400_/C vssd vccd _400_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_26_152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_20 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_31 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2027_A wire2027/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_64 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_331_ _331_/A _331_/B vssd vccd _331_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_19_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_75 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_86 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_262_ _262_/A _262_/B vssd vccd _262_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_52_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input381_A la_oenb_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_193_ _193_/A _193_/B vssd vccd _193_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_6_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire967 wire967/A vssd vccd _073_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input75_A la_data_out_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire978 wire978/A vssd vccd _061_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire989 wire989/A vssd vccd _093_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3700 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1127_A _386_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_529_ _529_/A _529_/B vssd vccd _529_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_33_2609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_18 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_29 mprj_dat_i_user[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3799 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output865_A _330_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1496_A wire1497/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1031 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1663_A wire1664/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__303__B _303_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3704 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1830_A wire1830/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1928_A wire1929/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] _282_/X vssd vccd _102_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_0_3544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3472 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2591 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3615 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4292 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3659 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4051 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__213__B _213_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_4145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput670 _039_/Y vssd vccd la_data_in_mprj[56] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_27_2958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_4095 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput681 _049_/Y vssd vccd la_data_in_mprj[66] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4178 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2102 wire2103/X vssd vccd _484_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput692 _059_/Y vssd vccd la_data_in_mprj[76] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_21_3203 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2113 wire2114/X vssd vccd wire2113/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2124 wire2125/X vssd vccd _474_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_3394 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2135 wire2135/A vssd vccd _468_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1401 wire1402/X vssd vccd _313_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2146 wire2147/X vssd vccd _457_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1412 wire1413/X vssd vccd _310_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2157 wire2158/X vssd vccd wire2157/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1423 wire1424/X vssd vccd wire1423/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2168 wire2168/A vssd vccd wire2168/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1434 wire1435/X vssd vccd wire1434/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2179 wire2179/A vssd vccd _309_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1445 wire1446/X vssd vccd wire1445/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1456 wire1456/A vssd vccd wire1456/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1467 wire1468/X vssd vccd _329_/B vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_input227_A la_iena_mprj[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1478 wire1479/X vssd vccd wire1478/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1489 wire1489/A vssd vccd wire1489/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_314_ _314_/A _314_/B vssd vccd _314_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_51_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4320 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4364 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_245_ _245_/A _245_/B vssd vccd _245_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput16 la_data_out_mprj[110] vssd vccd _479_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput27 la_data_out_mprj[120] vssd vccd input27/X vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput38 la_data_out_mprj[15] vssd vccd _384_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_6_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput49 la_data_out_mprj[25] vssd vccd _394_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
X_176_ _176_/A _176_/B vssd vccd _176_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1395 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1077_A _458_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1244_A wire1245/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1990 wire1991/X vssd vccd _579_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_450 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3828 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1411_A wire1411/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_494 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__A_N _619_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1509_A wire1510/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_290 _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1780_A wire1781/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1186 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1878_A wire1878/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_1484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4224 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput409 mprj_adr_o_core[29] vssd vccd wire1446/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_1211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_910 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__208__B _208_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_030_ _030_/A vssd vccd _030_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_22_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2247 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__224__A _224_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input177_A la_iena_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2094_A wire2095/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3434 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input344_A la_oenb_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3274 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input38_A la_data_out_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1220 wire1221/X vssd vccd wire1220/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1231 _345_/X vssd vccd wire1231/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1242 wire1243/X vssd vccd wire1242/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1253 _328_/X vssd vccd wire1253/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1264 wire1265/X vssd vccd wire1264/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1275 _314_/X vssd vccd wire1275/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1286 wire1287/X vssd vccd wire1286/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1297 wire1298/X vssd vccd wire1297/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_781 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_228_ _228_/A _228_/B vssd vccd _228_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_7_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_159_ _159_/A vssd vccd _159_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_7_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1194_A wire1195/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output730_A wire1042/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output828_A _580_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1361_A wire1361/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1459_A wire1460/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] _238_/X vssd vccd _058_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_3887 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1626_A wire1626/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4348 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1947 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__A _309_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1995_A wire1995/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2859 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_3371 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__044__A _044_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__387__A_N _515_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3826 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput206 la_iena_mprj[51] vssd vccd _214_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput217 la_iena_mprj[61] vssd vccd _224_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_4087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput228 la_iena_mprj[71] vssd vccd _234_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput239 la_iena_mprj[81] vssd vccd _244_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2107_A wire2107/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_798 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input294_A la_oenb_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1056 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_013_ _013_/A vssd vccd _013_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_29_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input461_A user_irq_ena[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3242 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_2574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_850 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1050 _500_/X vssd vccd wire1050/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1061 _474_/X vssd vccd wire1061/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1072 _463_/X vssd vccd wire1072/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1083 _427_/X vssd vccd wire1083/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1094 _419_/X vssd vccd wire1094/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__129__A _129_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3500 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1207_A _353_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output778_A wire1020/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output945_A wire1294/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1576_A wire1577/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3927 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4435 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3640 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__311__B _311_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_3734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1910_A wire1910/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] _264_/X vssd vccd _084_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_39_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4156 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1608 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3540 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__502__A _502_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2714 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_2747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2057_A wire2057/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__402__A_N _530_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1831 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_526 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_562_ _562_/A _562_/B vssd vccd _562_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_2598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input307_A la_oenb_mprj[27] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_493_ _621_/A _493_/B _493_/C vssd vccd _493_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_44_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_2898 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_202 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_3864 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1203 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output526_A wire1103/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1157_A _366_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1786 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1324_A _253_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_1280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output895_A _136_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_816 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] _201_/X vssd vccd _021_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_53_3655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1693_A wire1693/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__306__B _306_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1860_A wire1860/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1958_A wire1958/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2207 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__322__A _322_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4210 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__425__A_N _553_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1808 wire1808/A vssd vccd _244_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1819 wire1819/A vssd vccd _207_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_6_1241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1127 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_108 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_119 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3274 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2442 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__216__B _216_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_728 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[80\]_B wire1332/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4176 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__A _232_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input257_A la_iena_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2174_A wire2174/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2511 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2408 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input424_A mprj_dat_o_core[12] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3063 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input20_A la_data_out_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_614_ _614_/A _614_/B vssd vccd _614_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_37_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_545_ _545_/A _545_/B vssd vccd _545_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3926 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_476_ _604_/A _476_/B _476_/C vssd vccd _476_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_38_1084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output476_A wire1055/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_1235 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[71\]_B _234_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__448__A_N _576_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output643_A _014_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__142__A _142_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1732 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1274_A wire1275/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1826 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output810_A _564_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1441_A wire1441/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1539_A wire1539/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_4131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1706_A wire1707/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_3572 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_208 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput830 _582_/X vssd vccd la_oenb_core[85] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__052__A _052_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput841 _592_/X vssd vccd la_oenb_core[95] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput852 wire1264/X vssd vccd mprj_adr_o_user[13] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4119 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput863 wire1253/X vssd vccd mprj_adr_o_user[23] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput874 _309_/X vssd vccd mprj_adr_o_user[4] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_4299 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput885 _127_/Y vssd vccd mprj_dat_i_core[13] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput896 _137_/Y vssd vccd mprj_dat_i_core[23] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1605 wire1605/A vssd vccd _599_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1616 wire1616/A vssd vccd _457_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1627 wire1627/A vssd vccd _446_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1638 wire1638/A vssd vccd wire1638/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1649 wire1649/A vssd vccd wire1649/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_6_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3336 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_10 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_32 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_43 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_54 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_65 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_330_ _330_/A _330_/B vssd vccd _330_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_26_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_76 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_87 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_98 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__A _227_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_261_ _261_/A _261_/B vssd vccd _261_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_2370 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_192_ _192_/A _192_/B vssd vccd _192_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_48_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_2289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire968 wire968/A vssd vccd _072_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire979 wire979/A vssd vccd _110_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input374_A la_oenb_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input68_A la_data_out_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3712 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_528_ _528_/A _528_/B vssd vccd _528_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_50_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1022_A wire1023/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output593_A _084_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__137__A _137_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_459_ _587_/A _459_/B _459_/C vssd vccd _459_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_19 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output760_A wire1031/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output858_A wire1257/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1391_A wire1392/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1043 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1087 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1656_A wire1656/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__600__A _600_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1823_A wire1823/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_4196 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__047__A _047_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2690 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[35\]_B _198_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3627 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4063 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput660 _030_/Y vssd vccd la_data_in_mprj[47] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput671 _040_/Y vssd vccd la_data_in_mprj[57] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput682 _050_/Y vssd vccd la_data_in_mprj[67] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2103 wire2104/X vssd vccd wire2103/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput693 _060_/Y vssd vccd la_data_in_mprj[77] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_1111 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2114 wire2114/A vssd vccd wire2114/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2125 wire2125/A vssd vccd wire2125/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__510__A _510_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3215 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire2136 wire2136/A vssd vccd _467_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1402 wire1403/X vssd vccd wire1402/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2147 wire2148/X vssd vccd wire2147/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1413 wire1414/X vssd vccd wire1413/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2158 wire2158/A vssd vccd wire2158/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1424 wire1425/X vssd vccd wire1424/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2169 wire2170/X vssd vccd _449_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1435 wire1436/X vssd vccd wire1435/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1446 wire1446/A vssd vccd wire1446/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1457 wire1458/X vssd vccd _331_/B vssd vccd sky130_fd_sc_hd__buf_8
Xwire1468 wire1469/X vssd vccd wire1468/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1479 wire1480/X vssd vccd wire1479/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input122_A la_data_out_mprj[91] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2137_A wire2138/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2919 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_313_ _313_/A _313_/B vssd vccd _313_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_35_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_244_ _244_/A _244_/B vssd vccd _244_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_10_340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_4376 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput17 la_data_out_mprj[111] vssd vccd _480_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput28 la_data_out_mprj[121] vssd vccd _490_/C vssd vccd sky130_fd_sc_hd__buf_4
Xinput39 la_data_out_mprj[16] vssd vccd _385_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_10_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_175_ _175_/A _175_/B vssd vccd _175_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_6_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[3\] mprj_dat_i_user[3] max_length1311/X vssd vccd _117_/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[110\]_B _273_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output606_A _096_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1980 wire1980/A vssd vccd wire1980/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1991 wire1991/A vssd vccd wire1991/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_462 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1404_A wire1404/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_1831 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_280 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] _183_/X vssd vccd _003_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
XANTENNA_291 _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1773_A wire1774/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[17\]_B _180_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__314__B _314_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1940_A wire1940/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__330__A _330_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_3607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3568 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1278 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2580 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_A mprj_dat_i_user[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__505__A _505_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3446 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2087_A wire2087/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2035 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__A _240_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput490 _493_/X vssd vccd la_data_in_core[124] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3286 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input337_A la_oenb_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1210 _352_/X vssd vccd wire1210/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1221 wire1222/X vssd vccd wire1221/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1232 wire1233/X vssd vccd wire1232/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1243 _341_/X vssd vccd wire1243/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1254 wire1255/X vssd vccd wire1254/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1265 _318_/X vssd vccd wire1265/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1276 _313_/X vssd vccd wire1276/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1287 wire1288/X vssd vccd wire1287/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1298 _301_/X vssd vccd wire1298/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4162 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_227_ _227_/A _227_/B vssd vccd _227_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_45_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1160 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_158_ _158_/A vssd vccd _158_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_13_1171 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output556_A _438_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_089_ _089_/A vssd vccd _089_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_wire1187_A wire1188/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output723_A _600_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1354_A wire1355/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3899 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] _231_/X vssd vccd _051_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_22_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1521_A wire1521/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1619_A wire1619/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3615 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_292 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4040 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__309__B _309_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1890_A wire1891/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_958 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1988_A wire1989/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire974_A wire974/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3859 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3619 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4191 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__060__A _060_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput207 la_iena_mprj[52] vssd vccd _215_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput218 la_iena_mprj[62] vssd vccd _225_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_41_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput229 la_iena_mprj[72] vssd vccd _235_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_25_1020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1283 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2631 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2747 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2435 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_958 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2002_A wire2002/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__235__A _235_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input287_A la_oenb_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2034 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1068 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_012_ _012_/A vssd vccd _012_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_4_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1311 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input454_A mprj_sel_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input50_A la_data_out_mprj[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__481__A_N _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__401__C _401_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1040 _509_/X vssd vccd wire1040/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1051 _499_/X vssd vccd wire1051/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1062 _473_/X vssd vccd wire1062/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1073 _462_/X vssd vccd wire1073/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1084 _426_/X vssd vccd wire1084/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1095 _418_/X vssd vccd wire1095/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_3913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3826 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3534 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1102_A _411_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3556 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__145__A _145_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1299 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output840_A _591_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output938_A wire1244/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1471_A wire1471/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3939 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4447 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1736_A wire1737/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1226 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1903_A wire1904/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_4168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__055__A _055_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_2977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_604 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2840 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__502__B _502_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3668 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_561_ _561_/A _561_/B vssd vccd _561_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_1854 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input202_A la_iena_mprj[48] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_492_ _620_/A _492_/B _492_/C vssd vccd _492_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_44_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1411 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input98_A la_data_out_mprj[6] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3338 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__B _412_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3983 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output519_A wire1109/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4400 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1052_A _498_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__377__A_N _505_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3754 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output790_A wire1011/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_828 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_1339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1686_A wire1687/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__603__A _603_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1853_A wire1853/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_3703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__322__B _322_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_2219 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3736 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4222 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[2\]_A mprj_dat_i_user[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1809 wire1809/A vssd vccd _335_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_4288 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2820 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3598 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_109 mprj_dat_i_user[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_3144 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3286 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4111 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__A _513_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4144 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4188 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__232__B _232_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3307 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input152_A la_iena_mprj[118] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2167_A wire2168/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3075 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input417_A mprj_adr_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_613_ _613_/A _613_/B vssd vccd _613_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input13_A la_data_out_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_544_ _544_/A _544_/B vssd vccd _544_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_44_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_475_ _603_/A _475_/B _475_/C vssd vccd _475_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__407__B _407_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3640 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3684 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output469_A wire1061/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output636_A _008_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output803_A wire997/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1434_A wire1435/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_600 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput390 mprj_adr_o_core[11] vssd vccd wire1519/A vssd vccd sky130_fd_sc_hd__buf_6
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] _213_/X vssd vccd _033_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_53_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4116 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3551 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_636 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1183 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__317__B _317_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4474 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1027 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1970_A wire1970/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1336 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__A _333_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput820 _573_/X vssd vccd la_oenb_core[76] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput831 _583_/X vssd vccd la_oenb_core[86] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput842 _593_/X vssd vccd la_oenb_core[96] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput853 wire1262/X vssd vccd mprj_adr_o_user[14] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput864 _329_/X vssd vccd mprj_adr_o_user[24] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput875 _310_/X vssd vccd mprj_adr_o_user[5] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput886 _128_/Y vssd vccd mprj_dat_i_core[14] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput897 _138_/Y vssd vccd mprj_dat_i_core[24] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1606 wire1606/A vssd vccd _598_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input5_A la_data_out_mprj[100] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1617 wire1617/A vssd vccd _456_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2887 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1628 wire1628/A vssd vccd _445_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1639 wire1640/X vssd vccd _392_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_11 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_33 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_44 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__508__A _508_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_55 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_66 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_88 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_99 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__227__B _227_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3094 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_260_ _260_/A _260_/B vssd vccd _260_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_23_872 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_883 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_191_ _191_/A _191_/B vssd vccd _191_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire969 wire969/A vssd vccd _071_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__243__A _243_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input367_A la_oenb_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_irq_gates\[2\] user_irq_core[2] _293_/X vssd vccd _113_/A vssd vccd sky130_fd_sc_hd__nand2_1
XFILLER_43_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3262 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_231 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3920 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_527_ _527_/A _527_/B vssd vccd _527_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_15_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_458_ _586_/A _458_/B _458_/C vssd vccd _458_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__415__A_N _415_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output586_A wire1070/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_389_ _517_/A _389_/B _389_/C vssd vccd _389_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_12_1011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output753_A wire1037/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1055 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1099 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output920_A wire1205/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] _261_/X vssd vccd _081_/A vssd vccd
+ sky130_fd_sc_hd__nand2_8
XFILLER_29_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1649_A wire1649/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__600__B _600_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1816_A wire1816/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4060 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1209 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__063__A _063_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3639 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4031 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4075 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput650 _021_/Y vssd vccd la_data_in_mprj[38] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput661 _031_/Y vssd vccd la_data_in_mprj[48] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput672 _041_/Y vssd vccd la_data_in_mprj[58] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput683 _051_/Y vssd vccd la_data_in_mprj[68] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2104 wire2104/A vssd vccd wire2104/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2115 wire2116/X vssd vccd _479_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput694 _061_/Y vssd vccd la_data_in_mprj[78] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_1123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2126 wire2127/X vssd vccd _473_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__510__B _510_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_2651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2137 wire2138/X vssd vccd _466_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1403 wire1404/X vssd vccd wire1403/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2148 wire2148/A vssd vccd wire2148/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1167 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1414 wire1415/X vssd vccd wire1414/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2159 wire2160/X vssd vccd _453_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1425 wire1426/X vssd vccd wire1425/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1436 wire1436/A vssd vccd wire1436/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1447 wire1448/X vssd vccd _333_/B vssd vccd sky130_fd_sc_hd__buf_8
Xwire1458 wire1459/X vssd vccd wire1458/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1469 wire1470/X vssd vccd wire1469/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2032_A wire2032/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input115_A la_data_out_mprj[85] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__438__A_N _566_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__238__A _238_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_312_ _312_/A _312_/B vssd vccd _312_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_51_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_2488 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_243_ _243_/A _243_/B vssd vccd _243_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput18 la_data_out_mprj[112] vssd vccd _481_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_input80_A la_data_out_mprj[53] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput29 la_data_out_mprj[122] vssd vccd _491_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
X_174_ _174_/A _174_/B vssd vccd _174_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_6_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__404__C _404_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__420__B _420_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1690 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1970 wire1970/A vssd vccd wire1970/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output501_A wire1125/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1981 wire1982/X vssd vccd _583_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_1335 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1992 wire1993/X vssd vccd _578_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_15_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3808 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1132_A _381_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_4380 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_270 _215_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_281 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_292 wire1707/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] _176_/X vssd vccd _160_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_33_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_wb_dat_gates\[26\] mprj_dat_i_user[26] _294_/X vssd vccd _140_/A vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_53_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1599_A _477_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1766_A wire1766/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4204 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__611__A _611_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1443 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__330__B _330_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] wire1312/X vssd vccd _107_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_42_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2620 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__058__A _058_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[10\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__505__B _505_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1559 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__521__A _521_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput480 _484_/X vssd vccd la_data_in_core[115] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput491 _494_/X vssd vccd la_data_in_core[125] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__240__B _240_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2047 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1200 wire1201/X vssd vccd wire1200/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1211 wire1212/X vssd vccd wire1211/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1222 _348_/X vssd vccd wire1222/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1233 wire1234/X vssd vccd wire1233/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input232_A la_iena_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_2323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1244 wire1245/X vssd vccd wire1244/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1255 _327_/X vssd vccd wire1255/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1266 wire1267/X vssd vccd wire1266/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1277 _312_/X vssd vccd wire1277/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1288 _303_/X vssd vccd wire1288/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1299 wire1300/X vssd vccd wire1299/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_38_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_411 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_915 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3896 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3787 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_226_ _226_/A _226_/B vssd vccd _226_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA__415__B _415_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_4196 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_157_ _157_/A vssd vccd _157_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_6_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1183 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_088_ _088_/A vssd vccd _088_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output549_A wire1078/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1082_A wire1083/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_392 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output716_A _081_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4375 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1347_A wire1347/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4052 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3204 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__606__A _606_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1883_A wire1884/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__325__B _325_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire967_A wire967/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2558 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__341__A _341_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_819 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4264 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4034 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_318 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3300 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput208 la_iena_mprj[53] vssd vccd _216_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput219 la_iena_mprj[63] vssd vccd _226_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1251 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1295 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__516__A _516_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__235__B _235_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_011_ _011_/A vssd vccd _011_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_46_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input182_A la_iena_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1323 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2197_A wire2197/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__251__A _251_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3266 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input447_A mprj_dat_o_core[4] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input43_A la_data_out_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3062 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1030 _519_/X vssd vccd wire1030/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1041 _508_/X vssd vccd wire1041/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_856 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2383 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1052 _498_/X vssd vccd wire1052/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1063 _472_/X vssd vccd wire1063/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1074 _461_/X vssd vccd wire1074/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1085 wire1086/X vssd vccd wire1085/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2247 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1096 _417_/X vssd vccd wire1096/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output499_A wire1127/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_3693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_209_ _209_/A _209_/B vssd vccd _209_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_32_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1297_A wire1298/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output833_A _585_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__161__A _161_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1464_A wire1465/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_3620 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] wire1332/X vssd vccd wire976/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_3_4459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3664 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1806 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1631_A wire1631/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1729_A wire1730/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_1902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__336__A _336_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3603 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3636 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__071__A _071_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1070 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_560_ _560_/A _560_/B vssd vccd _560_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_45_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1866 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_491_ _619_/A _491_/B _491_/C vssd vccd _491_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_39_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2812 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2112_A wire2113/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__246__A _246_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3844 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1423 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input397_A mprj_adr_o_core[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__412__C _412_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4470 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_682 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4412 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1045_A _505_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1332 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_550 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3766 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1212_A wire1213/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output783_A wire1016/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__156__A _156_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output950_A wire1299/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1679_A wire1679/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__603__B _603_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_4201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1846_A wire1846/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3759 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[2\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3472 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_3544 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2832 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_2876 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__471__A_N _599_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3118 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__066__A _066_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_2428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2753 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__513__B _513_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1451 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_903 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3444 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3372 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2062_A wire2063/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input145_A la_iena_mprj[111] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_612_ _612_/A _612_/B vssd vccd _612_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_input312_A la_oenb_mprj[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1630 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_543_ _543_/A _543_/B vssd vccd _543_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_50_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_474_ _602_/A _474_/B _474_/C vssd vccd _474_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_4320 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__423__B _423_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4471 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output531_A wire1098/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1162_A wire1163/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput380 la_oenb_mprj[93] vssd vccd _590_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput391 mprj_adr_o_core[12] vssd vccd wire1517/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1427_A wire1428/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__494__A_N _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] _206_/X vssd vccd _026_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_18_3530 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_1090 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_648 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3416 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3487 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__614__A _614_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1963_A wire1964/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1348 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__333__B _333_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3720 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput810 _564_/X vssd vccd la_oenb_core[67] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput821 _574_/X vssd vccd la_oenb_core[77] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput832 _584_/X vssd vccd la_oenb_core[87] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput843 _594_/X vssd vccd la_oenb_core[97] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3764 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput854 wire1261/X vssd vccd mprj_adr_o_user[15] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput865 _330_/X vssd vccd mprj_adr_o_user[25] vssd vccd sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] _168_/X vssd vccd _152_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
Xoutput876 wire1278/X vssd vccd mprj_adr_o_user[6] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_3_4020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput887 _129_/Y vssd vccd mprj_dat_i_core[15] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput898 _139_/Y vssd vccd mprj_dat_i_core[25] vssd vccd sky130_fd_sc_hd__buf_8
Xwire1607 wire1607/A vssd vccd _597_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1618 wire1618/A vssd vccd _455_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_3352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1629 wire1629/A vssd vccd _444_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_2189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_12 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_34 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_56 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__B _508_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_67 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_78 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3972 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_190_ _190_/A _190_/B vssd vccd _190_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_22_394 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__524__A _524_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_3869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__243__B _243_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1860 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input262_A la_oenb_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_711 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3932 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3976 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2398 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__418__B _418_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_526_ _526_/A _526_/B vssd vccd _526_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_50_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2049 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_457_ _585_/A _457_/B _457_/C vssd vccd _457_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_53_1326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_388_ _516_/A _388_/B _388_/C vssd vccd _388_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output481_A _485_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output579_A wire1137/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_48_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1067 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output746_A _621_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1377_A wire1377/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3843 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output913_A wire1251/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1544_A wire1544/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4215 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1428 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1711_A wire1711/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1809_A wire1809/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__609__A _609_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_2857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__328__B _328_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire997_A wire998/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2523 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2567 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__344__A _344_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_10_2409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput640 _012_/Y vssd vccd la_data_in_mprj[29] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3403 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput651 _022_/Y vssd vccd la_data_in_mprj[39] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_4087 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput662 _032_/Y vssd vccd la_data_in_mprj[49] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput673 _042_/Y vssd vccd la_data_in_mprj[59] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput684 _052_/Y vssd vccd la_data_in_mprj[69] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2105 wire2106/X vssd vccd _483_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput695 _062_/Y vssd vccd la_data_in_mprj[79] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2116 wire2116/A vssd vccd wire2116/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2127 wire2127/A vssd vccd wire2127/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2138 wire2138/A vssd vccd wire2138/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1404 wire1404/A vssd vccd wire1404/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2149 wire2150/X vssd vccd _456_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1415 wire1416/X vssd vccd wire1415/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1426 wire1426/A vssd vccd wire1426/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_8_1179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1437 wire1438/X vssd vccd _307_/B vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1448 wire1449/X vssd vccd wire1448/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1459 wire1460/X vssd vccd wire1459/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__519__A _519_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__238__B _238_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input108_A la_data_out_mprj[79] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_311_ _311_/A _311_/B vssd vccd _311_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_242_ _242_/A _242_/B vssd vccd _242_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_52_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_180 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__254__A _254_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput19 la_data_out_mprj[113] vssd vccd _482_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_173_ _173_/A _173_/B vssd vccd _173_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_49_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input73_A la_data_out_mprj[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__420__C _420_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1960 wire1961/X vssd vccd wire1960/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1971 wire1971/A vssd vccd _590_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1982 wire1983/X vssd vccd wire1982/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1993 wire1993/A vssd vccd wire1993/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1125_A _388_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_260 _470_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_271 _216_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_282 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_509_ _509_/A _509_/B vssd vccd _509_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_37_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_293 wire1754/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_106 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output863_A wire1253/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__164__A _164_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[19\] mprj_dat_i_user[19] max_length1311/X vssd vccd _133_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XANTENNA_wire1494_A wire1495/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1498 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1661_A wire1662/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1759_A wire1760/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3712 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__611__B _611_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1926_A wire1927/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_1477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] _280_/X vssd vccd wire983/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_37_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2022 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_489 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__074__A _074_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_3986 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__521__B _521_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput470 wire1060/X vssd vccd la_data_in_core[106] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput481 _485_/X vssd vccd la_data_in_core[116] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput492 _495_/X vssd vccd la_data_in_core[126] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_40_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2059 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__405__A_N _405_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1201 _355_/X vssd vccd wire1201/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1212 wire1213/X vssd vccd wire1212/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1223 wire1224/X vssd vccd wire1223/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1234 _344_/X vssd vccd wire1234/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1245 _340_/X vssd vccd wire1245/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1256 _325_/X vssd vccd wire1256/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2142_A wire2142/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input225_A la_iena_mprj[69] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1267 _317_/X vssd vccd wire1267/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1278 wire1279/X vssd vccd wire1278/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1289 wire1290/X vssd vccd wire1289/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_34_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__249__A _249_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_979 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3886 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_225_ _225_/A _225_/B vssd vccd _225_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_11_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__415__C _415_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_156_ _156_/A vssd vccd _156_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1195 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_087_ _087_/A vssd vccd _087_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_49_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4503 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__B _431_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2279 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1075_A _460_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output611_A _101_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output709_A _074_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1242_A wire1243/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_2930 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1790 wire1790/A vssd vccd wire1790/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_795 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1507_A wire1508/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4064 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__606__B _606_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1876_A wire1877/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__622__A _622_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__341__B _341_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__428__A_N _556_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4171 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4046 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput209 la_iena_mprj[54] vssd vccd _217_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_3406 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__069__A _069_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_710 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__516__B _516_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_010_ _010_/A vssd vccd _010_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_10_2058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__532__A _532_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1335 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2092_A wire2093/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input175_A la_iena_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3278 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input342_A la_oenb_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input36_A la_data_out_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1020 wire1021/X vssd vccd wire1020/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1031 _518_/X vssd vccd wire1031/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2204 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1042 wire1043/X vssd vccd wire1042/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1053 _497_/X vssd vccd wire1053/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2395 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1064 _471_/X vssd vccd wire1064/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1075 _460_/X vssd vccd wire1075/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1086 _425_/X vssd vccd wire1086/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1097 _416_/X vssd vccd wire1097/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4340 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4362 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_208_ _208_/A _208_/B vssd vccd _208_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_45_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_975 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output561_A _442_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output659_A _029_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_139_ _139_/A vssd vccd _139_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1192_A wire1193/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output826_A _578_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3790 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3632 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1457_A wire1458/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3676 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] _236_/X vssd vccd _056_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_26_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1624_A wire1624/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3450 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__617__A _617_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1993_A wire1993/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_746 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__336__B _336_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1947 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2924 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[92\]_B wire1322/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_1611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__352__A _352_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3648 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1082 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_490_ _618_/A _490_/B _490_/C vssd vccd _490_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__527__A _527_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3823 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2105_A wire2106/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_3856 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_267 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1435 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input292_A la_oenb_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[83\]_B wire1331/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__262__A _262_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2065 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3042 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xmax_length1562 _416_/A_N vssd vccd wire1561/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_4482 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1038_A _511_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_562 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1205_A wire1206/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output776_A _533_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1791 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[74\]_B _237_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output943_A wire1229/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__172__A _172_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4406 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_4393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1741_A wire1741/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4246 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1839_A wire1839/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_4279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1058 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2888 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_3233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__347__A _347_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_3878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_554 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2587 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__082__A _082_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_436 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2310 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input138_A la_iena_mprj[105] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire2055_A wire2056/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_611_ _611_/A _611_/B vssd vccd _611_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_29_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1642 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_542_ _542_/A _542_/B vssd vccd _542_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_input305_A la_oenb_mprj[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__257__A _257_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_473_ _601_/A _473_/B _473_/C vssd vccd _473_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_44_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__423__C _423_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3810 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3771 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output524_A wire1142/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3854 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1155_A wire1156/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput370 la_oenb_mprj[84] vssd vccd wire1533/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput381 la_oenb_mprj[94] vssd vccd _591_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_7_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput392 mprj_adr_o_core[13] vssd vccd wire1514/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1322_A _255_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__167__A _167_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] _199_/X vssd vccd _019_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_1196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3428 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_2787 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1691_A wire1691/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3152 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1789_A wire1790/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__614__B _614_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_4203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1956_A wire1956/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput800 wire1000/X vssd vccd la_oenb_core[58] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput811 _565_/X vssd vccd la_oenb_core[68] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3732 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput822 _575_/X vssd vccd la_oenb_core[78] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput833 _585_/X vssd vccd la_oenb_core[88] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput844 _595_/X vssd vccd la_oenb_core[98] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput855 wire1260/X vssd vccd mprj_adr_o_user[16] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1201 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3776 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput866 _331_/X vssd vccd mprj_adr_o_user[26] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput877 wire1277/X vssd vccd mprj_adr_o_user[7] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput888 _130_/Y vssd vccd mprj_dat_i_core[16] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput899 _140_/Y vssd vccd mprj_dat_i_core[26] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_2834 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1608 input25/X vssd vccd _488_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1619 wire1619/A vssd vccd _454_/C vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_3317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_13 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XPHY_24 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__077__A _077_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_35 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_46 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_68 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_79 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3984 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_B _201_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_2259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__524__B _524_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[122\]_B _285_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_1585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__540__A _540_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_734 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2172_A wire2172/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input255_A la_iena_mprj[96] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3900 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3944 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input422_A mprj_dat_o_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[31\]_A mprj_dat_i_user[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_525_ _525_/A _525_/B vssd vccd _525_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__C _418_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_456_ _584_/A _456_/B _456_/C vssd vccd _456_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_3016 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_387_ _515_/A _387_/B _387_/C vssd vccd _387_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[29\]_B _192_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__434__B _434_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[113\]_B _276_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output474_A wire1135/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output739_A _615_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3855 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1272_A wire1273/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__A_N _589_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3899 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1537_A wire1537/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__609__B _609_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1704_A wire1705/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[22\]_A mprj_dat_i_user[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4084 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__625__A _625_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__344__B _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[104\]_B _267_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_2579 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1282 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2871 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3540 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2907 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput630 _148_/Y vssd vccd la_data_in_mprj[1] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__360__A _360_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput641 _149_/Y vssd vccd la_data_in_mprj[2] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput652 _150_/Y vssd vccd la_data_in_mprj[3] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput663 _151_/Y vssd vccd la_data_in_mprj[4] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput674 _152_/Y vssd vccd la_data_in_mprj[5] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput685 _153_/Y vssd vccd la_data_in_mprj[6] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2106 wire2107/X vssd vccd wire2106/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput696 _154_/Y vssd vccd la_data_in_mprj[7] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2117 wire2118/X vssd vccd _478_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire2128 wire2129/X vssd vccd _472_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire2139 wire2139/A vssd vccd _465_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1405 wire1406/X vssd vccd _312_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1416 wire1416/A vssd vccd wire1416/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1427 wire1428/X vssd vccd _336_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1438 wire1439/X vssd vccd wire1438/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1449 wire1450/X vssd vccd wire1449/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_39_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__519__B _519_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_wb_dat_gates\[13\]_A mprj_dat_i_user[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_3904 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_310_ _310_/A _310_/B vssd vccd _310_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_42_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2018_A wire2018/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__535__A _535_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_241_ _241_/A _241_/B vssd vccd _241_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_51_991 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_1057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_3612 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1300 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__254__B _254_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_172_ _172_/A _172_/B vssd vccd _172_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_49_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input372_A la_oenb_mprj[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__484__A_N _612_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input66_A la_data_out_mprj[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__270__A _270_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3752 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_911 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1950 wire1951/X vssd vccd _598_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1961 wire1962/X vssd vccd wire1961/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1972 wire1972/A vssd vccd _589_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1983 wire1983/A vssd vccd wire1983/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1994 wire1995/X vssd vccd _577_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1291 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_250 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_261 _469_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_508_ _508_/A _508_/B vssd vccd _508_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_272 wire1667/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1020_A wire1021/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_283 _352_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1118_A _395_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_294 wire1756/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output689_A _056_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_118 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_439_ _567_/A _439_/B _439_/C vssd vccd _439_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_31_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output856_A wire1258/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1487_A wire1488/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_892 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__180__A _180_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_4375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4228 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1654_A wire1654/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1248 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1919_A wire1920/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__339__B _339_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__355__A _355_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2387 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3998 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__090__A _090_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput471 wire1059/X vssd vccd la_data_in_core[107] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput482 _486_/X vssd vccd la_data_in_core[117] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput493 _496_/X vssd vccd la_data_in_core[127] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1202 wire1203/X vssd vccd wire1202/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1213 _351_/X vssd vccd wire1213/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1224 wire1225/X vssd vccd wire1224/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1235 wire1236/X vssd vccd wire1235/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1246 wire1247/X vssd vccd wire1246/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1257 _324_/X vssd vccd wire1257/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1268 wire1269/X vssd vccd wire1268/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1279 _311_/X vssd vccd wire1279/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_1718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input120_A la_data_out_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2135_A wire2135/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input218_A la_iena_mprj[62] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_796 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4544 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4408 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2877 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_479 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__265__A _265_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_2287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_224_ _224_/A _224_/B vssd vccd _224_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_7_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_155_ _155_/A vssd vccd _155_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_6_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_wb_dat_gates\[1\] mprj_dat_i_user[1] max_length1310/X vssd vccd _115_/A vssd
+ vccd sky130_fd_sc_hd__nand2_1
XFILLER_6_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_086_ _086_/A vssd vccd _086_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_23_4515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__C _431_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3983 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1068_A _467_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_3665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output604_A _094_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1780 wire1781/X vssd vccd _268_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1235_A wire1236/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1791 wire1792/X vssd vccd _262_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2986 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4032 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1402_A wire1403/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1642 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__175__A _175_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_wb_dat_gates\[31\] mprj_dat_i_user[31] max_length1310/X vssd vccd _145_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_37_1664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1815 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1771_A wire1772/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1869_A wire1870/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__622__B _622_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_2820 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1275 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__085__A _085_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2730 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2085_A wire2086/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input168_A la_iena_mprj[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input335_A la_oenb_mprj[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1010 _547_/X vssd vccd wire1010/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1021 _535_/X vssd vccd wire1021/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1032 _517_/X vssd vccd wire1032/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1043 _507_/X vssd vccd wire1043/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input29_A la_data_out_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1054 _481_/X vssd vccd wire1054/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1065 _470_/X vssd vccd wire1065/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1076 _459_/X vssd vccd wire1076/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1087 wire1088/X vssd vccd wire1087/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1098 _415_/X vssd vccd wire1098/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_3927 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__426__C _426_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3575 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_207_ _207_/A _207_/B vssd vccd _207_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_50_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_138_ _138_/A vssd vccd _138_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA__442__B _442_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output554_A _436_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_069_ _069_/A vssd vccd _069_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output721_A _598_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output819_A _572_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1352_A wire1353/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] _229_/X vssd vccd _049_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_39_3117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3484 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1617_A wire1617/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_593 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__617__B _617_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_2173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1986_A wire1987/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3172 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire972_A wire972/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__352__B _352_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[5\]_A mprj_dat_i_user[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_1107 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1050 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_3176 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1094 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_596 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__543__A _543_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input285_A la_oenb_mprj[122] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__262__B _262_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1111 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1155 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input452_A mprj_dat_o_core[9] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3076 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3087 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3806 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4494 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4327 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3724 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__B _437_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_574 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__418__A_N _546_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1100_A _413_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output769_A wire1051/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_4418 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output936_A wire1150/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1567_A _406_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3452 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1734_A wire1734/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3496 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1901_A wire1901/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_1109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_828 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__347__B _347_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1723 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_2419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__A _363_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_3227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_610_ _610_/A _610_/B vssd vccd _610_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_2_2355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_4013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2048_A wire2048/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_4193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__A _538_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_541_ _541_/A _541_/B vssd vccd _541_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_17_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2319 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input200_A la_iena_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__257__B _257_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_472_ _472_/A_N _472_/B _472_/C vssd vccd _472_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_17_4480 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4371 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input96_A la_data_out_mprj[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__273__A _273_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3866 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output517_A wire1111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput360 la_oenb_mprj[75] vssd vccd wire1542/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_42_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput371 la_oenb_mprj[85] vssd vccd wire1532/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_23_1357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput382 la_oenb_mprj[95] vssd vccd _592_/A vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1050_A _500_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1148_A wire1149/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput393 mprj_adr_o_core[14] vssd vccd wire1511/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_36_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_4255 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4108 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] _192_/X vssd vccd _012_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XANTENNA__390__A_N _518_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__183__A _183_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3186 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1684_A wire1685/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput801 wire999/X vssd vccd la_oenb_core[59] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput812 _566_/X vssd vccd la_oenb_core[69] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1851_A wire1851/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput823 _576_/X vssd vccd la_oenb_core[79] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1949_A wire1949/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3744 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput834 wire995/X vssd vccd la_oenb_core[89] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput845 _596_/X vssd vccd la_oenb_core[99] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_8_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput856 wire1258/X vssd vccd mprj_adr_o_user[17] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput867 _332_/X vssd vccd mprj_adr_o_user[27] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput878 wire1276/X vssd vccd mprj_adr_o_user[8] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput889 _131_/Y vssd vccd mprj_dat_i_core[17] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_3_4033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1257 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_4077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_3260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1609 wire1609/A vssd vccd _231_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_41_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_4008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__358__A _358_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_647 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_14 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_25 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_47 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_69 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3930 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2839 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__093__A _093_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_3996 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3232 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1283 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_768 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input150_A la_iena_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3912 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2165_A wire2166/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input248_A la_iena_mprj[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3956 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input415_A mprj_adr_o_core[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input11_A la_data_out_mprj[106] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_2163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__268__A _268_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[31\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_524_ _524_/A _524_/B vssd vccd _524_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_33_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_455_ _583_/A _455_/B _455_/C vssd vccd _455_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_53_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_386_ _514_/A _386_/B _386_/C vssd vccd _386_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_13_4196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3484 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__434__C _434_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_1096 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output467_A wire1063/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1098_A _415_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__450__B _450_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output634_A _006_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3867 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3709 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1265_A _318_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2052 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4156 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output801_A wire999/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3516 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1432_A wire1433/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1154 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput190 la_iena_mprj[37] vssd vccd _200_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_37_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__178__A _178_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_967 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[22\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_2205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4096 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1899_A wire1900/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_2563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_2536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_2547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1294 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2883 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput620 _109_/Y vssd vccd la_data_in_mprj[126] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput631 _003_/Y vssd vccd la_data_in_mprj[20] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3552 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__360__B _360_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput642 _013_/Y vssd vccd la_data_in_mprj[30] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_43_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput653 _023_/Y vssd vccd la_data_in_mprj[40] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput664 _033_/Y vssd vccd la_data_in_mprj[50] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput675 _043_/Y vssd vccd la_data_in_mprj[60] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput686 _053_/Y vssd vccd la_data_in_mprj[70] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2107 wire2107/A vssd vccd wire2107/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput697 _063_/Y vssd vccd la_data_in_mprj[80] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2118 wire2118/A vssd vccd wire2118/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2129 wire2129/A vssd vccd wire2129/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input3_A caravel_rstn vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1406 wire1407/X vssd vccd wire1406/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1417 wire1418/X vssd vccd _309_/B vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_2518 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1428 wire1429/X vssd vccd wire1428/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1439 wire1440/X vssd vccd wire1439/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3705 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__088__A _088_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_606 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[13\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_240_ _240_/A _240_/B vssd vccd _240_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA__535__B _535_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_171_ _171_/A _171_/B vssd vccd _171_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_3624 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1312 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3646 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input198_A la_iena_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3668 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__A _551_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input365_A la_oenb_mprj[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_510 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_irq_gates\[0\] user_irq_core[0] _291_/X vssd vccd _111_/A vssd vccd sky130_fd_sc_hd__nand2_1
XANTENNA_input59_A la_data_out_mprj[34] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3095 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3764 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1524 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1940 wire1940/A vssd vccd wire1940/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1951 wire1952/X vssd vccd wire1951/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1962 wire1962/A vssd vccd wire1962/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1973 wire1974/X vssd vccd _588_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1984 wire1985/X vssd vccd _582_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__429__C _429_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1995 wire1995/A vssd vccd wire1995/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_967 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_240 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_4236 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_251 _539_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_262 wire2134/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_507_ _507_/A _507_/B vssd vccd _507_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_37_2569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_273 wire1645/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_284 _351_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_295 _270_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__445__B _445_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1013_A wire1014/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_438_ _566_/A _438_/B _438_/C vssd vccd _438_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_output584_A wire1072/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_369_ _497_/A _369_/B _369_/C vssd vccd _369_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_18_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_175 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output751_A wire1039/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output849_A wire1271/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] wire1318/X vssd vccd _079_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_26_4387 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1647_A wire1647/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_4047 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_904 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_2013 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2300 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__355__B _355_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3900 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_2399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_4107 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_697 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_2153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput472 wire1058/X vssd vccd la_data_in_core[108] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput483 _487_/X vssd vccd la_data_in_core[118] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput494 wire1132/X vssd vccd la_data_in_core[12] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2451 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1203 wire1204/X vssd vccd wire1203/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1214 wire1215/X vssd vccd wire1214/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1225 _347_/X vssd vccd wire1225/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1236 wire1237/X vssd vccd wire1236/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1247 wire1248/X vssd vccd wire1247/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1258 wire1259/X vssd vccd wire1258/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1269 wire1270/X vssd vccd wire1269/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_252 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2030_A wire2030/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input113_A la_data_out_mprj[83] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2128_A wire2129/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4556 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__546__A _546_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_2266 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__265__B _265_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__451__A_N _579_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_1407 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_223_ _223_/A _223_/B vssd vccd _223_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_154_ _154_/A vssd vccd _154_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_13_1120 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__281__A _281_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_085_ _085_/A vssd vccd _085_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_3951 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3995 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3622 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1770 wire1770/A vssd vccd wire1770/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1781 wire1781/A vssd vccd wire1781/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1792 wire1792/A vssd vccd wire1792/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1130_A _383_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_1179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1228_A _346_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output799_A _554_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4088 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] _174_/X vssd vccd _158_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_15_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[24\] mprj_dat_i_user[24] _294_/X vssd vccd _138_/A vssd vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1597_A _478_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_4438 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__191__A _191_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1764_A wire1764/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1931_A wire1932/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] _285_/X vssd vccd wire982/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_6_2876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2646 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_3165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__474__A_N _602_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__366__A _366_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1774 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2629 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2078_A wire2078/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1000 wire1001/X vssd vccd wire1000/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1011 wire1012/X vssd vccd wire1011/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1022 wire1023/X vssd vccd wire1022/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input230_A la_iena_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1033 _516_/X vssd vccd wire1033/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input328_A la_oenb_mprj[46] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3892 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1044 _506_/X vssd vccd wire1044/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1055 _480_/X vssd vccd wire1055/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1066 _469_/X vssd vccd wire1066/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1077 _458_/X vssd vccd wire1077/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1088 _424_/X vssd vccd wire1088/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1099 _414_/X vssd vccd wire1099/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__276__A _276_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_206_ _206_/A _206_/B vssd vccd _206_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_3284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_137_ _137_/A vssd vccd _137_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_8_999 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2550 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__442__C _442_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_068_ _068_/A vssd vccd _068_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output547_A wire1080/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1080_A _429_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1178_A wire1179/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output714_A _079_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_4131 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1345_A wire1345/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1388 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] _222_/X vssd vccd _042_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_1_2740 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1512_A wire1513/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_3416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1716 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__A _186_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_4453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2450 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1881_A wire1882/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1979_A wire1980/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3512 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[5\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4042 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3188 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1825 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__096__A _096_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4504 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2258 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__543__B _543_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2594 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input180_A la_iena_mprj[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2195_A wire2195/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input278_A la_oenb_mprj[116] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_3105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1167 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3066 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_3149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input445_A mprj_dat_o_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_3099 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input41_A la_data_out_mprj[18] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_1493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_1274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_3736 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3627 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__437__C _437_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output497_A wire1129/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__B _453_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2667 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1295_A wire1296/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output831_A _583_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_4121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output929_A wire1174/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1462_A wire1463/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1439 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1727_A wire1728/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3282 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_380 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_512 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_545 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__363__B _363_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2767 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3425 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3458 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1984 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_3035 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1791 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__538__B _538_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_540_ _540_/A _540_/B vssd vccd _540_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_4069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_471_ _599_/A _471_/B _471_/C vssd vccd _471_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_32_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4312 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4492 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2110_A wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2208_A wire2209/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A _554_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input395_A mprj_adr_o_core[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__273__B _273_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input89_A la_data_out_mprj[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_3128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_4305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_961 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput350 la_oenb_mprj[66] vssd vccd wire1551/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput361 la_oenb_mprj[76] vssd vccd wire1541/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput372 la_oenb_mprj[86] vssd vccd wire1531/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput383 la_oenb_mprj[96] vssd vccd _593_/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput394 mprj_adr_o_core[15] vssd vccd wire1508/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_53_4103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__448__B _448_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1210_A _352_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output781_A _537_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1308_A wire1309/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output879_A wire1274/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2431 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3198 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2464 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput802 wire1048/X vssd vccd la_oenb_core[5] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput813 wire1047/X vssd vccd la_oenb_core[6] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput824 wire1046/X vssd vccd la_oenb_core[7] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_4249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput835 wire1045/X vssd vccd la_oenb_core[8] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput846 wire1044/X vssd vccd la_oenb_core[9] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput857 _323_/X vssd vccd mprj_adr_o_user[18] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1844_A wire1844/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput868 _333_/X vssd vccd mprj_adr_o_user[28] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput879 wire1274/X vssd vccd mprj_adr_o_user[9] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_3_4045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2104 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3322 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3272 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__358__B _358_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_2011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_2607 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_26 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_158 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_37 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_48 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_59 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3991 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3942 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_52_2244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_3244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1295 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2543 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_268 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_1369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_1831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1842 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input143_A la_iena_mprj[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2060_A wire2061/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1864 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1875 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_3968 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2158_A wire2158/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1886 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__549__A _549_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__268__B _268_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input310_A la_oenb_mprj[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input408_A mprj_adr_o_core[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_523_ _523_/A _523_/B vssd vccd _523_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_22_1391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_3864 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_454_ _582_/A _454_/B _454_/C vssd vccd _454_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__284__A _284_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_385_ _513_/A _385_/B _385_/C vssd vccd _385_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_16_1151 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1042 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3496 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3835 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__450__C _450_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3879 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_1628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1701 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1160_A wire1161/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_4229 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1258_A wire1259/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_2941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_290 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2816 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput180 la_iena_mprj[28] vssd vccd _191_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_42_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput191 la_iena_mprj[38] vssd vccd _201_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA__178__B _178_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1425_A wire1426/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] _204_/X vssd vccd _024_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_24_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3238 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__194__A _194_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1961_A wire1962/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2895 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3520 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput610 _100_/Y vssd vccd la_data_in_mprj[117] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput621 _110_/Y vssd vccd la_data_in_mprj[127] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput632 _004_/Y vssd vccd la_data_in_mprj[21] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput643 _014_/Y vssd vccd la_data_in_mprj[31] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput654 _024_/Y vssd vccd la_data_in_mprj[41] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput665 _034_/Y vssd vccd la_data_in_mprj[51] vssd vccd sky130_fd_sc_hd__buf_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] _166_/X vssd vccd _150_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xoutput676 _044_/Y vssd vccd la_data_in_mprj[61] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_3367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2108 wire2109/X vssd vccd _482_/B vssd vccd sky130_fd_sc_hd__buf_6
Xoutput687 _054_/Y vssd vccd la_data_in_mprj[71] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput698 _064_/Y vssd vccd la_data_in_mprj[81] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2119 wire2120/X vssd vccd _477_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_42_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1407 wire1408/X vssd vccd wire1407/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1418 wire1419/X vssd vccd wire1418/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1429 wire1430/X vssd vccd wire1429/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3717 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_170_ _170_/A _170_/B vssd vccd _170_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_52_1351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__551__B _551_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input260_A la_oenb_mprj[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_522 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input358_A la_oenb_mprj[73] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_566 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__380__A_N _508_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_599 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__279__A _279_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1930 wire1930/A vssd vccd wire1930/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1941 wire1942/X vssd vccd _602_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_1536 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1952 wire1952/A vssd vccd wire1952/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_935 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1963 wire1964/X vssd vccd _594_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1974 wire1974/A vssd vccd wire1974/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1985 wire1985/A vssd vccd wire1985/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4340 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1996 wire1997/X vssd vccd _576_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_230 _191_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_241 _166_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_4248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_506_ _506_/A _506_/B vssd vccd _506_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_252 _521_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_263 _467_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_274 _380_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_285 wire1428/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3558 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_296 wire1781/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_437_ _565_/A _437_/B _437_/C vssd vccd _437_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA__445__C _445_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1560 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_368_ _368_/A _368_/B vssd vccd _368_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_31_1413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output577_A _457_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1582 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_299_ _299_/A _299_/B vssd vccd _299_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__461__B _461_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output744_A _619_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1375_A wire1375/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4399 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2920 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] wire1325/X vssd vccd wire968/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_29_2098 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_2964 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1542_A wire1542/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__189__A _189_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1807_A wire1807/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_916 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_938 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire995_A _586_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_2470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_2481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_2323 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3956 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_676 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4119 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__B _371_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1729 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput473 wire1057/X vssd vccd la_data_in_core[109] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput484 _488_/X vssd vccd la_data_in_core[119] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput495 wire1131/X vssd vccd la_data_in_core[13] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_2535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1204 _354_/X vssd vccd wire1204/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1215 wire1216/X vssd vccd wire1215/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__099__A _099_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1226 wire1227/X vssd vccd wire1226/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1237 _343_/X vssd vccd wire1237/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1248 _339_/X vssd vccd wire1248/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1259 _322_/X vssd vccd wire1259/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_220 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__546__B _546_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input106_A la_data_out_mprj[77] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_908 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_993 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_222_ _222_/A _222_/B vssd vccd _222_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3422 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__562__A _562_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_1110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3444 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_153_ _153_/A vssd vccd _153_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_7_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input71_A la_data_out_mprj[45] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_084_ _084_/A vssd vccd _084_/Y vssd vccd sky130_fd_sc_hd__inv_4
XFILLER_45_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3963 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4324 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_3678 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1760 wire1760/A vssd vccd wire1760/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1771 wire1772/X vssd vccd _273_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1782 wire1783/X vssd vccd _267_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1793 wire1794/X vssd vccd _261_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_776 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__456__B _456_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_2345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1123_A _390_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_960 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_470 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output861_A _326_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[17\] mprj_dat_i_user[17] max_length1311/X vssd vccd _131_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XANTENNA_wire1492_A wire1493/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__191__B _191_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_3501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1757_A wire1758/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_3451 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1924_A wire1924/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_1058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] _278_/X vssd vccd wire984/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_39_3845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__366__B _366_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[95\]_B wire1319/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_4476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_805 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1001 _555_/X vssd vccd wire1001/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_878 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3860 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1012 _546_/X vssd vccd wire1012/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1023 _531_/X vssd vccd wire1023/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2282 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_2365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1034 _515_/X vssd vccd wire1034/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2218 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1045 _505_/X vssd vccd wire1045/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1056 _479_/X vssd vccd wire1056/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2140_A wire2140/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1067 _468_/X vssd vccd wire1067/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input223_A la_iena_mprj[67] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1078 _431_/X vssd vccd wire1078/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1089 _423_/X vssd vccd wire1089/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__557__A _557_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3809 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__276__B _276_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[86\]_B wire1328/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1227 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__A _292_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_205_ _205_/A _205_/B vssd vccd _205_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_11_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1552 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_136_ _136_/A vssd vccd _136_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_32_1574 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2562 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_4533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_067_ _067_/A vssd vccd _067_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_45_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4408 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_3061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1073_A _462_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4071 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2730 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_3497 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1590 wire1590/A vssd vccd _613_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_0_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__186__B _186_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1505_A wire1506/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_4465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[77\]_B _240_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_259 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1874_A wire1875/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2949 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_4225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_4308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2359 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__441__A_N _569_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_2433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1309 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2477 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2284 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1550 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4516 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3951 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3853 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_513 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3804 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3837 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_771 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input173_A la_iena_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2188_A wire2188/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1919 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1179 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3911 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2405 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3955 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input340_A la_oenb_mprj[57] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input438_A mprj_dat_o_core[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input34_A la_data_out_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3762 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__A _287_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_4004 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2927 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1614 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_579 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__453__C _453_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_output657_A _027_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_119_ _119_/A vssd vccd _119_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_wire1190_A wire1191/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2392 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_4100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__A_N _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output824_A wire1046/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1455_A wire1456/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] _234_/X vssd vccd _054_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_3_2847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1622_A wire1622/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__197__A _197_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3203 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1525 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2415 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1991_A wire1991/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_524 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_52_2437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2123 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_4138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_929 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_2539 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3069 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2335 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_470_ _598_/A _470_/B _470_/C vssd vccd _470_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_2_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_2793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4368 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[125\]_B _288_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__554__B _554_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2103_A wire2104/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input290_A la_oenb_mprj[127] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input388_A mprj_adr_o_core[0] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__487__A_N _615_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__570__A _570_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_4431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3982 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3616 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_1304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput340 la_oenb_mprj[57] vssd vccd _554_/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput351 la_oenb_mprj[67] vssd vccd wire1550/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput362 la_oenb_mprj[77] vssd vccd wire1540/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput373 la_oenb_mprj[87] vssd vccd wire1530/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput384 la_oenb_mprj[97] vssd vccd _594_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput395 mprj_adr_o_core[16] vssd vccd wire1504/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__448__C _448_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2880 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1061 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3403 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_4159 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_4279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1155 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1036_A _513_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2112 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_599_ _599_/A _599_/B vssd vccd _599_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_43_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__B _464_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[116\]_B _279_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4468 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1203_A wire1204/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output774_A wire1022/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_2590 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output941_A wire1235/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput803 wire997/X vssd vccd la_oenb_core[60] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput814 _567_/X vssd vccd la_oenb_core[70] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput825 _577_/X vssd vccd la_oenb_core[80] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput836 wire994/X vssd vccd la_oenb_core[90] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput847 _146_/Y vssd vccd mprj_ack_i_core vssd vccd sky130_fd_sc_hd__buf_8
Xoutput858 wire1257/X vssd vccd mprj_adr_o_user[19] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput869 _334_/X vssd vccd mprj_adr_o_user[29] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2909 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1837_A wire1838/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_3284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[25\]_A mprj_dat_i_user[25] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_1921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1965 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_126 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_16 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_2390 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XPHY_27 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_49 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_2089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1366 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4508 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[107\]_B wire1315/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__374__B _374_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_2808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_343 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2376 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3015 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2522 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2461 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2303 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_2555 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2599 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__549__B _549_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_1898 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2053_A wire2054/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input136_A la_iena_mprj[103] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_wb_dat_gates\[16\]_A mprj_dat_i_user[16] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_616 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_3409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_522_ _522_/A _522_/B vssd vccd _522_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_19_3832 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_2198 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input303_A la_oenb_mprj[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__565__A _565_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3876 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_453_ _581_/A _453_/B _453_/C vssd vccd _453_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3420 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_384_ _512_/A _384_/B _384_/C vssd vccd _384_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_1021 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1163 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1617 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4515 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_553 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_2308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_4377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output522_A wire1106/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_1101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__459__B _459_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1153_A _367_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput170 la_iena_mprj[19] vssd vccd _182_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput181 la_iena_mprj[29] vssd vccd _192_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_36_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_2193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput192 la_iena_mprj[39] vssd vccd _202_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_37_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1320_A _257_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1418_A wire1419/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_939 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_660 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] _197_/X vssd vccd _017_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
XFILLER_51_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__194__B _194_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1787_A wire1788/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2262 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1954_A wire1954/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput600 _091_/Y vssd vccd la_data_in_mprj[108] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput611 _101_/Y vssd vccd la_data_in_mprj[118] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput622 _159_/Y vssd vccd la_data_in_mprj[12] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput633 _005_/Y vssd vccd la_data_in_mprj[22] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3324 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput644 _015_/Y vssd vccd la_data_in_mprj[32] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput655 _025_/Y vssd vccd la_data_in_mprj[42] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_3576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xoutput666 _035_/Y vssd vccd la_data_in_mprj[52] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_3429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput677 _045_/Y vssd vccd la_data_in_mprj[62] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput688 _055_/Y vssd vccd la_data_in_mprj[72] vssd vccd sky130_fd_sc_hd__buf_8
Xwire2109 wire2109/A vssd vccd wire2109/X vssd vccd sky130_fd_sc_hd__buf_6
Xoutput699 _065_/Y vssd vccd la_data_in_mprj[82] vssd vccd sky130_fd_sc_hd__buf_8
Xwire1408 wire1408/A vssd vccd wire1408/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_42_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1419 wire1420/X vssd vccd wire1419/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__369__B _369_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_273 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1773 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_2427 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_4029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2741 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4452 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_641 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1926 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2351 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1071 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2170_A wire2170/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input253_A la_iena_mprj[94] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_8_3086 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_578 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1651 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input420_A mprj_cyc_o_core vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__279__B _279_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1920 wire1921/X vssd vccd wire1920/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1931 wire1932/X vssd vccd _606_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_3849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1942 wire1942/A vssd vccd wire1942/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1953 wire1954/X vssd vccd _597_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1964 wire1964/A vssd vccd wire1964/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1975 wire1975/A vssd vccd _587_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4330 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1986 wire1987/X vssd vccd _581_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1997 wire1997/A vssd vccd wire1997/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4352 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_220 _208_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_231 _191_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_505_ _505_/A _505_/B vssd vccd _505_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_50_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_242 _605_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_253 _521_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_264 _466_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_275 _522_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_286 _319_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_436_ _564_/A _436_/B _436_/C vssd vccd _436_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_18_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_297 wire1790/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_367_ _367_/A _367_/B vssd vccd _367_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_32_3873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_298_ _298_/A _298_/B vssd vccd _298_/X vssd vccd sky130_fd_sc_hd__and2_2
XANTENNA_output472_A wire1058/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__461__C _461_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3611 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output737_A _613_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1270_A _316_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_4141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3749 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1368_A wire1368/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4091 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__189__B _189_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1535_A wire1535/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2783 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1702_A wire1703/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_928 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2925 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__371__C _371_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_4052 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3419 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1391 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3143 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput463 wire1145/X vssd vccd la_data_in_core[0] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput474 wire1135/X vssd vccd la_data_in_core[10] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput485 wire1133/X vssd vccd la_data_in_core[11] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput496 wire1130/X vssd vccd la_data_in_core[14] vssd vccd sky130_fd_sc_hd__buf_8
Xwire1205 wire1206/X vssd vccd wire1205/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_25_2475 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1216 _350_/X vssd vccd wire1216/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1227 wire1228/X vssd vccd wire1227/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2328 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1238 wire1239/X vssd vccd wire1238/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1249 wire1250/X vssd vccd wire1249/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_4561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2260 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3893 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_2279 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2016_A wire2016/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3879 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_221_ _221_/A _221_/B vssd vccd _221_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_10_4146 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3592 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_152_ _152_/A vssd vccd _152_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3434 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__562__B _562_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3456 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1745 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_083_ _083_/A vssd vccd _083_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XANTENNA_input370_A la_oenb_mprj[84] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_1789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input64_A la_data_out_mprj[39] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_3975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_342 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2013 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4286 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_4369 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3635 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2057 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1750 wire1750/A vssd vccd wire1750/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1761 wire1762/X vssd vccd _278_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1772 wire1772/A vssd vccd wire1772/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1783 wire1783/A vssd vccd wire1783/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1794 wire1794/A vssd vccd wire1794/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_34_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__456__C _456_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1116_A _397_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output687_A _054_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_419_ _547_/A _419_/B _419_/C vssd vccd _419_/X vssd vccd sky130_fd_sc_hd__and3b_2
XFILLER_50_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2644 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__472__B _472_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_2519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2699 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output854_A wire1261/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1485_A wire1486/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_3513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1652_A wire1653/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_4028 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3463 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2604 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2041 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1026 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1917_A wire1918/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2659 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] _271_/X vssd vccd wire990/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_17_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_4157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__370__A_N _498_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__382__B _382_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[8\]_A mprj_dat_i_user[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1002 wire1003/X vssd vccd wire1002/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2344 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1013 wire1014/X vssd vccd wire1013/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_3933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3872 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1024 _530_/X vssd vccd wire1024/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1035 _514_/X vssd vccd wire1035/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_2377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1046 _504_/X vssd vccd wire1046/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1057 _478_/X vssd vccd wire1057/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1068 _467_/X vssd vccd wire1068/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1079 _430_/X vssd vccd wire1079/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2133_A wire2134/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input216_A la_iena_mprj[60] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_585 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3643 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__573__A _573_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_204_ _204_/A _204_/B vssd vccd _204_/X vssd vccd sky130_fd_sc_hd__and2_1
XFILLER_12_975 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3220 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__292__B _292_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_135_ _135_/A vssd vccd _135_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_49_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1586 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_066_ _066_/A vssd vccd _066_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_23_4304 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_3750 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_3708 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_4100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_3073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4050 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3360 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_3432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA__467__B _467_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1580 wire1580/A vssd vccd _623_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1591 wire1591/A vssd vccd _612_/A vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1233_A wire1234/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_53 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__393__A_N _521_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1400_A wire1400/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2029 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2906 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_2463 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1867_A wire1868/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_4011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_2868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1446 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1064 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2506 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_861 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__B _377_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_352 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_3963 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3540 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4296 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_271 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1873 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3584 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1895 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input166_A la_iena_mprj[15] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2083_A wire2084/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3923 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_3967 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_654 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4453 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input333_A la_oenb_mprj[50] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3680 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__A _568_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input27_A la_data_out_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__287__B _287_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1326 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_1298 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4152 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4016 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1751 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4196 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3304 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2349 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_3397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_242 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_253 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_118_ _118_/A vssd vccd _118_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_output552_A _434_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_4112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_049_ _049_/A vssd vccd _049_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_7_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1183_A wire1184/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_4134 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3591 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output817_A _570_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1350_A wire1351/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1448_A wire1449/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1007 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1187 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] _227_/X vssd vccd _047_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_1_3295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3117 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1984_A wire1985/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire970_A wire970/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_2293 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_2747 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2135 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1423 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3208 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_2461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2347 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_2286 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2082 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_4325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_3050 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3624 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1334 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input283_A la_oenb_mprj[120] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__570__B _570_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_1080 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_2691 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input450_A mprj_dat_o_core[7] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_4443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3731 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3994 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1513 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput330 la_oenb_mprj[48] vssd vccd _417_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__298__A _298_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput341 la_oenb_mprj[58] vssd vccd wire1556/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput352 la_oenb_mprj[68] vssd vccd wire1549/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput363 la_oenb_mprj[78] vssd vccd wire1539/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput374 la_oenb_mprj[88] vssd vccd wire1529/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_29_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput385 la_oenb_mprj[98] vssd vccd wire1528/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput396 mprj_adr_o_core[17] vssd vccd wire1500/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_35_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1145 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2703 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_3459 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_4425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1029_A _520_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_598_ _598_/A _598_/B vssd vccd _598_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_38_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__464__C _464_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3112 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_2157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__431__A_N _559_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output767_A wire1025/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_3178 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_4404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1398_A wire1399/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__480__B _480_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4207 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_1 la_data_out_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput804 wire996/X vssd vccd la_oenb_core[61] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_output934_A wire1154/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput815 _568_/X vssd vccd la_oenb_core[71] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput826 _578_/X vssd vccd la_oenb_core[81] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2930 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput837 _588_/X vssd vccd la_oenb_core[91] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_6_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1565_A _409_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3758 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput848 _305_/X vssd vccd mprj_adr_o_user[0] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1205 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_2963 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xoutput859 _306_/X vssd vccd mprj_adr_o_user[1] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4058 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1732_A wire1733/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[25\]_B _294_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_3092 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1955 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_17 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3922 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1378 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2989 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__390__B _390_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1854 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2534 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1800 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2567 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_2359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[16\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2046_A wire2046/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input129_A la_data_out_mprj[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_127 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1994 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_521_ _521_/A _521_/B vssd vccd _521_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_2_1476 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__565__B _565_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_4100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_452_ _580_/A _452_/B _452_/C vssd vccd _452_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_17_4280 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3888 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__454__A_N _582_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_383_ _511_/A _383_/B _383_/C vssd vccd _383_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_25_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_355 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3432 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input94_A la_data_out_mprj[66] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_359 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__A _581_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1175 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_3677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_2088 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_281 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3688 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__459__C _459_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output515_A wire1113/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput160 la_iena_mprj[125] vssd vccd _288_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2976 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput171 la_iena_mprj[1] vssd vccd _164_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput182 la_iena_mprj[2] vssd vccd _165_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_797 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput193 la_iena_mprj[3] vssd vccd _166_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1146_A wire1147/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3332 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__475__B _475_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1313_A _286_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_1529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] _190_/X vssd vccd _010_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_32_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2831 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1682_A wire1683/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_1117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput601 _092_/Y vssd vccd la_data_in_mprj[109] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput612 _102_/Y vssd vccd la_data_in_mprj[119] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput623 _160_/Y vssd vccd la_data_in_mprj[13] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput634 _006_/Y vssd vccd la_data_in_mprj[23] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput645 _016_/Y vssd vccd la_data_in_mprj[33] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput656 _026_/Y vssd vccd la_data_in_mprj[43] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3336 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput667 _036_/Y vssd vccd la_data_in_mprj[53] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2782 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput678 _046_/Y vssd vccd la_data_in_mprj[63] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput689 _056_/Y vssd vccd la_data_in_mprj[73] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1409 wire1410/X vssd vccd _311_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__369__C _369_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_937 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__477__A_N _477_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_970 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__385__B _385_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_2010 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1916 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3796 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1083 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_4413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2375 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input246_A la_iena_mprj[88] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2163_A wire2164/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1910 wire1910/A vssd vccd wire1910/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1921 wire1921/A vssd vccd wire1921/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1932 wire1933/X vssd vccd wire1932/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1943 wire1944/X vssd vccd _601_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1954 wire1954/A vssd vccd wire1954/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1965 wire1966/X vssd vccd _593_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1308 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1976 wire1976/A vssd vccd _586_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input413_A mprj_adr_o_core[3] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1987 wire1987/A vssd vccd wire1987/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__576__A _576_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1998 wire1999/X vssd vccd _575_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4364 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_210 _232_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_221 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3652 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_504_ _504_/A _504_/B vssd vccd _504_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_232 _191_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__295__B _295_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_243 _605_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_254 _521_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_3696 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_265 la_data_out_core[47] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_276 _557_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_287 _318_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_435_ _563_/A _435_/B _435_/C vssd vccd _435_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_37_1849 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2241 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_298 wire1888/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_366_ _366_/A _366_/B vssd vccd _366_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_31_2138 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_3885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_297_ _297_/A _297_/B vssd vccd _297_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_35_1595 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output465_A wire1065/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1096_A _417_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3706 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_3645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1263_A _319_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_1533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_3305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_49_561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2751 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2762 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2521 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1430_A wire1431/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1914 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_3020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_214 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_992 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_748 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_3097 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1897_A wire1897/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_2937 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_612 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_2374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_50_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_3373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3100 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_3205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3374 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput464 wire1066/X vssd vccd la_data_in_core[100] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput475 wire1056/X vssd vccd la_data_in_core[110] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_2651 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_3166 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput486 _489_/X vssd vccd la_data_in_core[120] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput497 wire1129/X vssd vccd la_data_in_core[15] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1206 wire1207/X vssd vccd wire1206/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input1_A caravel_clk vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1217 wire1218/X vssd vccd wire1217/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1228 _346_/X vssd vccd wire1228/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1239 wire1240/X vssd vccd wire1239/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_28_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2272 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3803 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1593 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_220_ _220_/A _220_/B vssd vccd _220_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_4125 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3571 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2009_A wire2009/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_151_ _151_/A vssd vccd _151_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XANTENNA_input196_A la_iena_mprj[42] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_177 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_3468 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1757 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_082_ _082_/A vssd vccd _082_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_45_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input363_A la_oenb_mprj[78] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input57_A la_data_out_mprj[32] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_398 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2025 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3553 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4298 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_701 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1740 wire1741/X vssd vccd _288_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_4_2069 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2924 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1751 wire1752/X vssd vccd _283_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1897 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1274 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1762 wire1762/A vssd vccd wire1762/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1773 wire1774/X vssd vccd _272_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2946 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1784 wire1784/A vssd vccd _266_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1795 wire1796/X vssd vccd _260_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_4003 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_266 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_789 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_737 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_418_ _546_/A _418_/B _418_/C vssd vccd _418_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_42_792 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1011_A wire1012/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_932 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output582_A wire1074/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1067 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_wire1109_A _404_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1813 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_3693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_349_ _349_/A _349_/B vssd vccd _349_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_35_1381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1478_A wire1479/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] wire1320/X vssd vccd wire963/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_3306 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3475 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1645_A wire1645/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_3124 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1812_A wire1812/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_4169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_2881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__382__C _382_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_wb_dat_gates\[8\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_3160 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2527 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_2481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2885 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xwire1003 _553_/X vssd vccd wire1003/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_user_to_mprj_in_gates\[8\]_B _171_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1014 _542_/X vssd vccd wire1014/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1025 _525_/X vssd vccd wire1025/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_3884 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1036 _513_/X vssd vccd wire1036/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1047 _503_/X vssd vccd wire1047/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1058 _477_/X vssd vccd wire1058/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1069 _466_/X vssd vccd wire1069/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1519 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input111_A la_data_out_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input209_A la_iena_mprj[54] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2126_A wire2127/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4367 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4378 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1354 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__573__B _573_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_203_ _203_/A _203_/B vssd vccd _203_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_10_3210 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_987 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3232 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_134_ _134_/A vssd vccd _134_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_065_ _065_/A vssd vccd _065_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_49_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_641 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_151 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_4281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_4156 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3383 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1059_A _476_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1570 wire1570/A vssd vccd _529_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_39_2409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1581 wire1581/A vssd vccd _622_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1592 wire1592/A vssd vccd _611_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_0_1018 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1226_A wire1227/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output797_A wire1004/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_4309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__B _483_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_2420 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_wb_dat_gates\[22\] mprj_dat_i_user[22] max_length1310/X vssd vccd _136_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_50_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2918 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1762_A wire1762/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2814 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3250 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3283 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2402 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] _283_/X vssd vccd _103_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_29_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__377__C _377_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_4501 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3920 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_331 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_53_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_876 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3817 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__B _393_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_3574 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_283 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_3596 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_1295 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2076_A wire2077/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_2379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input159_A la_iena_mprj[124] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_24_3979 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_3720 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_637 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2164 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__568__B _568_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1981 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3692 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_input326_A la_oenb_mprj[44] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3775 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_2197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_1391 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1316 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_1889 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__584__A _584_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_4164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4066 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2317 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_4028 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_1140 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2620 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3316 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1184 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1026 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1059 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_1985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_265 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_117_ _117_/A vssd vccd _117_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_29_3846 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_048_ _048_/A vssd vccd _048_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_4_961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output545_A wire1081/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1176_A wire1177/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1111 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output712_A _077_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__478__B _478_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1343_A wire1343/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1019 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_1199 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire2090 wire2090/A vssd vccd wire2090/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_26_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] _220_/X vssd vccd _040_/A vssd vccd
+ sky130_fd_sc_hd__nand2_2
XFILLER_36_3817 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_821 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1510_A wire1511/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_1505 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vccd vccd vssd
+ sky130_fd_sc_hd__diode_2
XFILLER_39_1549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_4117 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1977_A wire1978/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1435 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_4057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3378 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3389 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__388__B _388_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_681 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1048 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_301 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1382 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4397 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3062 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3636 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_2962 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1346 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4072 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_570 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_3961 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3360 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1660 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1693 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2193_A wire2193/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input276_A la_oenb_mprj[114] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3940 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4455 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__383__A_N _511_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_931 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input443_A mprj_dat_o_core[2] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_2237 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_4499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__579__A _579_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4240 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3848 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_3787 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput320 la_oenb_mprj[39] vssd vccd _536_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput331 la_oenb_mprj[49] vssd vccd _546_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_40_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput342 la_oenb_mprj[59] vssd vccd _556_/A vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA__298__B _298_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_1569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput353 la_oenb_mprj[69] vssd vccd wire1548/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput364 la_oenb_mprj[79] vssd vccd wire1538/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput375 la_oenb_mprj[89] vssd vccd _586_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_29_93 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput386 la_oenb_mprj[99] vssd vccd wire1527/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput397 mprj_adr_o_core[18] vssd vccd wire1497/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_48_489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_81 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_597_ _597_/A _597_/B vssd vccd _597_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_43_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2759 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2136 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output495_A wire1131/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2169 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3168 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_581 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output662_A _032_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_4416 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__480__C _480_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_3621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_2 la_data_out_core[10] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput805 _559_/X vssd vccd la_oenb_core[62] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_6_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput816 _569_/X vssd vccd la_oenb_core[72] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput827 _579_/X vssd vccd la_oenb_core[82] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput838 _589_/X vssd vccd la_oenb_core[92] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output927_A wire1182/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput849 wire1271/X vssd vccd mprj_adr_o_user[10] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_6_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1460_A wire1461/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_1490 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1558_A _420_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_2760 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2613 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1725_A wire1725/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_106 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3625 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_18 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_29 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4061 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_857 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1811 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1833 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1888 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_728 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2579 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_1709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1085 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_520_ _520_/A _520_/B vssd vccd _520_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_17_139 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2039_A wire2039/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_451_ _579_/A _451_/B _451_/C vssd vccd _451_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_35_2401 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_109 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_4292 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_3400 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_382_ _510_/A _382_/B _382_/C vssd vccd _382_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_15_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2206_A wire2207/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_305 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_153 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_367 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2489 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input393_A mprj_adr_o_core[14] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_349 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__581__B _581_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input87_A la_data_out_mprj[5] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_1187 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4263 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1548 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_4116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3792 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3404 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__102__A _102_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_721 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3437 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3448 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput150 la_iena_mprj[116] vssd vccd _279_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput161 la_iena_mprj[126] vssd vccd _289_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput172 la_iena_mprj[20] vssd vccd _183_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_4_2988 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput183 la_iena_mprj[30] vssd vccd _193_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4012 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output508_A wire1119/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3901 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput194 la_iena_mprj[40] vssd vccd _203_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XANTENNA_wire1041_A _508_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1139_A _375_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_3213 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_3344 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3235 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_3809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4201 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output877_A wire1277/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__491__B _491_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_2843 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1276 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_2865 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1129 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4224 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1675_A wire1675/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput602 _157_/Y vssd vccd la_data_in_mprj[10] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_4268 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput613 _158_/Y vssd vccd la_data_in_mprj[11] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput624 _161_/Y vssd vccd la_data_in_mprj[14] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput635 _007_/Y vssd vccd la_data_in_mprj[24] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput646 _017_/Y vssd vccd la_data_in_mprj[34] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput657 _027_/Y vssd vccd la_data_in_mprj[44] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1842_A wire1842/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput668 _037_/Y vssd vccd la_data_in_mprj[54] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1648 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xoutput679 _047_/Y vssd vccd la_data_in_mprj[64] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2794 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1225 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3119 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_3731 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_2629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_698 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_197 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_3921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2282 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_3871 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3713 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2387 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1412 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1900 wire1901/X vssd vccd wire1900/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input141_A la_iena_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1911 wire1912/X vssd vccd _612_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_3_4390 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1922 wire1923/X vssd vccd _609_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2156_A wire2157/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input239_A la_iena_mprj[81] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1933 wire1933/A vssd vccd wire1933/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__421__A_N _549_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1944 wire1944/A vssd vccd wire1944/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1955 wire1956/X vssd vccd _596_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1966 wire1966/A vssd vccd wire1966/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4321 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1977 wire1978/X vssd vccd _585_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1988 wire1989/X vssd vccd _580_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1999 wire2000/X vssd vccd wire1999/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__576__B _576_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input406_A mprj_adr_o_core[26] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_200 _262_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_211 _232_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_503_ _503_/A _503_/B vssd vccd _503_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_222 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_233 _186_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_244 _605_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_429 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_255 wire2071/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3528 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_266 mprj_dat_i_user[29] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_434_ _562_/A _434_/B _434_/C vssd vccd _434_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_277 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_288 _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_299 wire1904/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2253 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__592__A _592_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_1238 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_365_ _365_/A _365_/B vssd vccd _365_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_9_113 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2297 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_296_ _296_/A _296_/B vssd vccd _296_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_3296 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1449 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4347 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_3718 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1089_A _423_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[40\]_B _203_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3212 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3464 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1256_A _325_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_3245 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2741 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_2605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_2533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_3289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1589 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__486__B _486_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_2566 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1423_A wire1424/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_36_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_705 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_727 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3753 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_982 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_289 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3043 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1792_A wire1792/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_3341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_2348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3948 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_3385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1062 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__007__A _007_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_3331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] _164_/X vssd vccd _148_/A vssd vccd
+ sky130_fd_sc_hd__nand2_1
Xoutput465 wire1065/X vssd vccd la_data_in_core[101] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_B _194_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput476 wire1055/X vssd vccd la_data_in_core[111] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA__444__A_N _572_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput487 _490_/X vssd vccd la_data_in_core[121] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_9_2663 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput498 wire1128/X vssd vccd la_data_in_core[16] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3178 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1207 _353_/X vssd vccd wire1207/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1218 wire1219/X vssd vccd wire1218/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1229 wire1230/X vssd vccd wire1229/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_9_1995 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2499 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_4229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_713 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_746 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__396__B _396_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_757 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2284 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1561 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3815 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[98\]_B _261_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_14_4240 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3848 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_440 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_963 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_2573 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2437 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_150_ _150_/A vssd vccd _150_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_11_657 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_081_ _081_/A vssd vccd _081_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_12_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input189_A la_iena_mprj[36] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1471 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_845 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input356_A la_oenb_mprj[71] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3808 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_B _185_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2173 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_3532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_2577 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_2037 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__587__A _587_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_3565 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_1483 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1730 wire1731/X vssd vccd wire1730/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1741 wire1741/A vssd vccd wire1741/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1752 wire1752/A vssd vccd wire1752/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1763 wire1764/X vssd vccd _277_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1774 wire1774/A vssd vccd wire1774/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_20_1128 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1785 wire1786/X vssd vccd _265_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_245 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_768 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_4151 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1796 wire1796/A vssd vccd wire1796/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4184 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_749 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[89\]_B wire1325/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_417_ _417_/A_N _417_/B _417_/C vssd vccd _417_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_18_1035 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_81 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_3661 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1079 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_348_ _348_/A _348_/B vssd vccd _348_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_wire1004_A _552_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2679 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output575_A _455_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_3093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_1393 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_279_ _279_/A _279_/B vssd vccd _279_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_13_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__467__A_N _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output742_A _617_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_3410 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1373_A wire1374/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] wire1327/X vssd vccd wire970/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_22_3318 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_3487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1540_A wire1540/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3250 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1638_A wire1638/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__497__A _497_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_2560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2363 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_2396 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_4137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_568 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_4560 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1102 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4424 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2270 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_2194 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_988 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_3193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3218 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3172 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2539 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2493 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1004 _552_/X vssd vccd wire1004/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1015 _541_/X vssd vccd wire1015/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1026 _523_/X vssd vccd wire1026/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1037 _512_/X vssd vccd wire1037/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_47_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1048 _502_/X vssd vccd wire1048/X vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__200__A _200_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1059 _476_/X vssd vccd wire1059/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_3325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_4302 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3623 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input104_A la_data_out_mprj[75] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_1945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2119_A wire2120/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_3656 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_3509 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1978 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2381 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1989 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_202_ _202_/A _202_/B vssd vccd _202_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_51_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_1219 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1500 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_999 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3244 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_133_ _133_/A vssd vccd _133_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_10_2532 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2543 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4431 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_064_ _064_/A vssd vccd _064_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_653 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_174 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_4293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_1673 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1291 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2722 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__110__A _110_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_21_2650 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_3395 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1560 input33/X vssd vccd _495_/C vssd vccd sky130_fd_sc_hd__buf_6
Xwire1571 _400_/A_N vssd vccd _528_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1582 wire1582/A vssd vccd _621_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1593 wire1593/A vssd vccd _610_/A vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_1_2788 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1121_A _392_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_557 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output692_A _059_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_719 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire1219_A _349_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_2009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__483__C _483_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_3166 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_wb_dat_gates\[15\] mprj_dat_i_user[15] max_length1311/X vssd vccd _129_/A vssd
+ vccd sky130_fd_sc_hd__nand2_4
XFILLER_31_1021 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1490_A wire1491/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1065 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1755_A wire1756/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3262 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_3104 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_2149 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1922_A wire1923/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_3389 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2414 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2666 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_2458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__020__A _020_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1807 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] _276_/X vssd vccd wire986/A vssd
+ vccd sky130_fd_sc_hd__nand2_2
XFILLER_53_822 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_373 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_4081 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3932 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3976 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_1597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__393__C _393_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_2521 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4232 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_785 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_295 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1263 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_3109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2303 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3048 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2661 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_4444 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_wire2069_A wire2070/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_3660 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_2176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_2029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input221_A la_iena_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3798 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input319_A la_oenb_mprj[38] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_38_3133 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4012 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4132 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__584__B _584_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_888 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4078 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1628 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_2605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1038 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_116_ _116_/A vssd vccd _116_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_51_1997 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1385 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3858 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__105__A _105_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_047_ _047_/A vssd vccd _047_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_4_973 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_3571 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_461 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output538_A wire1091/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3529 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2892 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1071_A _464_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1217 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2080 wire2081/X vssd vccd wire2080/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire2091 wire2092/X vssd vccd _488_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1336_A input96/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_351 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1390 wire1390/A vssd vccd wire1390/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_36_3829 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_833 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__494__B _494_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[119\]_B _282_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_4265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_877 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1503_A wire1504/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_17_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2538 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_2549 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2841 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_3851 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2738 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_50_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1872_A wire1873/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_2601 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_3418 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_2645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1933 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_3070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_2801 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_A mprj_dat_i_user[28] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__388__C _388_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_2485 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_800 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_693 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_3317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2073 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_4305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_899 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_2941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_3074 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_357 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2974 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1358 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_4084 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_3973 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3372 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_1672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_3413 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2671 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xmax_length1310 _294_/X vssd vccd max_length1310/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_2409 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_49_1101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_3457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input171_A la_iena_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input269_A la_oenb_mprj[108] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire2186_A wire2187/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_921 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__579__B _579_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input436_A mprj_dat_o_core[23] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_user_wb_dat_gates\[19\]_A mprj_dat_i_user[19] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_3045 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput310 la_oenb_mprj[2] vssd vccd _499_/A vssd vccd sky130_fd_sc_hd__buf_4
Xinput321 la_oenb_mprj[3] vssd vccd _500_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_1_987 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_3799 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_413 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input32_A la_data_out_mprj[125] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_486 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput332 la_oenb_mprj[4] vssd vccd _501_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1318 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput343 la_oenb_mprj[5] vssd vccd _502_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4285 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_3089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput354 la_oenb_mprj[6] vssd vccd _503_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput365 la_oenb_mprj[7] vssd vccd _504_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_457 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1621 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput376 la_oenb_mprj[8] vssd vccd _505_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput387 la_oenb_mprj[9] vssd vccd _506_/A vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_21_1020 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput398 mprj_adr_o_core[19] vssd vccd wire1493/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__595__A _595_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_40_1665 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_596_ _596_/A _596_/B vssd vccd _596_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_32_803 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_93 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_3130 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_4449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2148 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_51_3185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_2402 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_3158 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output488_A _491_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_1469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3633 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output655_A _025_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_3 la_data_out_core[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_3081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput806 _560_/X vssd vccd la_oenb_core[63] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput817 _570_/X vssd vccd la_oenb_core[73] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_6_65 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput828 _580_/X vssd vccd la_oenb_core[83] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1286_A wire1287/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_7_4141 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_2943 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput839 _590_/X vssd vccd la_oenb_core[93] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output822_A _575_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2233 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4185 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3210 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_3473 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__489__B _489_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1453_A wire1454/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_23_2542 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1620_A wire1620/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_2669 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3637 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XPHY_19 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_652 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_4073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_685 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_379 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_1558 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_1569 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1211 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_1845 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_3733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1255 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_3777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_3176 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_206 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__399__B _399_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_44_1020 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_4561 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4503 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_2293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2124 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4536 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_3824 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1445 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_450_ _578_/A _450_/B _450_/C vssd vccd _450_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_26_685 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_381_ _509_/A _381_/B _381_/C vssd vccd _381_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_40_121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_346 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire2101_A wire2101/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_9_317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1122 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_4209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_379 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_4482 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input386_A la_oenb_mprj[99] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_3781 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_1199 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_4507 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_2829 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3760 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_4275 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2597 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1301 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3563 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1345 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput140 la_iena_mprj[107] vssd vccd _270_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_23_1115 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput151 la_iena_mprj[117] vssd vccd _280_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_49_777 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xinput162 la_iena_mprj[127] vssd vccd _290_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput173 la_iena_mprj[21] vssd vccd _184_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput184 la_iena_mprj[31] vssd vccd _194_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput195 la_iena_mprj[41] vssd vccd _204_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_18_4024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_3913 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_4035 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_2680 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_630 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2691 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4068 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_3957 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2611 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3356 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_4393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3269 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_2535 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_2081 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_579_ _579_/A _579_/B vssd vccd _579_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_4257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2677 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1211 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output772_A _529_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XPHY_190 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__491__C _491_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_2287 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4236 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_4186 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput603 _093_/Y vssd vccd la_data_in_mprj[110] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput614 _103_/Y vssd vccd la_data_in_mprj[120] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1668_A wire1669/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_25_4039 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput625 _162_/Y vssd vccd la_data_in_mprj[15] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_25_3305 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput636 _008_/Y vssd vccd la_data_in_mprj[25] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_29_3485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_1616 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xoutput647 _018_/Y vssd vccd la_data_in_mprj[35] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput658 _028_/Y vssd vccd la_data_in_mprj[45] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_45_2041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput669 _038_/Y vssd vccd la_data_in_mprj[55] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1835_A wire1836/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2350 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_3189 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_2394 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_2477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_909 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3445 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_4422 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_3710 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__373__A_N _501_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_110 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_121 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4308 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_655 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4488 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4529 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_309 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_2311 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_537 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_4404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__203__A _203_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_3933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2737 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_2355 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4448 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_4459 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3977 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1901 wire1901/A vssd vccd wire1901/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_41_3173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1424 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1912 wire1913/X vssd vccd wire1912/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1923 wire1924/X vssd vccd wire1923/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1934 wire1935/X vssd vccd _605_/B vssd vccd sky130_fd_sc_hd__buf_6
Xwire1945 wire1946/X vssd vccd _600_/B vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_917 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input134_A la_iena_mprj[101] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1956 wire1956/A vssd vccd wire1956/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2051_A wire2051/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1967 wire1968/X vssd vccd _592_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire2149_A wire2150/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1978 wire1978/A vssd vccd wire1978/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1989 wire1989/A vssd vccd wire1989/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_438 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_1793 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_201 _262_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_502_ _502_/A _502_/B vssd vccd _502_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_19_4388 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_212 _230_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input301_A la_oenb_mprj[21] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_22_1192 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_223 _205_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_234 _186_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_27_972 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_245 _570_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_460 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_256 wire2111/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1818 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_433_ _561_/A _433_/B _433_/C vssd vccd _433_/X vssd vccd sky130_fd_sc_hd__and3b_4
XANTENNA_267 wire2192/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_35_2221 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_278 _344_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_289 _570_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_441 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__592__B _592_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_4577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_364_ _364_/A _364_/B vssd vccd _364_/X vssd vccd sky130_fd_sc_hd__and2_2
XFILLER_35_2265 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_125 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2129 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_4017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3264 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_295_ _295_/A_N _295_/B vssd vccd _295_/X vssd vccd sky130_fd_sc_hd__and2b_2
XFILLER_26_4315 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_4409 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_4359 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1925 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_26_2902 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1407 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_46_2361 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1969 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3432 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_4019 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_output520_A wire1108/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_2269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output618_A _107_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_3476 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_3257 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1151_A wire1152/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1249_A wire1250/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA__486__C _486_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_1905 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__396__A_N _524_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_37_3721 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_3011 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire1416_A wire1416/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_3142 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_3765 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3164 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] _195_/X vssd vccd _015_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_18_3175 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_953 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_1317 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_4054 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3353 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_53_1653 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_1675 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1785_A wire1786/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_53_1686 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_1074 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4044 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_3861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_3725 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4077 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_3343 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4099 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__023__A _023_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput466 wire1064/X vssd vccd la_data_in_core[102] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput477 wire1054/X vssd vccd la_data_in_core[112] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_5_3229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput488 _491_/X vssd vccd la_data_in_core[122] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput499 wire1127/X vssd vccd la_data_in_core[17] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_47_1479 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2467 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_3493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1208 wire1209/X vssd vccd wire1208/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_5_1805 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_1170 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1001 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1219 _349_/X vssd vccd wire1219/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_45_1181 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2230 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1849 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_2241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_725 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_3841 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3780 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__396__C _396_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_1089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_769 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_780 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_3827 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2541 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_4252 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_975 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_4274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2405 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_4116 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_2585 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_3404 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_3584 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_2449 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4337 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_1103 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_1163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_629 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_080_ _080_/A vssd vccd _080_/Y vssd vccd sky130_fd_sc_hd__clkinv_4
XFILLER_17_1294 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_49_2913 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2195 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_97 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2099_A wire2100/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_3_857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_5_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2501 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4212 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_2681 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_input251_A la_iena_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_input349_A la_oenb_mprj[65] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2545 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_21_4256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_2589 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_1221 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1720 wire1721/X vssd vccd _294_/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA__587__B _587_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire1731 wire1731/A vssd vccd wire1731/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_3577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_3588 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1742 wire1743/X vssd vccd _287_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1753 wire1754/X vssd vccd _282_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1764 wire1764/A vssd vccd wire1764/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_46_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1775 wire1776/X vssd vccd _271_/A vssd vccd sky130_fd_sc_hd__buf_6
Xwire1786 wire1786/A vssd vccd wire1786/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_37_3017 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2959 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1797 wire1797/A vssd vccd _259_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_4163 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4196 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_3949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_430 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_4341 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3348 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_986 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_416_ _416_/A_N _416_/B _416_/C vssd vccd _416_/X vssd vccd sky130_fd_sc_hd__and3b_4
XFILLER_50_2505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_1047 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2073 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__108__A _108_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_30_945 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_2549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_2095 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
X_347_ _347_/A _347_/B vssd vccd _347_/X vssd vccd sky130_fd_sc_hd__and2_4
X_278_ _278_/A _278_/B vssd vccd _278_/X vssd vccd sky130_fd_sc_hd__and2_4
XANTENNA_output470_A wire1060/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_3960 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output568_A wire1138/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_13_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_3709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_3157 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_4123 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1199_A wire1200/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output735_A _611_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1733 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_1121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3527 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_4481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_48_1777 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1366_A wire1366/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2033 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_2618 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_4517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__497__B _497_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_wire1533_A wire1533/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_3137 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1365 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_2572 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_2331 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1700_A wire1701/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_514 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1746 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_547 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_4572 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_901 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire986_A wire986/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_4436 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3882 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3773 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_3724 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_433 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_14_1423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_53_1494 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__411__A_N _539_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_49_2209 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_1770 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2507 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_4109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_2821 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_3184 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_4532 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_2865 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_22_4576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1005 wire1006/X vssd vccd wire1005/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_40_2729 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1016 wire1017/X vssd vccd wire1016/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_38_4005 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1027 _522_/X vssd vccd wire1027/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1038 _511_/X vssd vccd wire1038/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire1049 _501_/X vssd vccd wire1049/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_0_4383 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_4325 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_205 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_1381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_51_4249 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_249 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_709 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_761 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1957 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_3668 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_4060 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2014_A wire2014/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_19_1345 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_51_2825 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_260 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_271 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2213 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4101 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2847 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2393 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_201_ _201_/A _201_/B vssd vccd _201_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_11_433 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_293 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_2869 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1512 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_4145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input299_A la_oenb_mprj[1] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
X_132_ _132_/A vssd vccd _132_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_8_949 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_477 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2511 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_3256 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_063_ _063_/A vssd vccd _063_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_10_3289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_4443 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_10_2577 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_4537 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input62_A la_data_out_mprj[37] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_48_1029 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_4487 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_3_665 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1917 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__598__A _598_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_43_2353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_809 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_4169 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xwire1550 wire1550/A vssd vccd _564_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_533 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xwire1561 wire1561/A vssd vccd _544_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2662 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xwire1572 wire1572/A vssd vccd _527_/A vssd vccd sky130_fd_sc_hd__buf_8
Xwire1583 wire1583/A vssd vccd _620_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_19_555 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1594 wire1594/A vssd vccd _609_/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_1_2756 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1009 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3893 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_1401 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_569 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_2179 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_2411 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA__434__A_N _562_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_32_3481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_2319 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_15_2499 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_1645 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output852_A wire1264/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1033 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1689 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1483_A wire1484/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_1077 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_4025 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_4036 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1541 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1650_A wire1651/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_3274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_3357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_2634 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_2426 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__301__A _301_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_39_4325 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_4_3070 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1933 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1915_A wire1916/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_42_1173 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_4369 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_0_2200 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] _269_/X vssd vccd _089_/A vssd
+ vccd sky130_fd_sc_hd__nand2_8
XFILLER_37_385 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3944 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_4200 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_13_3808 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_3988 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2533 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_4244 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_742 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_50_3581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_33_2588 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_797 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_2017 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4053 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_2315 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_4097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_2359 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_4423 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_2280 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_4373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2673 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__211__A _211_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_105 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2008 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1371 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_47_149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3101 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1869 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_3145 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input214_A la_iena_mprj[59] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_16_514 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_897 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__457__A_N _585_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_51_4024 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_3009 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_3189 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_4057 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_38_1765 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_51_2633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1921 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4505 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_234 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1353 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4549 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3241 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_115_ _115_/A vssd vccd _115_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_3105 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_1397 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_3285 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_4251 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
X_046_ _046_/A vssd vccd _046_/Y vssd vccd sky130_fd_sc_hd__clkinv_2
XFILLER_45_3149 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1861 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_3583 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_473 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3458 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__121__A _121_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_1135 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_3761 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_617 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_1229 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1064_A _471_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2070 wire2071/X vssd vccd wire2070/X vssd vccd sky130_fd_sc_hd__buf_6
Xwire2081 wire2081/A vssd vccd wire2081/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_36_4509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output600_A _091_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xwire2092 wire2093/X vssd vccd wire2092/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_43_1493 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1380 wire1380/A vssd vccd wire1380/X vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_21_2481 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_2492 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xwire1391 wire1392/X vssd vccd _337_/B vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_wire1231_A _345_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_1_1830 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1329_A _248_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_52_3109 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__494__C _494_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_1_1885 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_4277 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_2517 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4520 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_2853 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_4564 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_2717 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1698_A wire1699/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_15_2274 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_3863 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_3896 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_1453 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1865_A wire1866/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_790 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_4237 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3121 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2657 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_1945 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2813 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_6_3165 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_3007 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2993 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_wb_dat_gates\[28\]_B max_length1310/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_26_2381 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_2857 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_3465 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1649 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_52_4333 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_3329 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_193 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_4355 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_3621 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_52_4377 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1373 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_3752 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_4339 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1905 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3941 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_52_2997 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_3985 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__206__A _206_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_11_3384 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_3425 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xmax_length1311 _294_/X vssd vccd max_length1311/X vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_11_2683 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_49_1113 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_3469 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_20_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire2081_A wire2081/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_28_3881 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XANTENNA_input164_A la_iena_mprj[13] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_20_97 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_wire2179_A wire2179/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput300 la_oenb_mprj[20] vssd vccd _517_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_1_977 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_wb_dat_gates\[19\]_B max_length1311/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput311 la_oenb_mprj[30] vssd vccd wire1572/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput322 la_oenb_mprj[40] vssd vccd _409_/A_N vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_22_4192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput333 la_oenb_mprj[50] vssd vccd _547_/A vssd vccd sky130_fd_sc_hd__buf_4
XANTENNA_input331_A la_oenb_mprj[49] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput344 la_oenb_mprj[60] vssd vccd _557_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_29_51 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_input429_A mprj_dat_o_core[17] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_2_3552 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput355 la_oenb_mprj[70] vssd vccd wire1547/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_2_4297 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput366 la_oenb_mprj[80] vssd vccd wire1537/A vssd vccd sky130_fd_sc_hd__buf_6
XANTENNA_input25_A la_data_out_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xinput377 la_oenb_mprj[90] vssd vccd _587_/A vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_48_469 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1633 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput388 mprj_adr_o_core[0] vssd vccd wire1526/A vssd vccd sky130_fd_sc_hd__buf_6
Xinput399 mprj_adr_o_core[1] vssd vccd wire1489/A vssd vccd sky130_fd_sc_hd__buf_6
XFILLER_18_4217 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA__595__B _595_/B vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_18_4239 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1677 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_16_333 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
X_595_ _595_/A _595_/B vssd vccd _595_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_31_4417 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_377 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_837 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2414 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_4313 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2447 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1161 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_4 mprj_ack_i_user vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput807 _561_/X vssd vccd la_oenb_core[64] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput818 _571_/X vssd vccd la_oenb_core[74] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_49_3093 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output550_A _432_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_10_2182 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput829 _581_/X vssd vccd la_oenb_core[84] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_6_77 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_3509 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_29_3689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
X_029_ _029_/A vssd vccd _029_/Y vssd vccd sky130_fd_sc_hd__inv_2
XFILLER_42_4557 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1219 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1279_A _311_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_4_793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_4197 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_281 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_3222 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__489__C _489_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XANTENNA_output815_A _568_/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_45_2289 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_20_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1446_A wire1446/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_23_2565 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_2576 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] _225_/X vssd vccd _045_/A vssd vccd
+ sky130_fd_sc_hd__nand2_4
XFILLER_23_2587 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_27_609 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1936 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3605 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_19_193 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_4041 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_36_3649 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_664 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_50_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_1337 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_826 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_17_2314 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_53_3963 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_34_4085 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_697 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_50_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1504 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_4350 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_52_1515 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA_wire1982_A wire1983/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_34_2672 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XANTENNA__026__A _026_/A vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_50_1261 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_1223 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_3745 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1868 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_3133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_4001 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_43_3609 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_8_3216 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1267 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_47_3789 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_4181 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2421 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_41_4045 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_2465 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA__399__C _399_/C vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_41_4089 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_44_1032 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_4573 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2261 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2114 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_2136 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1953 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2147 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_417 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_4548 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_19_3836 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_39_3273 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_2_1457 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_130 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_35_3137 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_380_ _508_/A _380_/B _380_/C vssd vccd _380_/X vssd vccd sky130_fd_sc_hd__and3b_1
XFILLER_40_133 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_329 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_177 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_30_3793 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input281_A la_oenb_mprj[119] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_33_1481 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_11_3192 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_input379_A la_oenb_mprj[92] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_2207 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_46_3277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_3531 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_4107 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_3772 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_4287 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3625 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_2429 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_3636 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_7_1313 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_262 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_3669 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
Xinput130 la_data_out_mprj[99] vssd vccd _468_/C vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_2_4072 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
Xinput141 la_iena_mprj[108] vssd vccd _271_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_7_1357 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_24_2874 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput152 la_iena_mprj[118] vssd vccd _281_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_2153 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
Xinput163 la_iena_mprj[12] vssd vccd _175_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
Xinput174 la_iena_mprj[22] vssd vccd _185_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_40_1441 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput185 la_iena_mprj[32] vssd vccd _195_/B vssd vccd sky130_fd_sc_hd__clkbuf_4
XFILLER_48_277 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xinput196 la_iena_mprj[42] vssd vccd _205_/B vssd vccd sky130_fd_sc_hd__buf_4
XFILLER_18_3302 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_4047 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_40_1485 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_37_3969 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_4361 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_1980 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_141 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_601 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_2623 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_18_3368 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_4225 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
X_578_ _578_/A _578_/B vssd vccd _578_/X vssd vccd sky130_fd_sc_hd__and2_4
XFILLER_16_185 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_53_1802 vssd vccd vssd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_2093 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_645 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_output598_A _089_/Y vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_31_4269 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_31_2801 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_2981 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_32_689 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XPHY_180 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XPHY_191 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XANTENNA_output765_A wire1026/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_51_1581 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1396_A wire1397/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
XFILLER_29_4165 vssd vccd vssd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_4007 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_12_2299 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_9_4248 vssd vccd vssd vccd sky130_fd_sc_hd__decap_6
XANTENNA_output932_A wire1162/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput604 _094_/Y vssd vccd la_data_in_mprj[111] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput615 _104_/Y vssd vccd la_data_in_mprj[121] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_44_3929 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_4321 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput626 _163_/Y vssd vccd la_data_in_mprj[16] vssd vccd sky130_fd_sc_hd__buf_8
Xoutput637 _009_/Y vssd vccd la_data_in_mprj[26] vssd vccd sky130_fd_sc_hd__buf_8
XANTENNA_wire1563_A _415_/A_N vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
Xoutput648 _019_/Y vssd vccd la_data_in_mprj[36] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_28_1005 vssd vccd vssd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_3497 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xoutput659 _029_/Y vssd vccd la_data_in_mprj[46] vssd vccd sky130_fd_sc_hd__buf_8
XFILLER_42_4365 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_25_2605 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2053 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_28_1049 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_42_2941 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XFILLER_45_2097 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
XANTENNA_wire1730_A wire1731/X vssd vccd vccd vssd sky130_fd_sc_hd__diode_2
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VPWR VNB VPB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=1e+06u
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=5.88e+06u area=6.072e+11p
.ends

.subckt xres_buf A X VPWR VGND LVPWR LVGND
XFILLER_0_24 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_16 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XANTENNA_lvlshiftdown_A A VGND VPWR VPWR VGND sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
Xlvlshiftdown A VGND VPWR X VGND VPWR LVPWR sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_0_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
.ends

* Black-box entry subcircuit for user_analog_project_wrapper abstract view
.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
.ends

.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VPWR Q VNB VPB
X0 a_1178_261# a_1028_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_1028_413# a_1598_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1178_261# a_1028_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X4 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1136_413# a_193_47# a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X10 VGND a_1598_47# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X14 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_1224_47# a_27_47# a_1028_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1028_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1296_47# a_1178_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_1028_413# a_1598_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR a_1598_47# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 a_1028_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VPWR a_1178_261# a_1136_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 Q a_1598_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X36 Q a_1598_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 VPWR SET_B a_1028_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_33_199# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_33_199# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_27_47# a_33_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_109_47# a_33_199# a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VPWR X VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VPWR Y VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_47# C a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y A a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_277_47# B a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VPWR X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VPWR X VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_4 A B VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_8 A B VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VPWR X VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_4 A B C VGND VPWR X VNB VPB
X0 VPWR A a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_294_47# B a_185_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_185_47# A a_94_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C a_294_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_94_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C a_94_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_94_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_94_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_94_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_94_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VPWR X VNB VPB
X0 a_297_47# a_27_47# a_193_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_369_47# B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR D a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_193_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND D a_469_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_193_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR B a_193_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_193_413# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_193_413# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_469_47# C a_369_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VPWR X VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VPWR X VNB VPB
X0 VPWR A1 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_926_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A3 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_926_297# A2 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_102_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_496_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_102_21# B1 a_496_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_102_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_102_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_672_297# A3 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_496_47# B1 a_102_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_102_21# A3 a_672_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND a_102_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_102_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_496_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR B1 a_102_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_496_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_672_297# A2 a_926_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VPWR X VNB VPB
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VPWR Y VNB VPB
X0 a_316_297# C1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_420_297# B1 a_316_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A1 a_420_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_568_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_420_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_217_297# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_568_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VPWR X VNB VPB
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VPWR X VNB VPB
X0 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# A0 a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1259_199# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_1302_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_792_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1259_199# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND a_1259_199# a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 a_79_21# A1 a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_79_21# A0 a_1302_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR S a_792_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_792_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1302_47# a_1259_199# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 VPWR a_1259_199# a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_1302_297# a_1259_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_792_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X27 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_1302_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND S a_792_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X30 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_79_21# A1 a_1302_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 a_792_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_75_199# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_208_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_315_47# A2 a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B1 a_75_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_75_199# A1 a_315_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_75_199# C1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_544_297# B1 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_75_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_201_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_201_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_201_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_75_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VPWR X VNB VPB
X0 a_77_199# B2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_323_297# A2 a_227_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_227_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_227_47# B1 a_77_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_77_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B1 a_539_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_227_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_77_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_77_199# A3 a_323_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_227_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_227_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_539_297# B2 a_77_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VPWR Y VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VPWR Y VNB VPB
X0 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_215_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VPWR Y VNB VPB
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VPWR X VNB VPB
X0 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_475_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_762_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_475_47# B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_80_21# A2 a_762_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_80_21# B1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_475_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A1 a_934_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_934_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A1 a_475_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 Y A1 a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_181_47# A2 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_109_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VPWR Y VNB VPB
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_41_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR a_41_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_316_47# C a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_41_93# a_423_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_423_47# B a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A_N a_41_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VPWR Y VNB VPB
X0 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_633_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VPWR X VNB VPB
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VPWR Y VNB VPB
X0 a_281_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_475_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y D a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_475_297# C a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_281_297# C a_475_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_297# B a_281_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VPWR X VNB VPB
X0 a_585_47# B1 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A2 a_266_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_81_21# C1 a_585_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_266_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_368_297# A2 a_266_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_266_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_266_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_81_21# A3 a_368_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_81_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 VPWR a_86_235# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_86_235# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_86_235# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_86_235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_715_47# A1 a_86_235# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND A2 a_715_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_499_297# C1 a_427_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_86_235# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_86_235# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_607_297# B1 a_499_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_427_297# D1 a_86_235# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_607_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_607_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VPWR Y VNB VPB
X0 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_991_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_633_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND D a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_215_47# B a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_633_47# C a_991_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X29 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_991_47# C a_633_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VPWR Y VNB VPB
X0 Y A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_641_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_109_297# B1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_277_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_109_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A3 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_641_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_277_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_109_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y C1 a_641_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VPWR X VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 a_27_47# B1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_47# A2 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_717_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_277_297# B2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# B2 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_277_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_277_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_277_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR C1 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_27_47# C1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_27_47# B2 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A1 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_277_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_277_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR B1 a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A1 a_717_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_109_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_717_297# A2 a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_109_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VPWR X VNB VPB
X0 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR A1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_473_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND C1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_79_204# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_473_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_473_297# B1 a_727_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_79_204# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND B1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_79_204# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_1123_47# A1 a_79_204# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_555_297# B1 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A2 a_473_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A2 a_1123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_951_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR a_79_204# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_79_204# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_79_204# A1 a_951_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_79_204# C1 a_555_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_727_297# C1 a_79_204# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 X a_79_204# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VPWR X VNB VPB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VPWR X VNB VPB
X0 VGND A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND B2 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_804_297# B1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_79_21# A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_445_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_804_297# C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_445_297# B1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_1053_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_79_21# C1 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_1053_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 a_804_297# B2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_79_21# B1 a_1053_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_79_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_445_297# B2 a_804_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_445_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_445_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR A2 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VPWR A1 a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VPWR X VNB VPB
X0 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_815_47# B a_701_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR C a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_174_21# a_27_47# a_815_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_701_47# C a_617_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_174_21# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_174_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR a_27_47# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_617_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VPWR Y VNB VPB
X0 VGND a_91_199# Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_91_199# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_245_297# B a_161_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_91_199# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_161_297# a_91_199# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VPWR Y VNB VPB
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_449_297# C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VPWR Y VNB VPB
X0 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_462_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y B1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_28_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_28_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 VGND A2 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 VPWR A2 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_28_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_462_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 VPWR A1 a_28_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VPWR X VNB VPB
X0 VGND B1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_741_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_84_21# A1 a_741_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_901_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_483_297# B1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_84_21# B1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_483_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A1 a_483_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 a_84_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_483_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_901_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VPWR Y VNB VPB
X0 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# A2 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 Y B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_445_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_27_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 a_27_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y A1 a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_445_47# A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X28 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VPWR A3 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 VGND A3 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VPWR X VNB VPB
X0 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND D a_304_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_198_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_304_47# C a_198_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VPWR X VNB VPB
X0 a_30_297# C1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND C1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_44_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 X a_44_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_477_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_285_297# B1 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND D1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 a_770_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_30_297# D1 a_44_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A2 a_770_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 a_44_47# D1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_477_297# B1 a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_770_47# A1 a_44_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 a_477_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR a_44_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_285_297# C1 a_30_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_44_47# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_44_47# A1 a_770_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 VGND a_44_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 VPWR A2 a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 X a_44_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_44_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_6 A VGND VPWR Y VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VPWR Y VNB VPB
X0 a_465_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_204_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y B1 a_204_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_109_297# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VPWR X VNB VPB
X0 a_174_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_174_21# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_476_47# a_27_47# a_174_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_174_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_174_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_548_47# a_505_280# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 X a_174_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR D a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND D a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_505_280# a_174_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_505_280# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND a_174_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_505_280# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_639_47# C a_548_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt housekeeping VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1] irq[2]
+ mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13] mask_rev_in[14]
+ mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18] mask_rev_in[19]
+ mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23] mask_rev_in[24]
+ mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28] mask_rev_in[29]
+ mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4] mask_rev_in[5]
+ mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0] mgmt_gpio_in[10]
+ mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14] mgmt_gpio_in[15]
+ mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19] mgmt_gpio_in[1]
+ mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23] mgmt_gpio_in[24]
+ mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28] mgmt_gpio_in[29]
+ mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32] mgmt_gpio_in[33]
+ mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37] mgmt_gpio_in[3]
+ mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7] mgmt_gpio_in[8]
+ mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11] mgmt_gpio_oeb[12]
+ mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16] mgmt_gpio_oeb[17]
+ mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20] mgmt_gpio_oeb[21]
+ mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25] mgmt_gpio_oeb[26]
+ mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2] mgmt_gpio_oeb[30]
+ mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34] mgmt_gpio_oeb[35]
+ mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4] mgmt_gpio_oeb[5]
+ mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9] mgmt_gpio_out[0]
+ mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13] mgmt_gpio_out[14]
+ mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18] mgmt_gpio_out[19]
+ mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22] mgmt_gpio_out[23]
+ mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27] mgmt_gpio_out[28]
+ mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31] mgmt_gpio_out[32]
+ mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36] mgmt_gpio_out[37]
+ mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6] mgmt_gpio_out[7]
+ mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb pad_flash_csb
+ pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb pad_flash_io0_oeb
+ pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb pll90_sel[0]
+ pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1] pll_div[2]
+ pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0] pll_trim[10]
+ pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16] pll_trim[17]
+ pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22] pll_trim[23]
+ pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5] pll_trim[6]
+ pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2]
+ pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1 serial_data_2
+ serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb
+ spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i VGND
XFILLER_39_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_350 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6914_ _7081_/CLK _6914_/D fanout478/X VGND VPWR _6914_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_82_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6845_ _6951_/CLK _6845_/D fanout474/X VGND VPWR _6845_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6776_ _6777_/CLK _6776_/D fanout483/X VGND VPWR _7195_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3988_ hold151/X hold99/X _3989_/S VGND VPWR _3988_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5727_ _6909_/Q _5814_/B1 _5724_/X _5726_/X VGND VPWR _5727_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_148_352 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5658_ _5664_/A _5658_/B _5666_/B VGND VPWR _5658_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_191_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4609_ _4607_/A _4753_/B VGND VPWR _4609_/Y VGND VPWR sky130_fd_sc_hd__nand2b_2
XFILLER_190_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5589_ _7098_/Q _7097_/Q VGND VPWR _5979_/A VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_2_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold340 _4055_/X VGND VPWR _6491_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold351 _6463_/Q VGND VPWR hold351/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _4236_/X VGND VPWR _6628_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _6718_/Q VGND VPWR hold373/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _4108_/X VGND VPWR _6523_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _7196_/A VGND VPWR hold395/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _4061_/X VGND VPWR _6494_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 hold1577/X VGND VPWR _5172_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _5383_/X VGND VPWR _6938_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1073 _6611_/Q VGND VPWR _4211_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1084 _5485_/X VGND VPWR _7029_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 _6516_/Q VGND VPWR _4099_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 _5652_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_23 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4960_ _4947_/C _4959_/Y _5018_/A _4775_/B VGND VPWR _5088_/D VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_51_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3911_ _3164_/Y _7158_/Q _3868_/S _3911_/B1 VGND VPWR _3911_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_17_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4891_ _4810_/A _4947_/C _4902_/B _4490_/B _4878_/C VGND VPWR _5029_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_177_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6630_ _6632_/CLK _6630_/D fanout454/X VGND VPWR _6630_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3842_ _3866_/S VGND VPWR _3851_/C VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_20_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6561_ _6653_/CLK _6561_/D fanout452/X VGND VPWR _6561_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_192_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3773_ _3773_/A _3773_/B _3773_/C VGND VPWR _3794_/A VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_118_503 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_514 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5512_ hold145/X hold99/X _5513_/S VGND VPWR _5512_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6492_ _6527_/CLK hold90/X fanout484/X VGND VPWR _7183_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_145_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5443_ hold928/X _5548_/A1 _5444_/S VGND VPWR _5443_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5374_ _5374_/A0 _5524_/A1 _5381_/S VGND VPWR _5374_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7113_ _7113_/CLK _7113_/D fanout459/X VGND VPWR _7113_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4325_ hold431/X _5544_/A1 _4327_/S VGND VPWR _4325_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7044_ _7069_/CLK hold78/X fanout482/X VGND VPWR _7044_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4256_ _4256_/A _4322_/B VGND VPWR _4261_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_3207_ _6917_/Q VGND VPWR _3207_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4187_ _6638_/Q _6307_/B VGND VPWR _4195_/S VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_95_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_762 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6828_ _6908_/CLK _6828_/D fanout475/X VGND VPWR _6828_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6759_ _6953_/CLK _6759_/D fanout459/X VGND VPWR _6759_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_148_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold170 _7174_/A VGND VPWR hold170/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 _5297_/X VGND VPWR _6862_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold192 _6559_/Q VGND VPWR hold192/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_311 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4110_ _4110_/A0 _5473_/A1 hold38/X VGND VPWR _4110_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5090_ _4672_/B _4496_/Y _4542_/B VGND VPWR _5090_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_96_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4041_ hold968/X _6355_/A1 _4043_/S VGND VPWR _4041_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_578 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5992_ _6818_/Q _5953_/X _5960_/X _7071_/Q _5991_/X VGND VPWR _5992_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4943_ _4673_/A _4619_/Y _4995_/B _4941_/X _5071_/A VGND VPWR _4944_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_178_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4874_ _4542_/A _4947_/B _4652_/Y _4694_/Y _4873_/X VGND VPWR _4875_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6613_ _6654_/CLK _6613_/D fanout454/X VGND VPWR _6613_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_20_434 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3825_ _6874_/Q _5310_/A _5229_/A _6802_/Q _3824_/X VGND VPWR _3826_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6544_ _6709_/CLK _6544_/D fanout445/X VGND VPWR _6544_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3756_ _7064_/Q _5523_/A _4286_/A _6681_/Q VGND VPWR _3756_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_9_490 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clkbuf_3_5_0_csclk/A VGND VPWR clkbuf_3_5_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
X_6475_ _6707_/CLK _6475_/D fanout445/X VGND VPWR _6475_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_118_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3687_ _6662_/Q _4262_/A _3684_/X _3686_/X VGND VPWR _3688_/C VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_133_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5426_ hold700/X _5513_/A1 _5426_/S VGND VPWR _5426_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput220 _7183_/X VGND VPWR mgmt_gpio_out[18] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput231 _7193_/X VGND VPWR mgmt_gpio_out[28] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput242 _7175_/X VGND VPWR mgmt_gpio_out[3] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput253 _3948_/Y VGND VPWR pad_flash_io0_oeb VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput264 _6739_/Q VGND VPWR pll_div[2] VGND VPWR sky130_fd_sc_hd__buf_12
X_5357_ hold305/X _5465_/A1 _5363_/S VGND VPWR _5357_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput275 _6431_/Q VGND VPWR pll_trim[13] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput286 _6425_/Q VGND VPWR pll_trim[23] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput297 _6751_/Q VGND VPWR pwr_ctrl_out[0] VGND VPWR sky130_fd_sc_hd__buf_12
X_4308_ hold748/X _6356_/A1 _4309_/S VGND VPWR _4308_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5288_ hold459/X _5528_/A1 _5291_/S VGND VPWR _5288_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7027_ _7085_/CLK _7027_/D fanout477/X VGND VPWR _7027_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4239_ _4239_/A0 _6353_/A1 _4243_/S VGND VPWR _4239_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_718 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xwire347 _3437_/Y VGND VPWR _3447_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_149_491 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire358 _3392_/Y VGND VPWR _3410_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_137_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout480 fanout485/X VGND VPWR fanout480/X VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_93_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3610_ _6909_/Q _5346_/A _4102_/A input64/X _3609_/X VGND VPWR _3611_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4590_ _4591_/A _4664_/B VGND VPWR _4747_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_3541_ _6854_/Q _5283_/A _5319_/A _6886_/Q _3540_/X VGND VPWR _3552_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold906 _6976_/Q VGND VPWR hold906/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold917 _5296_/X VGND VPWR _6861_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 _6992_/Q VGND VPWR hold928/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold939 _5530_/X VGND VPWR _7069_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6260_ _6633_/Q _5946_/X _5955_/X _6553_/Q VGND VPWR _6260_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3472_ _3472_/A _3472_/B _3472_/C VGND VPWR _3485_/A VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_143_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5211_ _5211_/A hold17/X VGND VPWR hold18/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6191_ _6650_/Q _5973_/A _5948_/X _6695_/Q _6190_/X VGND VPWR _6191_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5142_ _5142_/A _5142_/B _5142_/C _5142_/D VGND VPWR _5142_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_96_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5073_ _5073_/A _5073_/B _5073_/C VGND VPWR _5074_/C VGND VPWR sky130_fd_sc_hd__and3_1
X_4024_ hold351/X _5494_/A1 _4025_/S VGND VPWR _4024_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_65_662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5975_ _5975_/A _5975_/B _5975_/C _5975_/D VGND VPWR _5975_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_4926_ _4992_/A _4926_/B VGND VPWR _5068_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_52_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4857_ _4810_/A _4496_/Y _4856_/Y _4887_/A VGND VPWR _4878_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_193_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3808_ _6938_/Q _5382_/A _4304_/A _6695_/Q VGND VPWR _3808_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_176_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4788_ _4689_/A _4616_/Y _4658_/C VGND VPWR _5106_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_181_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6527_ _6527_/CLK _6527_/D fanout484/X VGND VPWR _6527_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_180_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3739_ input15/X _3381_/Y _5148_/A _6738_/Q _3738_/X VGND VPWR _3742_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6458_ _6747_/CLK _6458_/D fanout448/X VGND VPWR _6458_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5409_ _5409_/A hold17/X VGND VPWR _5417_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_121_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6389_ _6400_/A _6400_/B VGND VPWR _6389_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_48_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_618 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_464 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5760_ _6991_/Q _5627_/X _5635_/X _6831_/Q VGND VPWR _5760_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4711_ _4701_/Y _4710_/Y _4627_/A VGND VPWR _4711_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_148_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5691_ _5681_/Y _5690_/Y _6787_/Q _5652_/Y VGND VPWR _5691_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4642_ _4642_/A _4673_/B VGND VPWR _4644_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_162_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4573_ _4965_/B _4724_/A VGND VPWR _5041_/B VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold703 _5289_/X VGND VPWR _6855_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _6824_/Q VGND VPWR hold714/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6312_ _6312_/A0 _6312_/A1 _6315_/S VGND VPWR _7137_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3524_ _3562_/A _3546_/A VGND VPWR _4202_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_116_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold725 _4296_/X VGND VPWR _6688_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold736 _6568_/Q VGND VPWR hold736/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _5255_/X VGND VPWR _6825_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _6543_/Q VGND VPWR hold758/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 _6356_/X VGND VPWR _7154_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6562_/Q _5953_/X _5960_/X _6672_/Q _6242_/X VGND VPWR _6243_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3455_ _3455_/A _3577_/B VGND VPWR _4102_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_103_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6174_ _7062_/Q _5954_/X _5976_/D _6881_/Q _6156_/X VGND VPWR _6175_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3386_ _7017_/Q _5463_/A _3370_/Y _7009_/Q VGND VPWR _3386_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_97_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5125_ _4413_/Y _4946_/X _5124_/X _4823_/X VGND VPWR _5126_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_111_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1403 _6798_/Q VGND VPWR _5225_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1414 _6572_/Q VGND VPWR hold1414/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 _6583_/Q VGND VPWR hold1425/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1436 _7138_/Q VGND VPWR _6313_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _6595_/Q VGND VPWR _4192_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _5089_/B _5089_/C _5142_/A _5056_/D VGND VPWR _5058_/D VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1458 _6729_/Q VGND VPWR _3702_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _6573_/Q VGND VPWR _4167_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4007_ hold744/X _5540_/A1 _4007_/S VGND VPWR _4007_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A VGND VPWR clkbuf_2_1_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_53_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_698 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5958_ _5968_/A _5981_/A _5979_/C VGND VPWR _5958_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_52_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4909_ _4969_/A _5051_/B VGND VPWR _4909_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_5889_ _6458_/Q _5645_/X _5646_/X _6653_/Q _5888_/X VGND VPWR _5896_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_csclk clkbuf_2_3_0_csclk/A VGND VPWR clkbuf_3_5_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_136_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold30 hold30/A VGND VPWR hold30/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold53/X VGND VPWR hold54/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A VGND VPWR hold52/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A VGND VPWR hold63/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A VGND VPWR hold74/X VGND VPWR sky130_fd_sc_hd__buf_12
Xhold85 hold85/A VGND VPWR hold85/X VGND VPWR sky130_fd_sc_hd__buf_12
Xhold96 hold96/A VGND VPWR hold96/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_676 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_5 _5310_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3240_ _6415_/Q _3264_/B VGND VPWR _3867_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_140_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3171_ _6487_/Q VGND VPWR _3837_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_13_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6930_ _7006_/CLK _6930_/D fanout457/X VGND VPWR _6930_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_82_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6861_ _6951_/CLK _6861_/D fanout474/X VGND VPWR _6861_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_6_csclk clkbuf_3_1_0_csclk/X VGND VPWR _7036_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5812_ _7001_/Q _5643_/X _5664_/X _6929_/Q VGND VPWR _5812_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_6792_ _7054_/CLK _6792_/D fanout461/X VGND VPWR _6792_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_34_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5743_ _6902_/Q _5621_/X _5658_/X _6886_/Q VGND VPWR _5743_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_188_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5674_ _6963_/Q _5642_/X _5928_/A2 _6835_/Q _5673_/X VGND VPWR _5681_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4625_ _4625_/A _4625_/B VGND VPWR _4969_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_128_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold500 _4260_/X VGND VPWR _6658_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _6807_/Q VGND VPWR hold511/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _4556_/A _4562_/A _4972_/A VGND VPWR _4557_/A VGND VPWR sky130_fd_sc_hd__and3_1
Xhold522 _5434_/X VGND VPWR _6984_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _6479_/Q VGND VPWR hold533/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _3573_/A _3571_/B VGND VPWR _4292_/A VGND VPWR sky130_fd_sc_hd__nor2_2
Xhold544 _5525_/X VGND VPWR _7064_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold555 _6539_/Q VGND VPWR hold555/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _7155_/Q VGND VPWR hold566/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _4561_/B _4993_/A VGND VPWR _4582_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold577 _5408_/X VGND VPWR _6961_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold588 _7027_/Q VGND VPWR hold588/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ _6221_/X _6226_/B _6226_/C _6226_/D VGND VPWR _6226_/X VGND VPWR sky130_fd_sc_hd__and4b_1
Xhold599 _5509_/X VGND VPWR _7050_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3438_ _7069_/Q _5523_/A _5328_/A _6896_/Q VGND VPWR _3438_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_103_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6157_ _6929_/Q _5938_/X _5952_/X _6961_/Q VGND VPWR _6157_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_58_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1200 _5410_/X VGND VPWR _6962_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3369_ _3373_/B hold75/X VGND VPWR _5463_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1211 _7010_/Q VGND VPWR _5464_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1222 _5437_/X VGND VPWR _6986_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5108_ _5108_/A _5108_/B _5108_/C VGND VPWR _5135_/B VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1233 _7079_/Q VGND VPWR _5542_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 _4257_/X VGND VPWR _6655_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6982_/Q _5945_/X _5975_/C _6838_/Q _6087_/X VGND VPWR _6089_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1255 _6645_/Q VGND VPWR _4245_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _4215_/X VGND VPWR _6614_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1277 _6742_/Q VGND VPWR _5155_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _5039_/A _5039_/B _5039_/C _5039_/D VGND VPWR _5122_/A VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1288 _4009_/X VGND VPWR _6450_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _6737_/Q VGND VPWR _5149_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_618 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput120 wb_adr_i[29] VGND VPWR _3900_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VPWR _3899_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_dat_i[19] VGND VPWR _6333_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_dat_i[29] VGND VPWR _6338_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VPWR input164/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_48_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_679 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4410_ _4498_/A _4459_/B VGND VPWR _4948_/A VGND VPWR sky130_fd_sc_hd__nand2_4
X_5390_ hold658/X _5513_/A1 _5390_/S VGND VPWR _5390_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4341_ _4753_/A _4607_/A VGND VPWR _4690_/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_98_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7060_ _7078_/CLK hold88/X fanout482/X VGND VPWR _7060_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_99_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4272_ hold355/X _5494_/A1 _4273_/S VGND VPWR _4272_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6011_ _6971_/Q _5947_/X _5965_/X _6795_/Q _6010_/X VGND VPWR _6014_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_3223_ _6543_/Q VGND VPWR _3223_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_100_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6913_ _6969_/CLK _6913_/D fanout475/X VGND VPWR _6913_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6844_ _6884_/CLK _6844_/D fanout475/X VGND VPWR _6844_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_112 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6775_ _6777_/CLK hold92/X fanout483/X VGND VPWR hold91/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3987_ hold630/X _5469_/A1 _3989_/S VGND VPWR _3987_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5726_ _6901_/Q _5621_/X _5648_/X _6853_/Q _5725_/X VGND VPWR _5726_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5657_ _5664_/A _5657_/B _5660_/C VGND VPWR _5657_/X VGND VPWR sky130_fd_sc_hd__and3b_2
XFILLER_175_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4608_ _4607_/A _4753_/B VGND VPWR _4608_/X VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_163_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5588_ _6508_/Q _7098_/Q _7097_/Q VGND VPWR _5594_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_151_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold330 _5336_/X VGND VPWR _6897_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold341 _6785_/Q VGND VPWR hold341/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _4591_/A _4552_/A _4549_/A VGND VPWR _4959_/B VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_2_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold352 _4024_/X VGND VPWR _6463_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_123 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold363 _6948_/Q VGND VPWR hold363/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _4332_/X VGND VPWR _6718_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold385 _6996_/Q VGND VPWR hold385/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _5201_/X VGND VPWR _6777_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _6556_/Q _5971_/B _5949_/X _6676_/Q _6208_/X VGND VPWR _6225_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7189_ _7189_/A VGND VPWR _7189_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_100_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1030 _4028_/X VGND VPWR _6466_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _6780_/Q VGND VPWR _5205_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_362 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1052 _5172_/X VGND VPWR _6755_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_684 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1063 _6893_/Q VGND VPWR _5332_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 _4211_/X VGND VPWR _6611_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _7021_/Q VGND VPWR _5476_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1096 _4099_/X VGND VPWR _6516_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_203 _5667_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_96 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6926_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_64_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3910_ _3910_/A _3910_/B VGND VPWR _6635_/D VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_32_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4890_ _4542_/A _4496_/Y _4892_/B _4381_/Y _4697_/Y VGND VPWR _4895_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_3841_ _3837_/B _3867_/B _3840_/X _3860_/B VGND VPWR _3866_/S VGND VPWR sky130_fd_sc_hd__o31a_4
XFILLER_32_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6560_ _6653_/CLK _6560_/D fanout452/X VGND VPWR _6560_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3772_ _6540_/Q _4127_/A _3769_/X _3771_/X VGND VPWR _3773_/C VGND VPWR sky130_fd_sc_hd__a211o_1
X_5511_ hold403/X _5538_/A1 _5513_/S VGND VPWR _5511_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6491_ _6527_/CLK _6491_/D fanout484/X VGND VPWR _7182_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_157_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5442_ hold379/X _5538_/A1 _5444_/S VGND VPWR _5442_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_173_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5373_ _5373_/A hold17/X VGND VPWR _5381_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7112_ _7131_/CLK _7112_/D fanout459/X VGND VPWR _7112_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4324_ hold265/X _5534_/A1 _4327_/S VGND VPWR _4324_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7043_ _7079_/CLK _7043_/D fanout478/X VGND VPWR _7043_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4255_ _4255_/A0 hold60/X _4255_/S VGND VPWR _4255_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3206_ _6925_/Q VGND VPWR _3206_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4186_ _3410_/Y _4186_/A1 _4186_/S VGND VPWR _6590_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk _6888_/CLK VGND VPWR _6969_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xclkbuf_3_1_0_csclk clkbuf_3_1_0_csclk/A VGND VPWR clkbuf_3_1_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_82_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_546 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_387 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_590 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6827_ _6884_/CLK _6827_/D fanout475/X VGND VPWR _6827_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_51_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6758_ _6953_/CLK _6758_/D fanout460/X VGND VPWR _6758_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_183_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5709_ _6948_/Q _5637_/X _5660_/X _6804_/Q VGND VPWR _5709_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_149_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6689_ _6707_/CLK _6689_/D fanout448/X VGND VPWR _6689_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_12_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold160 _6863_/Q VGND VPWR hold160/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _4074_/X VGND VPWR _6500_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _7043_/Q VGND VPWR hold182/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold193 _4150_/X VGND VPWR _6559_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_43 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_323 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_175 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4040_ hold796/X _6354_/A1 _4043_/S VGND VPWR _4040_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5991_ _7010_/Q _5940_/X _5947_/X _6970_/Q _5990_/X VGND VPWR _5991_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_18_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4942_ _4942_/A _4942_/B _4942_/C VGND VPWR _5071_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_178_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4873_ _4542_/A _4496_/Y _4700_/Y _4627_/B _4872_/X VGND VPWR _4873_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_757 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6612_ _6671_/CLK _6612_/D _6383_/A VGND VPWR _6612_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3824_ _6768_/Q _5190_/A _5190_/B _4274_/A _6670_/Q VGND VPWR _3824_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_6543_ _6735_/CLK _6543_/D fanout445/X VGND VPWR _6543_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3755_ _6427_/Q _3981_/A _4220_/A _6620_/Q _3754_/X VGND VPWR _3760_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6474_ _6735_/CLK _6474_/D _3946_/B VGND VPWR _6474_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3686_ _6996_/Q _5445_/A _5211_/A _6788_/Q _3685_/X VGND VPWR _3686_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_118_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput210 _3216_/Y VGND VPWR mgmt_gpio_oeb[7] VGND VPWR sky130_fd_sc_hd__buf_12
X_5425_ hold906/X _5548_/A1 _5426_/S VGND VPWR _5425_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput221 _7184_/X VGND VPWR mgmt_gpio_out[19] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput232 _7194_/X VGND VPWR mgmt_gpio_out[29] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput243 _7176_/X VGND VPWR mgmt_gpio_out[4] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput254 _7198_/X VGND VPWR pad_flash_io1_do VGND VPWR sky130_fd_sc_hd__buf_12
X_5356_ _5356_/A0 hold667/X _5363_/S VGND VPWR _5356_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput265 _6740_/Q VGND VPWR pll_div[3] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput276 _6432_/Q VGND VPWR pll_trim[14] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6748_/Q VGND VPWR pll_trim[24] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_101_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput298 _6752_/Q VGND VPWR pwr_ctrl_out[1] VGND VPWR sky130_fd_sc_hd__buf_12
X_4307_ hold956/X _6355_/A1 _4309_/S VGND VPWR _4307_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5287_ hold912/X _5509_/A1 _5291_/S VGND VPWR _5287_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7026_ _7026_/CLK _7026_/D fanout465/X VGND VPWR _7026_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4238_ _4238_/A _4322_/B VGND VPWR _4243_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_87_479 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4169_ _3486_/Y _4169_/A1 _4171_/S VGND VPWR _6575_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_74_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire348 _3826_/Y VGND VPWR _3827_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_136_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_554 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout470 _6390_/A VGND VPWR fanout470/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_48_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout481 fanout485/X VGND VPWR fanout481/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_171_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3540_ _6918_/Q _5355_/A _6352_/A _7155_/Q VGND VPWR _3540_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_128_665 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold907 _5425_/X VGND VPWR _6976_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _6880_/Q VGND VPWR hold918/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold929 _5443_/X VGND VPWR _6992_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3471_ _6943_/Q _5382_/A _5274_/A _6847_/Q _3457_/X VGND VPWR _3472_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_182_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5210_ hold341/X _5540_/A1 _5210_/S VGND VPWR _5210_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_143_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6190_ _6645_/Q _5976_/C _5971_/D _6565_/Q VGND VPWR _6190_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5141_ _4542_/A _4946_/X _5058_/C _5140_/X VGND VPWR _5142_/D VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_96_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5072_ _4565_/X _4741_/A _4650_/Y _5088_/C VGND VPWR _5073_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_96_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4023_ _4023_/A0 _6355_/A1 _4025_/S VGND VPWR _4023_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5974_ _5946_/X _5970_/X _5974_/C _5974_/D VGND VPWR _5977_/A VGND VPWR sky130_fd_sc_hd__and4bb_1
XFILLER_40_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4925_ _5088_/A _4925_/B _5114_/A VGND VPWR _5103_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_21_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4856_ _4856_/A _4911_/B VGND VPWR _4856_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_3807_ _3807_/A _3807_/B _3807_/C _3807_/D VGND VPWR _3827_/B VGND VPWR sky130_fd_sc_hd__nor4_1
X_4787_ _4644_/Y _4714_/X _4782_/Y VGND VPWR _4791_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_20_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6526_ _6527_/CLK hold7/X fanout484/X VGND VPWR _6526_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3738_ _6651_/Q _4250_/A _4133_/A _6546_/Q VGND VPWR _3738_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_109_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6457_ _6747_/CLK _6457_/D fanout447/X VGND VPWR _6457_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3669_ _6940_/Q _5382_/A _4172_/A _6580_/Q _3668_/X VGND VPWR _3670_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5408_ hold576/X _5513_/A1 _5408_/S VGND VPWR _5408_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6388_ _6400_/A _6400_/B VGND VPWR _6388_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_133_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5339_ hold618/X _5543_/A1 _5345_/S VGND VPWR _5339_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_125_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7009_ _7017_/CLK _7009_/D fanout461/X VGND VPWR _7009_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_75_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_302 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_471 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_722 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_131 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4710_ _4710_/A _4969_/B VGND VPWR _4710_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_5690_ _5690_/A _5690_/B _5690_/C _5690_/D VGND VPWR _5690_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_187_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4641_ _4739_/A _4661_/B VGND VPWR _4673_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_147_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4572_ _4672_/A _4947_/B VGND VPWR _4574_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_116_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold704 _6839_/Q VGND VPWR hold704/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ _3640_/Y _6311_/A1 _6315_/S VGND VPWR _7136_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold715 _5254_/X VGND VPWR _6824_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ _3523_/A _3523_/B _3523_/C _3523_/D VGND VPWR _3582_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_155_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold726 _6999_/Q VGND VPWR hold726/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold737 _4161_/X VGND VPWR _6568_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_763 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold748 _6698_/Q VGND VPWR hold748/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 _4131_/X VGND VPWR _6543_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _6652_/Q _5973_/A _5948_/X _6697_/Q _6241_/X VGND VPWR _6242_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3454_ _3454_/A _3454_/B VGND VPWR _3577_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_115_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6173_ _6817_/Q _5971_/B _5949_/X _6937_/Q _6172_/X VGND VPWR _6175_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3385_ _6945_/Q _5382_/A _5436_/A _6993_/Q VGND VPWR _3385_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5124_ _4672_/B _4496_/Y _4810_/A VGND VPWR _5124_/X VGND VPWR sky130_fd_sc_hd__a21o_1
Xhold1404 _6469_/Q VGND VPWR _4031_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1415 _6573_/Q VGND VPWR hold1415/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1426 _6584_/Q VGND VPWR hold1426/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _6592_/Q VGND VPWR _4189_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _4413_/Y _4496_/Y _5092_/B _5054_/X VGND VPWR _5056_/D VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_57_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1448 _7137_/Q VGND VPWR _6312_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _6732_/Q VGND VPWR _3488_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ hold892/X _5548_/A1 _4007_/S VGND VPWR _4006_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5957_ _5969_/A _5968_/A _5969_/C VGND VPWR _5975_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_178_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4908_ _4845_/X _4907_/X _4465_/B VGND VPWR _4915_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_166_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5888_ _7154_/Q _5625_/X _5642_/X _6718_/Q VGND VPWR _5888_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4839_ _5068_/A _4964_/B _5039_/C _4838_/X _4541_/X VGND VPWR _4839_/X VGND VPWR
+ sky130_fd_sc_hd__a41o_1
XFILLER_166_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6509_ _7131_/CLK _6509_/D fanout460/X VGND VPWR _6509_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_134_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_340 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3224__1 net399_2/A VGND VPWR _7157_/CLK VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_76_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold20 hold20/A VGND VPWR hold20/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold31 hold31/A VGND VPWR hold31/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VPWR hold42/X VGND VPWR sky130_fd_sc_hd__buf_8
Xhold53 hold53/A VGND VPWR hold53/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A VGND VPWR hold64/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A VGND VPWR hold75/X VGND VPWR sky130_fd_sc_hd__buf_8
Xhold86 hold86/A VGND VPWR hold86/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A VGND VPWR hold97/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_688 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_708 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _5310_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_153_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3170_ _6635_/Q VGND VPWR _3170_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6860_ _7079_/CLK _6860_/D fanout478/X VGND VPWR _6860_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_179_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5811_ _6937_/Q _5654_/X _5808_/X _5809_/X _5810_/X VGND VPWR _5811_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_179_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6791_ _6953_/CLK _6791_/D fanout459/X VGND VPWR _6791_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5742_ _6870_/Q _5628_/X _5634_/X _6974_/Q _5741_/X VGND VPWR _5748_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5673_ _6947_/Q _5637_/X _5638_/X _6955_/Q VGND VPWR _5673_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4624_ _4620_/Y _4645_/B VGND VPWR _4942_/B VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_163_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold501 _6602_/Q VGND VPWR hold501/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4555_ _4724_/A _4650_/A VGND VPWR _5088_/C VGND VPWR sky130_fd_sc_hd__nand2_2
Xhold512 _5235_/X VGND VPWR _6807_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _6441_/Q VGND VPWR hold523/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _4043_/X VGND VPWR _6479_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _6747_/Q VGND VPWR hold545/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3506_ _3554_/A _3692_/A VGND VPWR _4250_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_1_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold556 _4126_/X VGND VPWR _6539_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ _4690_/B _4626_/B VGND VPWR _4689_/A VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold567 _6357_/X VGND VPWR _7155_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _6699_/Q VGND VPWR hold578/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold589 _5483_/X VGND VPWR _7027_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ _6225_/A _6225_/B _6225_/C _6225_/D VGND VPWR _6225_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_3437_ _6912_/Q _5346_/A _3432_/X _3434_/X _3436_/X VGND VPWR _3437_/Y VGND VPWR
+ sky130_fd_sc_hd__a2111oi_1
X_6156_ _7086_/Q _5976_/B _5971_/C _7046_/Q VGND VPWR _6156_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3368_ _3543_/A hold85/X VGND VPWR _5373_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1201 _6786_/Q VGND VPWR _5212_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _5464_/X VGND VPWR _7010_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 _6954_/Q VGND VPWR _5401_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5107_ _4611_/Y _4644_/Y _4663_/Y _4969_/Y VGND VPWR _5108_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_57_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1234 _5542_/X VGND VPWR _7079_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3299_ _3347_/A hold72/X VGND VPWR _3311_/C VGND VPWR sky130_fd_sc_hd__nor2_2
X_6087_ _6926_/Q _5938_/X _5952_/X _6958_/Q VGND VPWR _6087_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_73_706 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1245 _6660_/Q VGND VPWR _4263_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _4245_/X VGND VPWR _6645_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 _6890_/Q VGND VPWR _5329_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _5155_/X VGND VPWR _6742_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _5114_/B _5115_/A _5038_/C VGND VPWR _5038_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_73_739 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1289 _6675_/Q VGND VPWR _4281_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6989_ _7082_/CLK _6989_/D fanout480/X VGND VPWR _6989_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_41_647 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_371 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput110 wb_adr_i[1] VGND VPWR _4556_/A VGND VPWR sky130_fd_sc_hd__buf_8
Xinput121 wb_adr_i[2] VGND VPWR _4625_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput132 wb_dat_i[0] VGND VPWR _6323_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput143 wb_dat_i[1] VGND VPWR _6327_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_544 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VPWR _6329_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VPWR _6316_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_63_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_173 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4340_ _4753_/A _4607_/A VGND VPWR _4562_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_153_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4271_ _4271_/A0 _6355_/A1 _4273_/S VGND VPWR _4271_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3222_ _6789_/Q VGND VPWR _3222_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_97_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6010_ _6891_/Q _5946_/X _5955_/X _6803_/Q VGND VPWR _6010_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_79_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6912_ _6951_/CLK _6912_/D fanout474/X VGND VPWR _6912_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_35_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6843_ _7067_/CLK _6843_/D fanout477/X VGND VPWR _6843_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_62_271 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6774_ _7082_/CLK _6774_/D fanout483/X VGND VPWR _7193_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3986_ hold620/X _6357_/A1 _3989_/S VGND VPWR _3986_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5725_ _6869_/Q _5628_/X _5658_/X _6885_/Q VGND VPWR _5725_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_148_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5656_ _6930_/Q _5654_/X _5655_/X _6794_/Q _5653_/X VGND VPWR _5669_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4607_ _4607_/A _4970_/A VGND VPWR _4673_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_5587_ _7098_/Q _7097_/Q VGND VPWR _5968_/A VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_117_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold320 _5521_/X VGND VPWR _7061_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _6905_/Q VGND VPWR hold331/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4538_ _4424_/Y _4500_/Y _4504_/X _4537_/Y _5023_/A VGND VPWR _4538_/X VGND VPWR
+ sky130_fd_sc_hd__o41a_1
XFILLER_116_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold342 _5210_/X VGND VPWR _6785_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold353 _7012_/Q VGND VPWR hold353/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold364 _5394_/X VGND VPWR _6948_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _6515_/Q VGND VPWR hold375/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_135 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold386 _5448_/X VGND VPWR _6996_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4469_ _4469_/A _4672_/A VGND VPWR _4472_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold397 _7078_/Q VGND VPWR hold397/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _7035_/Q _5601_/X _5959_/X _6716_/Q VGND VPWR _6208_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7188_ _7188_/A VGND VPWR _7188_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6139_ _6984_/Q _5945_/X _5975_/C _6840_/Q _6138_/X VGND VPWR _6140_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1020 _4135_/X VGND VPWR _6546_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1031 _6451_/Q VGND VPWR _4010_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _5205_/X VGND VPWR _6780_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1053 _6447_/Q VGND VPWR _4005_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_374 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_78 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1064 _5332_/X VGND VPWR _6893_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1075 _6909_/Q VGND VPWR _5350_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _5476_/X VGND VPWR _7021_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 _6949_/Q VGND VPWR _5395_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _5971_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_45_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_744 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_csclk clkbuf_3_1_0_csclk/X VGND VPWR _6632_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_174_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3840_ _7167_/Q _3875_/C _6485_/Q VGND VPWR _3840_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_20_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_499 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3771_ _6794_/Q _3326_/Y _4032_/A _6470_/Q _3770_/X VGND VPWR _3771_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_157_140 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5510_ hold483/X _5528_/A1 _5513_/S VGND VPWR _5510_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6490_ _6527_/CLK _6490_/D fanout481/X VGND VPWR _7181_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5441_ hold439/X _5528_/A1 _5444_/S VGND VPWR _5441_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5372_ hold654/X _5513_/A1 _5372_/S VGND VPWR _5372_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7111_ _7131_/CLK _7111_/D fanout459/X VGND VPWR _7111_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4323_ _4323_/A0 hold667/X _4327_/S VGND VPWR _4323_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7086_/CLK _7042_/D fanout483/X VGND VPWR _7042_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4254_ hold389/X _5494_/A1 _4255_/S VGND VPWR _4254_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3205_ _6933_/Q VGND VPWR _3205_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4185_ _3447_/Y _4185_/A1 _4186_/S VGND VPWR _6589_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_399 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6826_ _6908_/CLK _6826_/D fanout475/X VGND VPWR _6826_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_50_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6757_ _6953_/CLK _6757_/D fanout460/X VGND VPWR _6757_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3969_ hold1/X hold4/X _3975_/S VGND VPWR hold5/A VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_109_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_460 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5708_ _6836_/Q _5928_/A2 _5697_/X _5707_/X VGND VPWR _5711_/B VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_164_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_516 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6688_ _6707_/CLK _6688_/D fanout448/X VGND VPWR _6688_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5639_ _6946_/Q _5637_/X _5638_/X _6954_/Q _5636_/X VGND VPWR _5639_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_136_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold150 _5389_/X VGND VPWR _6944_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _5298_/X VGND VPWR _6863_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _7148_/Q VGND VPWR hold172/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold183 _5501_/X VGND VPWR _7043_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _6678_/Q VGND VPWR hold194/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_688 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_699 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5990_ _6938_/Q _5961_/X _5976_/D _6874_/Q VGND VPWR _5990_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_91_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4941_ _4996_/C _4941_/B _5073_/B _4941_/D VGND VPWR _4941_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_17_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4872_ _4872_/A _4872_/B _4872_/C _4872_/D VGND VPWR _4872_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_20_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6611_ _6668_/CLK _6611_/D fanout452/X VGND VPWR _6611_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3823_ _6655_/Q _4256_/A _4172_/A _6578_/Q _3822_/X VGND VPWR _3826_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6542_ _6709_/CLK _6542_/D fanout445/X VGND VPWR _6542_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_118_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3754_ _6811_/Q _5238_/A hold67/A _6466_/Q VGND VPWR _3754_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6473_ _6704_/CLK _6473_/D fanout448/X VGND VPWR _6473_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3685_ _6852_/Q _5283_/A _4208_/A _6611_/Q VGND VPWR _3685_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5424_ hold882/X _5538_/A1 _5426_/S VGND VPWR _5424_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput200 _3191_/Y VGND VPWR mgmt_gpio_oeb[32] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput211 _3215_/Y VGND VPWR mgmt_gpio_oeb[8] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput222 _3932_/X VGND VPWR mgmt_gpio_out[1] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput233 _7174_/X VGND VPWR mgmt_gpio_out[2] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput244 _7177_/X VGND VPWR mgmt_gpio_out[5] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5355_ _5355_/A _5541_/B VGND VPWR _5363_/S VGND VPWR sky130_fd_sc_hd__and2_4
Xoutput255 _3950_/A VGND VPWR pad_flash_io1_ieb VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput266 _6741_/Q VGND VPWR pll_div[4] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput277 _6433_/Q VGND VPWR pll_trim[15] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput288 _6749_/Q VGND VPWR pll_trim[25] VGND VPWR sky130_fd_sc_hd__buf_12
X_4306_ hold818/X _6354_/A1 _4309_/S VGND VPWR _4306_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput299 _6753_/Q VGND VPWR pwr_ctrl_out[2] VGND VPWR sky130_fd_sc_hd__buf_12
X_5286_ hold333/X _5526_/A1 _5291_/S VGND VPWR _5286_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7025_ _7086_/CLK hold31/X fanout484/X VGND VPWR _7025_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4237_ hold842/X _5546_/A1 _4237_/S VGND VPWR _4237_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4168_ _6312_/A0 _4168_/A1 _4171_/S VGND VPWR _6574_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_558 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4099_ _4099_/A0 _4098_/X _4101_/S VGND VPWR _4099_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_539 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_583 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6809_ _7078_/CLK _6809_/D fanout481/X VGND VPWR _6809_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_184_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire349 _3670_/Y VGND VPWR _3699_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_136_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VPWR _7037_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_151_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_566 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout460 fanout462/X VGND VPWR fanout460/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout471 _6396_/A VGND VPWR _6390_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout482 fanout485/X VGND VPWR fanout482/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_46_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_753 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6884_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_30_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk _6888_/CLK VGND VPWR _7070_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_155_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_677 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold908 _6808_/Q VGND VPWR hold908/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold919 _5317_/X VGND VPWR _6880_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ _6839_/Q _5265_/A _5463_/A _7015_/Q _3458_/X VGND VPWR _3472_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5140_ _4542_/D _4672_/B _4518_/C _4821_/X VGND VPWR _5140_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_170_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5071_ _5071_/A _5071_/B _5071_/C VGND VPWR _5077_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_84_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4022_ _4022_/A0 _5492_/A1 _4025_/S VGND VPWR _4022_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_111_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5973_ _5973_/A _5973_/B VGND VPWR _5974_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_80_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4924_ _4456_/Y _4562_/Y _4673_/A _4689_/B _4768_/C VGND VPWR _4999_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4855_ _4782_/A _4630_/X _4515_/Y VGND VPWR _4855_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3806_ _6680_/Q _4286_/A _3585_/Y input98/X _3805_/X VGND VPWR _3807_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4786_ _4673_/A _4689_/B _4781_/X _5108_/B _4785_/X VGND VPWR _4791_/A VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_165_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6525_ _6527_/CLK _6525_/D fanout484/X VGND VPWR _6525_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3737_ _7048_/Q _5505_/A _5274_/A _6843_/Q _3736_/X VGND VPWR _3742_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_180_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6456_ _6704_/CLK _6456_/D fanout447/X VGND VPWR _6456_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3668_ _6462_/Q _4020_/A _4328_/A _6717_/Q VGND VPWR _3668_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_173_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5407_ hold137/X hold99/X _5408_/S VGND VPWR _5407_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6387_ _6401_/A _6401_/B VGND VPWR _6387_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_88_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3599_ _6683_/Q _4286_/A _4268_/A _6668_/Q _3598_/X VGND VPWR _3604_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5338_ _5338_/A0 hold667/X _5345_/S VGND VPWR _5338_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_544 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5269_ hold223/X _5494_/A1 _5273_/S VGND VPWR _5269_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_75_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7008_ _7033_/CLK _7008_/D fanout464/X VGND VPWR _7008_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_56_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_314 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_647 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_658 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_439 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_678 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4640_ _4673_/A _4626_/Y _4639_/Y VGND VPWR _5062_/A VGND VPWR sky130_fd_sc_hd__a21o_1
X_4571_ _4496_/Y _4570_/Y _5099_/A _4559_/X _4548_/X VGND VPWR _4589_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_6310_ _3700_/Y _6310_/A1 _6315_/S VGND VPWR _7135_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_116_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold705 _5271_/X VGND VPWR _6839_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3522_ _6838_/Q _5265_/A _3381_/Y input30/X _3521_/X VGND VPWR _3523_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold716 _6872_/Q VGND VPWR hold716/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 _5451_/X VGND VPWR _6999_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold738 _6873_/Q VGND VPWR hold738/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold749 _4308_/X VGND VPWR _6698_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _6647_/Q _5976_/C _5971_/D _6567_/Q VGND VPWR _6241_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3453_ _3453_/A hold64/X _3454_/A VGND VPWR _5164_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_131_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6172_ _6449_/Q _5601_/X _5959_/X _6969_/Q VGND VPWR _6172_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3384_ _7033_/Q hold49/A _5505_/A _7054_/Q VGND VPWR _3384_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5123_ _5123_/A VGND VPWR _5123_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xhold1405 _6963_/Q VGND VPWR _5411_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _6575_/Q VGND VPWR hold1416/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 _6588_/Q VGND VPWR hold1427/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1438 _6594_/Q VGND VPWR _4191_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _4413_/Y _4672_/B _5057_/A _5057_/B VGND VPWR _5054_/X VGND VPWR sky130_fd_sc_hd__o211a_1
Xhold1449 _6722_/Q VGND VPWR _4988_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ _4005_/A0 _5469_/A1 _4007_/S VGND VPWR _4005_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_65_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5956_ _5978_/A _5964_/A _5969_/C VGND VPWR _5976_/C VGND VPWR sky130_fd_sc_hd__and3_4
X_4907_ _4887_/B _4907_/B VGND VPWR _4907_/X VGND VPWR sky130_fd_sc_hd__and2b_1
X_5887_ _5887_/A1 _6279_/S _5885_/X _5886_/X VGND VPWR _7116_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_21_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4838_ _4453_/B _4570_/Y _4837_/X _4925_/B VGND VPWR _4838_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_119_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_708 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4769_ _4769_/A _4999_/A _4769_/C _4769_/D VGND VPWR _4770_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_181_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6508_ _7113_/CLK _6508_/D fanout460/X VGND VPWR _6508_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_119_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6439_ _6747_/CLK _6439_/D fanout447/X VGND VPWR _6439_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_134_488 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold10/A VGND VPWR hold10/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_352 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold21 hold21/A VGND VPWR hold21/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VPWR hold32/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold43 hold43/A VGND VPWR hold43/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A VGND VPWR hold54/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A VGND VPWR hold65/X VGND VPWR sky130_fd_sc_hd__buf_6
Xhold76 hold76/A VGND VPWR hold76/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A VGND VPWR hold87/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A VGND VPWR hold98/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_7 _5391_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_556 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5810_ _6873_/Q _5628_/X _5658_/X _6889_/Q _5801_/X VGND VPWR _5810_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_6790_ _7006_/CLK _6790_/D fanout457/X VGND VPWR _6790_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5741_ _6982_/Q _5624_/X _5654_/X _6934_/Q VGND VPWR _5741_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5672_ _5672_/A1 _6103_/B1 _5670_/Y _5671_/X VGND VPWR _7106_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_175_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4623_ _4653_/B _4638_/A VGND VPWR _4623_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_136_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4554_ _4574_/A _4554_/B VGND VPWR _4559_/B VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold502 _4200_/X VGND VPWR _6602_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold513 _6871_/Q VGND VPWR hold513/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _3998_/X VGND VPWR _6441_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ hold74/X _3562_/B VGND VPWR _4044_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold535 _6883_/Q VGND VPWR hold535/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_606 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold546 _5160_/X VGND VPWR _6747_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4485_ _4690_/B _4626_/B VGND VPWR _4911_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold557 hold557/A VGND VPWR hold557/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _6926_/Q VGND VPWR hold568/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold579 _4309_/X VGND VPWR _6699_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6456_/Q _5944_/X _5975_/A _6600_/Q _6205_/X VGND VPWR _6225_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3436_ _7000_/Q _5445_/A _3964_/A _6424_/Q _3435_/X VGND VPWR _3436_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_131_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6155_ _7033_/Q _5944_/X _5975_/A _6849_/Q VGND VPWR _6155_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3367_ _3370_/A _3511_/A VGND VPWR _3367_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_85_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1202 _5212_/X VGND VPWR _6786_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5106_ _5106_/A _5106_/B _5106_/C _5106_/D VGND VPWR _5109_/B VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1213 _6994_/Q VGND VPWR _5446_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1224 _5401_/X VGND VPWR _6954_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6086_ _6974_/Q _5947_/X _5965_/X _6798_/Q _6085_/X VGND VPWR _6089_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1235 _6619_/Q VGND VPWR _4221_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3298_ _3975_/S hold71/X _3298_/B1 VGND VPWR _3298_/Y VGND VPWR sky130_fd_sc_hd__o21ai_2
XFILLER_57_247 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1246 _4263_/X VGND VPWR _6660_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _6475_/Q VGND VPWR _4039_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5114_/C _5086_/C _5037_/C _5115_/B VGND VPWR _5038_/C VGND VPWR sky130_fd_sc_hd__nand4_1
Xhold1268 _5329_/X VGND VPWR _6890_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 _6460_/Q VGND VPWR _4021_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6988_ _7049_/CLK _6988_/D fanout456/X VGND VPWR _6988_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_53_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_659 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5939_ _7098_/Q _7097_/Q VGND VPWR _5981_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_178_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_547 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_700 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_704 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput100 wb_adr_i[10] VGND VPWR _4337_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput111 wb_adr_i[20] VGND VPWR _4566_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput122 wb_adr_i[30] VGND VPWR input122/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_103_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput133 wb_dat_i[10] VGND VPWR _6330_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VPWR _6336_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VPWR _6341_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_sel_i[1] VGND VPWR _6319_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_76_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_718 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_152 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4270_ _4270_/A0 _5492_/A1 _4273_/S VGND VPWR _4270_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3221_ _6797_/Q VGND VPWR _3221_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_121_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6911_ _6967_/CLK _6911_/D fanout474/X VGND VPWR _6911_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6842_ _7026_/CLK _6842_/D fanout463/X VGND VPWR _6842_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_35_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6773_ _6777_/CLK _6773_/D fanout479/X VGND VPWR _7192_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3985_ hold770/X _6356_/A1 _3989_/S VGND VPWR _3985_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5724_ _6997_/Q _5643_/X _5667_/X _6813_/Q VGND VPWR _5724_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_50_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5655_ _5638_/A _5667_/C _5666_/C VGND VPWR _5655_/X VGND VPWR sky130_fd_sc_hd__and3b_4
X_4606_ _4607_/A _4970_/A VGND VPWR _4975_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_5586_ _5586_/A VGND VPWR _7097_/D VGND VPWR sky130_fd_sc_hd__inv_2
Xhold310 _4224_/X VGND VPWR _6622_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold321 _6964_/Q VGND VPWR hold321/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _5068_/A _4925_/B _4537_/C _4537_/D VGND VPWR _4537_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_132_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold332 _5345_/X VGND VPWR _6905_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 _7004_/Q VGND VPWR hold343/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold354 _5466_/X VGND VPWR _7012_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _7195_/A VGND VPWR hold365/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _4817_/A _4965_/B VGND VPWR _5041_/A VGND VPWR sky130_fd_sc_hd__nand2_2
Xhold376 _4097_/X VGND VPWR _6515_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _6956_/Q VGND VPWR hold387/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold398 _5540_/X VGND VPWR _7078_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _7152_/Q _5958_/X _5978_/X _6481_/Q VGND VPWR _6207_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_89_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3419_ _6808_/Q _5229_/A hold86/A _7061_/Q VGND VPWR _3419_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_7187_ _7187_/A VGND VPWR _7187_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4399_ _4551_/A _4813_/A VGND VPWR _4459_/A VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_98_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6138_ _6928_/Q _5938_/X _5952_/X _6960_/Q VGND VPWR _6138_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_58_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1010 _4252_/X VGND VPWR _6651_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _6600_/Q VGND VPWR _4198_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1032 _4010_/X VGND VPWR _6451_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 _6499_/Q VGND VPWR _4072_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1054 _4005_/X VGND VPWR _6447_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6069_ _6821_/Q _5953_/X _5960_/X _7074_/Q _6068_/X VGND VPWR _6069_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1065 _7013_/Q VGND VPWR _5467_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1076 _5350_/X VGND VPWR _6909_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 _6989_/Q VGND VPWR _5440_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 _5395_/X VGND VPWR _6949_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _3251_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_54_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3770_ _7010_/Q _5463_/A _4316_/A _6705_/Q VGND VPWR _3770_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_157_152 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5440_ _5440_/A0 _5545_/A1 _5444_/S VGND VPWR _5440_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_66_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5371_ hold114/X hold99/X _5372_/S VGND VPWR _5371_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7110_ _7131_/CLK _7110_/D fanout456/X VGND VPWR _7110_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4322_ _4322_/A _4322_/B VGND VPWR _4327_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_7041_ _7051_/CLK hold3/X fanout477/X VGND VPWR _7041_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4253_ hold888/X _5493_/A1 _4255_/S VGND VPWR _4253_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3204_ _6941_/Q VGND VPWR _3204_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_79_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4184_ _3486_/Y _4184_/A1 _4186_/S VGND VPWR _6588_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_353 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VPWR _3937_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_6825_ _7070_/CLK _6825_/D fanout473/X VGND VPWR _6825_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_168_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6756_ _6769_/CLK _6756_/D fanout469/X VGND VPWR _7173_/A VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3968_ hold247/X _5465_/A1 _3980_/S VGND VPWR _3968_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_149_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5707_ _6844_/Q _5902_/A2 _5905_/A2 _6796_/Q _5695_/X VGND VPWR _5707_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6687_ _6707_/CLK _6687_/D fanout448/X VGND VPWR _6687_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_176_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3899_ input123/X input122/X _3899_/C _3899_/D VGND VPWR _3901_/C VGND VPWR sky130_fd_sc_hd__and4bb_1
XFILLER_164_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_528 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5638_ _5638_/A _5657_/B _5666_/C VGND VPWR _5638_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_117_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5569_ _6508_/Q _5567_/Y _7092_/Q VGND VPWR _7092_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_151_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold140 _5218_/X VGND VPWR _6792_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A VGND VPWR hold151/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _6958_/Q VGND VPWR hold162/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _3979_/X VGND VPWR hold21/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _6902_/Q VGND VPWR hold184/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _4284_/X VGND VPWR _6678_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_288 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_397 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_20 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4940_ _4948_/B _4562_/Y _4673_/A _4644_/Y _4738_/Y VGND VPWR _4941_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4871_ _4947_/B _4456_/Y _4694_/Y _4627_/B VGND VPWR _4872_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_178_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6610_ _6668_/CLK _6610_/D _6400_/A VGND VPWR _6610_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3822_ _6604_/Q _4202_/A _4262_/A _6660_/Q VGND VPWR _3822_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_20_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6541_ _6709_/CLK _6541_/D fanout445/X VGND VPWR _6541_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_146_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3753_ _6915_/Q _5355_/A hold49/A _7027_/Q _3752_/X VGND VPWR _3760_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6472_ _6735_/CLK _6472_/D _3946_/B VGND VPWR _6472_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_173_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3684_ input54/X _5193_/A _5229_/A _6804_/Q VGND VPWR _3684_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5423_ hold437/X _5528_/A1 _5426_/S VGND VPWR _5423_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput201 _3190_/Y VGND VPWR mgmt_gpio_oeb[33] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput212 _3214_/Y VGND VPWR mgmt_gpio_oeb[9] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput223 _7185_/X VGND VPWR mgmt_gpio_out[20] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput234 _7195_/X VGND VPWR mgmt_gpio_out[30] VGND VPWR sky130_fd_sc_hd__buf_12
X_5354_ hold675/X _5540_/A1 _5354_/S VGND VPWR _5354_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput245 _3929_/X VGND VPWR mgmt_gpio_out[6] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput256 _3950_/Y VGND VPWR pad_flash_io1_oeb VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput267 _6735_/Q VGND VPWR pll_ena VGND VPWR sky130_fd_sc_hd__buf_12
X_4305_ _4305_/A0 _5491_/A1 _4309_/S VGND VPWR _4305_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput278 _6418_/Q VGND VPWR pll_trim[16] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_59_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput289 _6436_/Q VGND VPWR pll_trim[2] VGND VPWR sky130_fd_sc_hd__buf_12
X_5285_ hold293/X _5465_/A1 _5291_/S VGND VPWR _5285_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7024_ _7085_/CLK _7024_/D fanout482/X VGND VPWR _7024_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4236_ hold361/X _5518_/A1 _4237_/S VGND VPWR _4236_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4167_ _3640_/Y _4167_/A1 _4171_/S VGND VPWR _6573_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4098_ hold291/X _5548_/A1 _5202_/B VGND VPWR _4098_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_82_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_58 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_4_csclk clkbuf_leaf_4_csclk/A VGND VPWR _6654_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6808_ _7085_/CLK _6808_/D fanout482/X VGND VPWR _6808_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6739_ _6739_/CLK _6739_/D _3946_/B VGND VPWR _6739_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_136_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_636 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout450 fanout486/X VGND VPWR fanout450/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_171_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout461 fanout462/X VGND VPWR fanout461/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout472 fanout486/X VGND VPWR _6396_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_120_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout483 fanout484/X VGND VPWR fanout483/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_34_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_710 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_765 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_623 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold909 _5236_/X VGND VPWR _6808_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5070_ _4542_/B _4428_/Y _4846_/B _4619_/Y _4771_/C VGND VPWR _5071_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4021_ _4021_/A0 _6353_/A1 _4025_/S VGND VPWR _4021_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5972_ _5600_/A _5978_/A _5981_/B _5934_/X _5967_/X VGND VPWR _5973_/B VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_64_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4923_ _4921_/A _5043_/A _4747_/A _4747_/B _4740_/B VGND VPWR _4923_/Y VGND VPWR
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_178_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4854_ _4542_/B _4947_/B _4902_/B _4616_/Y VGND VPWR _4877_/B VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_60_381 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3805_ _6834_/Q _5265_/A _4328_/A _6715_/Q VGND VPWR _3805_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4785_ _4902_/B _4689_/B _4784_/X _4967_/A VGND VPWR _4785_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_118_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6524_ _6527_/CLK _6524_/D fanout484/X VGND VPWR _6524_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3736_ _6676_/Q _4280_/A _4139_/A _6551_/Q VGND VPWR _3736_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_119_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6455_ _6747_/CLK _6455_/D fanout447/X VGND VPWR _6455_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3667_ _7012_/Q _5463_/A _5182_/S _6759_/Q _3666_/X VGND VPWR _3670_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_659 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5406_ hold710/X _5469_/A1 _5408_/S VGND VPWR _5406_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6386_ _6401_/A _6400_/B VGND VPWR _6386_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_133_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3598_ input46/X hold37/A _5523_/A _7066_/Q VGND VPWR _3598_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_133_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5337_ _5337_/A _5541_/B VGND VPWR _5345_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_735 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5268_ hold369/X _5526_/A1 _5273_/S VGND VPWR _5268_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_556 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7007_ _7017_/CLK _7007_/D fanout461/X VGND VPWR _7007_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4219_ hold982/X _5546_/A1 _4219_/S VGND VPWR _4219_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_75_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5199_ hold91/X hold42/X _5201_/S VGND VPWR hold92/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4570_ _4570_/A _4959_/B VGND VPWR _4570_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_3521_ _7083_/Q _5541_/A _4172_/A _6582_/Q VGND VPWR _3521_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold706 _6927_/Q VGND VPWR hold706/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 _5308_/X VGND VPWR _6872_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _6740_/Q VGND VPWR hold728/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ _6240_/A _6240_/B _6240_/C VGND VPWR _6240_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_143_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold739 _5309_/X VGND VPWR _6873_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ _3714_/B _3562_/B VGND VPWR _5154_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_115_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6171_ _7025_/Q _5937_/X _5975_/D _6889_/Q _6155_/X VGND VPWR _6175_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3383_ _7025_/Q hold29/A _5409_/A _6969_/Q VGND VPWR _3383_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_124_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_532 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5122_ _5122_/A _5122_/B _5122_/C VGND VPWR _5123_/A VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1406 _5411_/X VGND VPWR hold14/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1417 _7160_/Q VGND VPWR hold8/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _4948_/A _4672_/B _4523_/Y _4824_/X _4953_/Y VGND VPWR _5092_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
Xhold1428 _6589_/Q VGND VPWR hold1428/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1439 _6593_/Q VGND VPWR _4190_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4004_ hold79/X _5519_/A1 _4007_/S VGND VPWR hold80/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5955_ _5978_/A _5981_/B _5969_/C VGND VPWR _5955_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4906_ _4381_/Y _4900_/Y _4869_/B VGND VPWR _4906_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5886_ _5552_/B _7115_/Q _6103_/B1 VGND VPWR _5886_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_139_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4837_ _5114_/A _5089_/A _5018_/A _4837_/D VGND VPWR _4837_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_4768_ _4768_/A _4768_/B _4768_/C _4768_/D VGND VPWR _4769_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_147_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6507_ _7131_/CLK _6507_/D fanout460/X VGND VPWR _6507_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3719_ _6443_/Q _3999_/A _5145_/A _6736_/Q _3718_/X VGND VPWR _3720_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4699_ _4460_/A _4611_/B _4628_/Y _4967_/B _4625_/A VGND VPWR _4706_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_134_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6438_ _6747_/CLK _6438_/D fanout447/X VGND VPWR _6438_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_88_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6369_ _6383_/A _6396_/B VGND VPWR _6369_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_96_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_csclk clkbuf_opt_2_0_csclk/X VGND VPWR _6882_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold11 hold11/A VGND VPWR hold11/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VPWR hold22/X VGND VPWR sky130_fd_sc_hd__buf_6
Xhold33 hold33/A VGND VPWR hold33/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A VGND VPWR hold44/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A VGND VPWR hold55/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VPWR hold66/X VGND VPWR sky130_fd_sc_hd__buf_8
Xhold77 hold77/A VGND VPWR hold77/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A VGND VPWR hold88/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VPWR hold99/X VGND VPWR sky130_fd_sc_hd__buf_12
Xclkbuf_leaf_37_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7078_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_90_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VPWR clkbuf_0_mgmt_gpio_in[4]/X VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XPHY_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 hold29/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_152_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_120 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_568 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5740_ _6990_/Q _5627_/X _5635_/X _6830_/Q VGND VPWR _5740_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_188_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5671_ _6786_/Q _5652_/Y _5610_/Y VGND VPWR _5671_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_175_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4622_ _4653_/B _4638_/A VGND VPWR _4645_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_4553_ _4947_/C _4553_/B VGND VPWR _4554_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_144_732 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold503 _7030_/Q VGND VPWR hold503/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold514 _5307_/X VGND VPWR _6871_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold525 _6649_/Q VGND VPWR hold525/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ _3504_/A _3504_/B _3504_/C _3504_/D VGND VPWR _3504_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
Xhold536 _5321_/X VGND VPWR _6883_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4562_/A _4972_/A VGND VPWR _4484_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold547 _7190_/A VGND VPWR hold547/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_618 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold558 _7048_/Q VGND VPWR hold558/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold569 _5369_/X VGND VPWR _6926_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6681_/Q _5934_/X _5975_/B _6615_/Q _6222_/X VGND VPWR _6225_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3435_ _6984_/Q _5427_/A _3381_/Y input32/X VGND VPWR _3435_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6154_ _6178_/A0 _6153_/X _6304_/S VGND VPWR _6154_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3366_ _3571_/A _3379_/A VGND VPWR _5274_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1203 _6930_/Q VGND VPWR _5374_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _4616_/Y _4970_/Y _5010_/Y _4613_/Y VGND VPWR _5106_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_57_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1214 _5446_/X VGND VPWR _6994_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6085_ _6894_/Q _5946_/X _5955_/X _6806_/Q VGND VPWR _6085_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold1225 _6751_/Q VGND VPWR _5167_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3297_ hold1003/X _3975_/S VGND VPWR _3297_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold1236 _4221_/X VGND VPWR _6619_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _6970_/Q VGND VPWR _5419_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _4500_/A _4902_/B _4494_/Y _4882_/C _4909_/Y VGND VPWR _5115_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_57_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_440 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1258 _4039_/X VGND VPWR _6475_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1269 _6630_/Q VGND VPWR _4239_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6987_ _7085_/CLK _6987_/D fanout477/X VGND VPWR _6987_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_41_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5938_ _5979_/A _5981_/A _5981_/B VGND VPWR _5938_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_179_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5869_ _6697_/Q _5637_/X _5645_/X _6457_/Q VGND VPWR _5869_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_166_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_716 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput101 wb_adr_i[11] VGND VPWR _4337_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput112 wb_adr_i[21] VGND VPWR _4702_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_76_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput123 wb_adr_i[31] VGND VPWR input123/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VPWR _6332_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_103_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput145 wb_dat_i[21] VGND VPWR _6339_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_dat_i[31] VGND VPWR _6344_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VPWR _6318_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3220_ _6805_/Q VGND VPWR _3220_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_67_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_708 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6910_ _7081_/CLK _6910_/D fanout478/X VGND VPWR _6910_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_47_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6841_ _6865_/CLK _6841_/D fanout464/X VGND VPWR _6841_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6772_ _7082_/CLK _6772_/D fanout479/X VGND VPWR _7191_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3984_ hold993/X _6355_/A1 _3989_/S VGND VPWR _3984_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5723_ _6981_/Q _5624_/X _5654_/X _6933_/Q _5717_/Y VGND VPWR _5723_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5654_ _5664_/A _5667_/C _5660_/C VGND VPWR _5654_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4605_ _4753_/A _4753_/B VGND VPWR _4625_/B VGND VPWR sky130_fd_sc_hd__nand2b_2
XFILLER_163_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5585_ _5567_/Y _6508_/Q _7097_/Q VGND VPWR _5586_/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold300 _5429_/X VGND VPWR _6979_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold311 _7046_/Q VGND VPWR hold311/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4536_ _5010_/A _4969_/A _4881_/B VGND VPWR _4537_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
Xhold322 _5412_/X VGND VPWR _6964_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _6852_/Q VGND VPWR hold333/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _5457_/X VGND VPWR _7004_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _6668_/Q VGND VPWR hold355/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _5200_/X VGND VPWR _6776_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4467_ _4498_/A _4531_/B _4579_/B VGND VPWR _5027_/A VGND VPWR sky130_fd_sc_hd__nand3_1
Xhold377 _6683_/Q VGND VPWR hold377/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold388 _5403_/X VGND VPWR _6956_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold399 _6940_/Q VGND VPWR hold399/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6610_/Q _5943_/X _5981_/X _6656_/Q VGND VPWR _6206_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3418_ _7053_/Q _5505_/A _3367_/Y input27/X VGND VPWR _3418_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7186_ _7186_/A VGND VPWR _7186_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4398_ _4415_/A _4415_/B VGND VPWR _4813_/A VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_98_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1000 _4173_/X VGND VPWR _6578_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6137_ _6976_/Q _5947_/X _5965_/X _6800_/Q _6136_/X VGND VPWR _6140_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3349_ hold75/A hold28/X VGND VPWR hold29/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1011 _6610_/Q VGND VPWR _4210_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1022 _4198_/X VGND VPWR _6600_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _6615_/Q VGND VPWR _4216_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _4072_/X VGND VPWR _6499_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6068_ _6909_/Q _5973_/A _5948_/X _6949_/Q _6067_/X VGND VPWR _6068_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1055 _7026_/Q VGND VPWR _5482_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1066 _5467_/X VGND VPWR _7013_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 _6842_/Q VGND VPWR _5275_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _5440_/X VGND VPWR _6989_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _5041_/B _4681_/Y _4710_/Y _4627_/A VGND VPWR _5021_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_26_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1099 _6802_/Q VGND VPWR _5230_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_206 _5490_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_273 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_744 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_418 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5370_ hold706/X _5469_/A1 _5372_/S VGND VPWR _5370_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4321_ hold580/X _6357_/A1 _4321_/S VGND VPWR _4321_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_245 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7040_ _7081_/CLK _7040_/D fanout477/X VGND VPWR _7040_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4252_ _4252_/A0 _5492_/A1 _4255_/S VGND VPWR _4252_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3203_ _6949_/Q VGND VPWR _3203_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_101_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4183_ _4192_/A0 _4183_/A1 _4186_/S VGND VPWR _6587_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_192 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6824_ _6920_/CLK _6824_/D fanout473/X VGND VPWR _6824_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6755_ _6755_/CLK _6755_/D _6360_/A VGND VPWR _6755_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3967_ hold8/X hold11/X _3975_/S VGND VPWR hold12/A VGND VPWR sky130_fd_sc_hd__mux2_8
X_5706_ _5706_/A _5706_/B _5706_/C _5706_/D VGND VPWR _5706_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
X_6686_ _6707_/CLK _6686_/D fanout448/X VGND VPWR _6686_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3898_ _4334_/B _4334_/C VGND VPWR _4702_/C VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_191_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5637_ _5664_/A _5658_/B _5657_/B VGND VPWR _5637_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_148_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5568_ _6506_/Q _5610_/B VGND VPWR _5568_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_117_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold130 _5180_/X VGND VPWR _6761_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _6856_/Q VGND VPWR hold141/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ _4886_/B _4953_/A VGND VPWR _4522_/B VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold152 _6998_/Q VGND VPWR hold152/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _5405_/X VGND VPWR _6958_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5499_/A0 hold6/X hold77/A VGND VPWR _5499_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold174 hold21/X VGND VPWR hold174/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _5342_/X VGND VPWR _6902_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _6814_/Q VGND VPWR hold196/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7169_ _3945_/A1 _7169_/D _6399_/X VGND VPWR _7169_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_86_674 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_32 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4870_ _4870_/A _5027_/B _4870_/C VGND VPWR _4872_/C VGND VPWR sky130_fd_sc_hd__and3_1
X_3821_ _6810_/Q _5238_/A _4208_/A _6609_/Q _3820_/X VGND VPWR _3826_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6540_ _6735_/CLK _6540_/D fanout445/X VGND VPWR _6540_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3752_ _6995_/Q _5445_/A _5373_/A _6931_/Q VGND VPWR _3752_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_146_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6471_ _6739_/CLK _6471_/D _3946_/B VGND VPWR _6471_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3683_ _6482_/Q _4044_/A _4268_/A _6667_/Q _3682_/X VGND VPWR _3688_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_173_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5422_ _5422_/A0 _5545_/A1 _5426_/S VGND VPWR _5422_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_173_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput202 _3189_/Y VGND VPWR mgmt_gpio_oeb[34] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_173_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput213 _3933_/X VGND VPWR mgmt_gpio_out[0] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput224 _7186_/X VGND VPWR mgmt_gpio_out[21] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput235 _7196_/X VGND VPWR mgmt_gpio_out[31] VGND VPWR sky130_fd_sc_hd__buf_12
X_5353_ hold673/X _5521_/A1 _5354_/S VGND VPWR _5353_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput246 _7178_/X VGND VPWR mgmt_gpio_out[7] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput257 _6745_/Q VGND VPWR pll90_sel[0] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput268 _6742_/Q VGND VPWR pll_sel[0] VGND VPWR sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A _6352_/B VGND VPWR _4309_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_87_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput279 _6419_/Q VGND VPWR pll_trim[17] VGND VPWR sky130_fd_sc_hd__buf_12
X_5284_ _5284_/A0 _5524_/A1 _5291_/S VGND VPWR _5284_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7023_ _7086_/CLK hold57/X fanout482/X VGND VPWR hold56/A VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_87_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4235_ hold461/X _5544_/A1 _4237_/S VGND VPWR _4235_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4166_ _3700_/Y _4166_/A1 _4171_/S VGND VPWR _6572_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_460 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4097_ hold375/X _4096_/X _4101_/S VGND VPWR _4097_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_82_176 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6807_ _7078_/CLK _6807_/D fanout481/X VGND VPWR _6807_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_11_416 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4999_ _4999_/A _4999_/B _4999_/C VGND VPWR _5001_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_6738_ _6739_/CLK _6738_/D _3946_/B VGND VPWR _6738_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_315 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6669_ _6677_/CLK _6669_/D fanout452/X VGND VPWR _6669_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_164_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_648 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout440 _6396_/B VGND VPWR _6400_/B VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout451 fanout452/X VGND VPWR _6400_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout462 fanout466/X VGND VPWR fanout462/X VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_59_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout473 fanout474/X VGND VPWR fanout473/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout484 fanout485/X VGND VPWR fanout484/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_74_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_292 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_703 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4020_ _4020_/A _5490_/B VGND VPWR _4025_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_49_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_614 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5971_ _5971_/A _5971_/B _5971_/C _5971_/D VGND VPWR _5974_/C VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_18_593 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_658 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4922_ _4582_/B _4576_/B _4737_/A _4965_/B VGND VPWR _4922_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_100_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4853_ _4947_/B _4948_/C _4902_/B _4689_/B VGND VPWR _4872_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_178_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3804_ _7055_/Q hold86/A _4157_/A _6565_/Q _3803_/X VGND VPWR _3807_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_4784_ _4625_/B _4702_/Y _4703_/Y _4716_/Y _4646_/Y VGND VPWR _4784_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
Xclkbuf_opt_2_0_csclk _6601_/CLK VGND VPWR clkbuf_opt_2_0_csclk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6523_ _6990_/CLK _6523_/D fanout478/X VGND VPWR _6523_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3735_ _6787_/Q _5211_/A _4151_/A _6561_/Q _3734_/X VGND VPWR _3742_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6454_ _6655_/CLK _6454_/D _6383_/A VGND VPWR _6454_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3666_ _6472_/Q _4032_/A _4322_/A _6712_/Q VGND VPWR _3666_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_106_318 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5405_ hold162/X hold60/X _5408_/S VGND VPWR _5405_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_161_435 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6385_ _6401_/A _6401_/B VGND VPWR _6385_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3597_ _6869_/Q _5301_/A _4250_/A _6653_/Q _3596_/X VGND VPWR _3597_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5336_ hold329/X _5540_/A1 _5336_/S VGND VPWR _5336_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_671 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5267_ hold297/X _5465_/A1 _5273_/S VGND VPWR _5267_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_568 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7006_ _7006_/CLK _7006_/D fanout458/X VGND VPWR _7006_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4218_ hold495/X _5518_/A1 _4219_/S VGND VPWR _4218_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5198_ hold443/X _5528_/A1 _5201_/S VGND VPWR _5198_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_324 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4149_ hold317/X _5518_/A1 _4150_/S VGND VPWR _4149_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_332 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_135 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3520_ _3562_/A _3577_/B VGND VPWR _4172_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_7_762 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold707 _5370_/X VGND VPWR _6927_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _6920_/Q VGND VPWR hold718/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _5152_/X VGND VPWR _6740_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3451_ _3454_/A hold84/X VGND VPWR _3562_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_41_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6170_ _7070_/Q _5934_/X _5975_/B _6873_/Q _6169_/X VGND VPWR _6175_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3382_ _6857_/Q _5283_/A _5427_/A _6985_/Q VGND VPWR _3382_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_130_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_csclk clkbuf_3_1_0_csclk/X VGND VPWR _6653_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_124_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5121_ _5087_/D _5118_/X _5120_/X _5116_/Y VGND VPWR _5129_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_57_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1407 _7150_/Q VGND VPWR _3963_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1418 _6597_/Q VGND VPWR hold1418/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _4551_/A _5041_/Y _4957_/Y VGND VPWR _5142_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_97_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1429 _6571_/Q VGND VPWR hold1429/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4003_ hold646/X _5509_/A1 _4007_/S VGND VPWR _4003_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_65_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5954_ _5978_/A _5966_/A _5981_/B VGND VPWR _5954_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4905_ _5080_/A _4905_/B _5131_/A VGND VPWR _4916_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_5885_ _6542_/Q _5652_/Y _5875_/X _5884_/X _6303_/S VGND VPWR _5885_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4836_ _4810_/A _4810_/B _4834_/X _4835_/Y _5088_/B VGND VPWR _4837_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_166_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4767_ _4764_/X _4767_/B _4767_/C _4996_/B VGND VPWR _4768_/D VGND VPWR sky130_fd_sc_hd__and4b_1
X_6506_ _7131_/CLK _6506_/D fanout459/X VGND VPWR _6506_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3718_ _6875_/Q _5310_/A _5463_/A _7011_/Q VGND VPWR _3718_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_4_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_273 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4698_ _4984_/A _4970_/A _4698_/C VGND VPWR _4967_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_107_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6437_ _7155_/CLK _6437_/D fanout449/X VGND VPWR _6437_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3649_ _7081_/Q _5541_/A _3999_/A _6444_/Q VGND VPWR _3649_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_134_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6368_ _6401_/A _6401_/B VGND VPWR _6368_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5319_ _5319_/A _5541_/B VGND VPWR _5327_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6299_ _6694_/Q _5954_/X _5976_/D _6623_/Q _6280_/X VGND VPWR _6300_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold12 hold12/A VGND VPWR hold9/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VPWR hold23/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold34 hold34/A VGND VPWR hold34/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold45 hold45/A VGND VPWR hold45/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A VGND VPWR hold56/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A VGND VPWR hold67/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A VGND VPWR hold78/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold89 hold89/A VGND VPWR hold89/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_90_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_379 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _5328_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_152_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5670_ _5670_/A _5670_/B VGND VPWR _5670_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_175_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4621_ _4846_/B _4616_/Y _4619_/Y _4673_/A VGND VPWR _4621_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_129_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4552_ _4552_/A _4664_/A VGND VPWR _4574_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_156_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold504 _5486_/X VGND VPWR _7030_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _6879_/Q VGND VPWR hold515/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _6862_/Q _5292_/A _5418_/A _6974_/Q _3502_/X VGND VPWR _3504_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4483_ _4984_/A _4636_/A VGND VPWR _4483_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xhold526 _4249_/X VGND VPWR _6649_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold537 _6803_/Q VGND VPWR hold537/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _5195_/X VGND VPWR _6771_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold559 _5507_/X VGND VPWR _7048_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ _6701_/Q _5971_/A _5979_/X _6471_/Q VGND VPWR _6222_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3434_ _6960_/Q _5400_/A _3999_/A _6448_/Q _3433_/X VGND VPWR _3434_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_171_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6153_ _7124_/Q _6152_/X _6303_/S VGND VPWR _6153_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3365_ _3373_/B _3511_/A VGND VPWR _3365_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
X_5104_ _5004_/A _5077_/A _5099_/X _5138_/B _5103_/Y VGND VPWR _5129_/D VGND VPWR
+ sky130_fd_sc_hd__a41o_1
Xhold1204 _5374_/X VGND VPWR _6930_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _6942_/Q _5961_/X _6080_/X _6083_/X VGND VPWR _6089_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_97_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1215 _6978_/Q VGND VPWR _5428_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3296_ _3292_/A hold70/X _6488_/Q VGND VPWR hold71/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1226 _5167_/X VGND VPWR _6751_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _6690_/Q VGND VPWR _4299_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _5419_/X VGND VPWR _6970_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _4899_/B _5118_/B _5083_/C _5035_/D VGND VPWR _5037_/C VGND VPWR sky130_fd_sc_hd__and4b_1
Xhold1259 _6510_/Q VGND VPWR _4087_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_452 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6986_ _7049_/CLK _6986_/D fanout457/X VGND VPWR _6986_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_41_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5937_ _5979_/A _5964_/A _5981_/A VGND VPWR _5937_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_15_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5868_ _6687_/Q _5632_/X _5638_/X _6707_/Q VGND VPWR _5868_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_139_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4819_ _4413_/Y _4902_/A _4562_/Y _4542_/B VGND VPWR _5057_/A VGND VPWR sky130_fd_sc_hd__o22a_1
X_5799_ _6507_/Q _7111_/Q _6103_/B1 VGND VPWR _5799_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_166_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput102 wb_adr_i[12] VGND VPWR _4336_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput113 wb_adr_i[22] VGND VPWR _4334_/C VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput124 wb_adr_i[3] VGND VPWR _4753_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_193_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput135 wb_dat_i[12] VGND VPWR _6335_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_dat_i[22] VGND VPWR _6342_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput157 wb_dat_i[3] VGND VPWR _6333_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_sel_i[3] VGND VPWR _6320_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_91_539 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6840_ _6997_/CLK _6840_/D fanout463/X VGND VPWR _6840_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6771_ _7082_/CLK _6771_/D fanout479/X VGND VPWR _7190_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3983_ hold828/X _6354_/A1 _3989_/S VGND VPWR _3983_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5722_ _7013_/Q _5630_/X _5719_/X _5720_/X _5721_/X VGND VPWR _5722_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6683_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5653_ _6850_/Q _5648_/X _5652_/B _6914_/Q _5651_/Y VGND VPWR _5653_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_694 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_508 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_154 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4604_ _4753_/A _4753_/B VGND VPWR _4970_/A VGND VPWR sky130_fd_sc_hd__and2b_2
X_5584_ _5584_/A VGND VPWR _7096_/D VGND VPWR sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7076_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold301 _6939_/Q VGND VPWR hold301/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4535_ _4535_/A _4535_/B _4535_/C _4535_/D VGND VPWR _4537_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_116_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold312 _5504_/X VGND VPWR _7046_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _7058_/Q VGND VPWR hold323/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _5286_/X VGND VPWR _6852_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _6693_/Q VGND VPWR hold345/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4466_ _4493_/B VGND VPWR _4846_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_104_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold356 _4272_/X VGND VPWR _6668_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold367 _6753_/Q VGND VPWR hold367/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _4290_/X VGND VPWR _6683_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold389 _6653_/Q VGND VPWR hold389/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6466_/Q _5937_/X _5975_/D _6626_/Q VGND VPWR _6205_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3417_ _7131_/Q _6761_/Q _6762_/Q VGND VPWR _3417_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_131_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7185_ _7185_/A VGND VPWR _7185_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4397_ _4739_/A _4396_/A _4400_/B VGND VPWR _4415_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_6136_ _6896_/Q _5946_/X _5955_/X _6808_/Q VGND VPWR _6136_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_58_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3348_ _3586_/A _3714_/B VGND VPWR _5211_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1001 _6666_/Q VGND VPWR _4270_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _4210_/X VGND VPWR _6610_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1023 _6676_/Q VGND VPWR _4282_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1034 _4216_/X VGND VPWR _6615_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ _6901_/Q _5976_/C _5971_/D _6829_/Q VGND VPWR _6067_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3279_ hold62/X hold81/A _6488_/Q VGND VPWR hold63/A VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_39_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1045 _6820_/Q VGND VPWR _5250_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1056 _5482_/X VGND VPWR _7026_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1067 _6834_/Q VGND VPWR _5266_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5018_ _5018_/A _5112_/C _5018_/C _5018_/D VGND VPWR _5021_/C VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1078 _5275_/X VGND VPWR _6842_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 _6805_/Q VGND VPWR _5233_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_731 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_207 _5171_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6969_ _6969_/CLK _6969_/D fanout474/X VGND VPWR _6969_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_146 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold890 _6738_/Q VGND VPWR hold890/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_580 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1590 _7181_/A VGND VPWR hold1590/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_698 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4320_ hold740/X _6356_/A1 _4321_/S VGND VPWR _4320_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_153_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4251_ _4251_/A0 _6353_/A1 _4255_/S VGND VPWR _4251_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3202_ _6957_/Q VGND VPWR _3202_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_141_588 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4182_ _3640_/Y _4182_/A1 _4186_/S VGND VPWR _6586_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_94_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6823_ _6951_/CLK _6823_/D fanout474/X VGND VPWR _6823_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6754_ _7011_/CLK _6754_/D fanout456/X VGND VPWR _6754_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3966_ _3966_/A0 _5491_/A1 _3980_/S VGND VPWR _3966_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_148_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5705_ _6820_/Q _5818_/A2 _5814_/B1 _6908_/Q _5704_/X VGND VPWR _5706_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6685_ _6707_/CLK _6685_/D fanout448/X VGND VPWR _6685_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3897_ _4702_/A _4566_/A VGND VPWR _4374_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_5636_ _6970_/Q _5634_/X _5635_/X _6826_/Q VGND VPWR _5636_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_191_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_327 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5567_ _6506_/Q _6508_/Q VGND VPWR _5567_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold120 _6412_/Q VGND VPWR _3292_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _7014_/Q VGND VPWR hold131/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _4515_/Y _4518_/B _4518_/C _4518_/D VGND VPWR _4522_/A VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_117_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold142 _5290_/X VGND VPWR _6856_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold153 _5450_/X VGND VPWR _6998_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ hold602/X _5543_/A1 hold77/X VGND VPWR _5498_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold164 _7008_/Q VGND VPWR hold164/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _5318_/X VGND VPWR _6881_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _6684_/Q VGND VPWR hold186/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4551_/A _4813_/A _4579_/B VGND VPWR _4948_/B VGND VPWR sky130_fd_sc_hd__nand3_4
Xhold197 _5243_/X VGND VPWR _6814_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7168_ _3945_/A1 _7168_/D _6398_/X VGND VPWR _7168_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_58_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6119_ _7052_/Q _5971_/A _5979_/X _6991_/Q _6105_/X VGND VPWR _6125_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7099_ _7113_/CLK _7099_/D fanout464/X VGND VPWR _7099_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_85_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_46 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_706 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3820_ _7071_/Q _5532_/A _4139_/A _6550_/Q VGND VPWR _3820_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_32_288 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3751_ _3751_/A _3751_/B _3751_/C _3751_/D VGND VPWR _3761_/C VGND VPWR sky130_fd_sc_hd__nor4_1
X_6470_ _6735_/CLK _6470_/D _3946_/B VGND VPWR _6470_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3682_ _6567_/Q _4157_/A _4250_/A _6652_/Q VGND VPWR _3682_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_145_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5421_ hold880/X _5484_/A1 _5426_/S VGND VPWR _5421_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_161_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput203 _3922_/X VGND VPWR mgmt_gpio_oeb[35] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput214 _3926_/X VGND VPWR mgmt_gpio_out[10] VGND VPWR sky130_fd_sc_hd__buf_12
X_5352_ hold449/X _5538_/A1 _5354_/S VGND VPWR _5352_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput225 _7187_/X VGND VPWR mgmt_gpio_out[22] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput236 _3923_/X VGND VPWR mgmt_gpio_out[32] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput247 _3928_/X VGND VPWR mgmt_gpio_out[8] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput258 _6746_/Q VGND VPWR pll90_sel[1] VGND VPWR sky130_fd_sc_hd__buf_12
X_4303_ hold838/X _5546_/A1 _4303_/S VGND VPWR _4303_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput269 _6743_/Q VGND VPWR pll_sel[1] VGND VPWR sky130_fd_sc_hd__buf_12
X_5283_ _5283_/A hold17/X VGND VPWR _5291_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_99_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7022_ _7051_/CLK _7022_/D fanout476/X VGND VPWR _7022_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4234_ hold413/X _5534_/A1 _4237_/S VGND VPWR _4234_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4165_ _3762_/Y _4165_/A1 _4171_/S VGND VPWR _6571_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_472 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4096_ hold168/X hold42/X _5202_/B VGND VPWR _4096_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6806_ _7051_/CLK _6806_/D fanout476/X VGND VPWR _6806_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4998_ _5068_/C _5069_/C _4998_/C VGND VPWR _5001_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_11_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3949_ _6403_/Q _3949_/B VGND VPWR _3950_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_6737_ _6739_/CLK _6737_/D _3946_/B VGND VPWR _6737_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6668_ _6668_/CLK _6668_/D fanout452/X VGND VPWR _6668_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_176_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5619_ _5664_/A _5666_/B _5666_/C VGND VPWR _5619_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_191_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6599_ _6654_/CLK _6599_/D fanout454/X VGND VPWR _6599_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_117_360 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_503 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout430 hold16/X VGND VPWR _4322_/B VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout441 _6396_/B VGND VPWR _6401_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xfanout452 fanout455/X VGND VPWR fanout452/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout463 fanout465/X VGND VPWR fanout463/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_58_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout474 fanout475/X VGND VPWR fanout474/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xfanout485 fanout486/X VGND VPWR fanout485/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_171_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_623 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_764 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_715 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5970_ _5600_/A _5969_/A _5981_/C _5943_/X _5965_/X VGND VPWR _5970_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_80_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4921_/A _5043_/A VGND VPWR _4921_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_33_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_350 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4852_ _4947_/B _4456_/Y _4902_/B _4628_/Y VGND VPWR _4852_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_3803_ input43/X _4058_/S _4102_/A input61/X VGND VPWR _3803_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_20_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4783_ _4846_/B _4644_/Y _4663_/Y _4782_/Y VGND VPWR _5108_/B VGND VPWR sky130_fd_sc_hd__o22a_1
X_6522_ _6990_/CLK _6522_/D fanout478/X VGND VPWR _6522_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3734_ _6656_/Q _4256_/A _4298_/A _6691_/Q VGND VPWR _3734_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_146_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6453_ _6655_/CLK _6453_/D _6383_/A VGND VPWR _6453_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_134_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3665_ _6436_/Q _3372_/Y _4280_/A _6677_/Q _3664_/X VGND VPWR _3670_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5404_ hold221/X _5494_/A1 _5408_/S VGND VPWR _5404_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6384_ _6401_/A _6400_/B VGND VPWR _6384_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3596_ _6861_/Q _5292_/A _3593_/X _3595_/X VGND VPWR _3596_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_5335_ hold940/X _5548_/A1 _5336_/S VGND VPWR _5335_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5266_ _5266_/A0 hold666/X _5273_/S VGND VPWR _5266_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7005_ _7017_/CLK _7005_/D fanout466/X VGND VPWR _7005_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4217_ hold662/X _5544_/A1 _4219_/S VGND VPWR _4217_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5197_ _5197_/A0 _5545_/A1 _5201_/S VGND VPWR _5197_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4148_ hold453/X _5544_/A1 _4150_/S VGND VPWR _4148_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4079_ hold742/X hold42/X _4083_/S VGND VPWR _4079_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_70_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_764 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold708 _6919_/Q VGND VPWR hold708/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 _5362_/X VGND VPWR _6920_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3450_ _7118_/Q _6760_/Q _6762_/Q VGND VPWR _3450_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_3381_ _3511_/A hold66/A VGND VPWR _3381_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
X_5120_ _4906_/Y _5120_/B _5120_/C VGND VPWR _5120_/X VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_34_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5051_ _5051_/A _5051_/B VGND VPWR _5089_/C VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold1408 _7005_/Q VGND VPWR _5458_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1419 _6586_/Q VGND VPWR hold1419/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4002_ hold886/X _5484_/A1 _4007_/S VGND VPWR _4002_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5953_ _5969_/A _5969_/C _5981_/C VGND VPWR _5953_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_40_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4904_ _4359_/Y _4900_/Y _4850_/Y VGND VPWR _5131_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_21_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5884_ _6547_/Q _5655_/X _5879_/X _5881_/X _5883_/X VGND VPWR _5884_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4835_ _4551_/B _4554_/B _4574_/A VGND VPWR _4835_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_21_578 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4766_ _4627_/A _4626_/Y _4643_/Y _4948_/C _4672_/B VGND VPWR _4767_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_6505_ _6537_/CLK _6505_/D fanout464/X VGND VPWR _7178_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3717_ hold28/X _3717_/B VGND VPWR _5145_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_107_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4697_ _4911_/B _4703_/B VGND VPWR _4697_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_20_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6436_ _6747_/CLK _6436_/D fanout447/X VGND VPWR _6436_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3648_ _3957_/A _4102_/A _3585_/Y input97/X _3647_/X VGND VPWR _3651_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6367_ _6383_/A _6367_/B VGND VPWR _6367_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_88_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3579_ _6870_/Q _5301_/A _4014_/A _6459_/Q _3578_/X VGND VPWR _3580_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5318_ _5318_/A0 hold22/X _5318_/S VGND VPWR _5318_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6298_ _6559_/Q _5971_/B _5949_/X _6679_/Q _6297_/X VGND VPWR _6300_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_556 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold13 hold9/X VGND VPWR hold13/X VGND VPWR sky130_fd_sc_hd__buf_6
Xhold24 hold24/A VGND VPWR hold24/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ hold287/X _5534_/A1 _5255_/S VGND VPWR _5249_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold35 hold35/A VGND VPWR hold35/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold46 hold46/A VGND VPWR hold46/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A VGND VPWR hold57/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A VGND VPWR hold68/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VPWR hold79/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XPHY_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_88 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_372 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4716_/A _4975_/A VGND VPWR _4620_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_187_185 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4551_ _4551_/A _4551_/B VGND VPWR _5088_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_144_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3502_ hold79/A _3999_/A _4256_/A _6659_/Q VGND VPWR _3502_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold505 _6553_/Q VGND VPWR hold505/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _4482_/A _4482_/B VGND VPWR _4972_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_171_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold516 _5316_/X VGND VPWR _6879_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 _6425_/Q VGND VPWR hold527/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 _5231_/X VGND VPWR _6803_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ _6561_/Q _5953_/X _5960_/X _6671_/Q _6220_/X VGND VPWR _6221_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_116_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold549 _6891_/Q VGND VPWR hold549/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _7032_/Q hold49/A _5463_/A _7016_/Q VGND VPWR _3433_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_131_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6152_ _6140_/Y _6151_/X _6792_/Q _6226_/B VGND VPWR _6152_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3364_ _3714_/A hold74/X VGND VPWR _5436_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_106_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5103_ _5103_/A _5103_/B _5103_/C VGND VPWR _5103_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_6083_ _6862_/Q _5943_/X _5981_/X _6918_/Q _6079_/X VGND VPWR _6083_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1205 _7002_/Q VGND VPWR _5455_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3295_ _3295_/A _3323_/B VGND VPWR _3295_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold1216 _5428_/X VGND VPWR _6978_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1227 _6898_/Q VGND VPWR _5338_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5034_ _5034_/A _5034_/B _5085_/B _5034_/D VGND VPWR _5035_/D VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1238 _4299_/X VGND VPWR _6690_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _7063_/Q VGND VPWR _5524_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_464 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6985_ _7033_/CLK _6985_/D fanout464/X VGND VPWR _6985_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_13_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5936_ _5968_/A _5981_/B _5969_/C VGND VPWR _5971_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_179_642 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5867_ _7153_/Q _5625_/X _5661_/X _6621_/Q VGND VPWR _5867_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_179_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4818_ _4902_/A _4456_/Y _4562_/Y _4948_/C VGND VPWR _4818_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_166_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5798_ _3227_/Y _5651_/Y _5787_/Y _5797_/Y _5552_/B VGND VPWR _5798_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4749_ _4413_/Y _4581_/B _4611_/Y _4616_/Y VGND VPWR _5099_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_147_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6419_ _7049_/CLK _6419_/D fanout457/X VGND VPWR _6419_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_103_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput103 wb_adr_i[13] VGND VPWR _4336_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput114 wb_adr_i[23] VGND VPWR _4334_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput125 wb_adr_i[4] VGND VPWR _4642_/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xinput136 wb_dat_i[13] VGND VPWR _6338_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput147 wb_dat_i[23] VGND VPWR _6345_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput158 wb_dat_i[4] VGND VPWR _6336_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_57_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput169 wb_stb_i VGND VPWR _3899_/D VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_29_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clkbuf_3_1_0_csclk/X VGND VPWR _6668_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_188_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_542 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_581 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_754 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6770_ _7080_/CLK _6770_/D fanout479/X VGND VPWR _7189_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3982_ _3982_/A0 _6353_/A1 _3989_/S VGND VPWR _3982_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_15_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_450 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5721_ _6949_/Q _5637_/X _5645_/X _7029_/Q VGND VPWR _5721_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_148_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5652_ _5899_/B _5652_/B VGND VPWR _5652_/Y VGND VPWR sky130_fd_sc_hd__nand2b_4
X_4603_ _4607_/A _4993_/B VGND VPWR _4682_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_129_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5583_ _5582_/Y _5664_/A _5583_/S VGND VPWR _5584_/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_175_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4534_ _4782_/A _4881_/B _5088_/A VGND VPWR _4535_/D VGND VPWR sky130_fd_sc_hd__a21boi_1
Xhold302 _5384_/X VGND VPWR _6939_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold313 _7062_/Q VGND VPWR hold313/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 _5518_/X VGND VPWR _7058_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _7049_/Q VGND VPWR hold335/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _4302_/X VGND VPWR _6693_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _4489_/A _4465_/B VGND VPWR _4493_/B VGND VPWR sky130_fd_sc_hd__and2_1
Xhold357 _6980_/Q VGND VPWR hold357/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold368 _5169_/X VGND VPWR _6753_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_439 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold379 _6991_/Q VGND VPWR hold379/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _6204_/A0 _6203_/X _6279_/S VGND VPWR _7127_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3416_ _3714_/B _3571_/B VGND VPWR _5182_/S VGND VPWR sky130_fd_sc_hd__nor2_8
X_7184_ _7184_/A VGND VPWR _7184_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4396_ _4396_/A _4396_/B VGND VPWR _4415_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_6135_ _6944_/Q _5961_/X _6131_/X _6134_/X VGND VPWR _6140_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3347_ _3347_/A _3356_/B VGND VPWR _3714_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_140_770 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_301 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1002 _4270_/X VGND VPWR _6666_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1013 _6519_/Q VGND VPWR _4104_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1024 _4282_/X VGND VPWR _6676_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6066_ _6066_/A _6066_/B _6066_/C VGND VPWR _6075_/C VGND VPWR sky130_fd_sc_hd__nor3_2
Xhold1035 _6551_/Q VGND VPWR _4141_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ hold83/X VGND VPWR _3453_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
Xhold1046 _5250_/X VGND VPWR _6820_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _6973_/Q VGND VPWR _5422_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _5106_/B _5064_/B _5062_/D VGND VPWR _5018_/D VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1068 _5266_/X VGND VPWR _6834_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1079 _6813_/Q VGND VPWR _5242_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_404 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6968_ _7069_/CLK _6968_/D fanout482/X VGND VPWR _6968_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5919_ _7038_/Q _5614_/X _5917_/X _5918_/X VGND VPWR _5919_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_6899_ _7080_/CLK _6899_/D fanout479/X VGND VPWR _6899_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_166_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_712 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold880 _6972_/Q VGND VPWR hold880/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold891 _5150_/X VGND VPWR _6738_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_269 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1580 _7100_/Q VGND VPWR _5596_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_592 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1591 _6528_/Q VGND VPWR hold812/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_158 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4250_ _4250_/A _5490_/B VGND VPWR _4255_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_3201_ _6965_/Q VGND VPWR _3201_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4181_ _3700_/Y _4181_/A1 _4186_/S VGND VPWR _6585_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_687 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6822_ _6884_/CLK _6822_/D fanout475/X VGND VPWR _6822_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_51_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_297 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6753_ _7011_/CLK _6753_/D fanout459/X VGND VPWR _6753_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3965_ _3251_/A hold664/X _3975_/S VGND VPWR _3965_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5704_ _6996_/Q _5643_/X _5652_/B _6916_/Q _5651_/Y VGND VPWR _5704_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6684_ _6714_/CLK _6684_/D fanout470/X VGND VPWR _6684_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3896_ _5552_/B _3887_/Y _5959_/A _5966_/A _3895_/X VGND VPWR _6509_/D VGND VPWR
+ sky130_fd_sc_hd__a41o_1
X_5635_ _5638_/A _5657_/B _5666_/C VGND VPWR _5635_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_163_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5566_ _3176_/Y _5564_/B _5565_/X VGND VPWR _7091_/D VGND VPWR sky130_fd_sc_hd__a21boi_1
Xhold110 _7006_/Q VGND VPWR hold110/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold121 _3292_/X VGND VPWR hold121/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _5468_/X VGND VPWR _7014_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _4953_/A _5042_/B VGND VPWR _4518_/C VGND VPWR sky130_fd_sc_hd__nand2_1
X_5497_ _5497_/A0 hold667/X hold77/A VGND VPWR _5497_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold143 _6985_/Q VGND VPWR hold143/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _7144_/Q VGND VPWR hold154/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _5461_/X VGND VPWR _7008_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold176 _7070_/Q VGND VPWR hold176/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4408_/B _4448_/B VGND VPWR _4579_/B VGND VPWR sky130_fd_sc_hd__and2b_4
Xhold187 _4291_/X VGND VPWR _6684_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _7037_/Q VGND VPWR hold198/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7167_ _3945_/A1 _7167_/D _6397_/X VGND VPWR _7167_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4379_ _4360_/B _4379_/B VGND VPWR _4384_/A VGND VPWR sky130_fd_sc_hd__nand2b_1
X_6118_ _6823_/Q _5953_/X _5960_/X _7076_/Q _6117_/X VGND VPWR _6118_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7098_ _7113_/CLK _7098_/D fanout462/X VGND VPWR _7098_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_18_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6049_ _6049_/A _6049_/B _6049_/C _6049_/D VGND VPWR _6049_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_37_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_614 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6714_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_134_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_698 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VPWR _6527_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_32_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3750_ input12/X _3358_/Y _4208_/A _6610_/Q _3749_/X VGND VPWR _3751_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3681_ _6836_/Q _5265_/A _5319_/A _6884_/Q _3680_/X VGND VPWR _3688_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_328 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5420_ hold634/X _5543_/A1 _5426_/S VGND VPWR _5420_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput204 _3921_/X VGND VPWR mgmt_gpio_oeb[36] VGND VPWR sky130_fd_sc_hd__buf_12
X_5351_ hold485/X _5528_/A1 _5354_/S VGND VPWR _5351_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput215 _7179_/X VGND VPWR mgmt_gpio_out[11] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput226 _7188_/X VGND VPWR mgmt_gpio_out[23] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput237 _3924_/X VGND VPWR mgmt_gpio_out[33] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput248 _3946_/Y VGND VPWR pad_flash_clk_oeb VGND VPWR sky130_fd_sc_hd__buf_12
X_4302_ hold345/X _5518_/A1 _4303_/S VGND VPWR _4302_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput259 _6747_/Q VGND VPWR pll90_sel[2] VGND VPWR sky130_fd_sc_hd__buf_12
X_5282_ hold624/X _5513_/A1 _5282_/S VGND VPWR _5282_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7021_ _7082_/CLK _7021_/D fanout483/X VGND VPWR _7021_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4233_ _4233_/A0 hold667/X _4237_/S VGND VPWR _4233_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4164_ _3828_/Y _4164_/A1 _4171_/S VGND VPWR _6570_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_665 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4095_ hold393/X _4094_/X _4101_/S VGND VPWR _4095_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6805_ _7085_/CLK _6805_/D fanout477/X VGND VPWR _6805_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_168_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4997_ _5073_/A _5103_/A _4997_/C _4997_/D VGND VPWR _4998_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_23_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6736_ _6739_/CLK _6736_/D _3946_/B VGND VPWR _6736_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3948_ _3948_/A VGND VPWR _3948_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_164_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6667_ _6668_/CLK _6667_/D fanout452/X VGND VPWR _6667_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3879_ _6642_/Q _3962_/B _3879_/B1 VGND VPWR _6642_/D VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_176_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5618_ _7093_/Q _7092_/Q VGND VPWR _5666_/C VGND VPWR sky130_fd_sc_hd__and2b_2
X_6598_ _7137_/CLK _6598_/D VGND VPWR _6598_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_5549_ _5549_/A0 hold22/X _5549_/S VGND VPWR hold23/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_372 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_407 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout420 hold13/X VGND VPWR _5534_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
Xfanout431 _5505_/B VGND VPWR _5541_/B VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout442 _3268_/Y VGND VPWR _6396_/B VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xfanout453 fanout454/X VGND VPWR _6401_/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xfanout464 fanout465/X VGND VPWR fanout464/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout475 fanout486/X VGND VPWR fanout475/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout486 input75/X VGND VPWR fanout486/X VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_101_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A VGND VPWR _7150_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_69_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4920_ _5023_/B _4920_/B _4964_/C VGND VPWR _5069_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_178_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4851_ _4413_/Y _4496_/Y _4616_/Y _4689_/A VGND VPWR _4877_/A VGND VPWR sky130_fd_sc_hd__o22a_1
X_3802_ input4/X _3381_/Y _4044_/A _6480_/Q _3801_/X VGND VPWR _3807_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4782_ _4782_/A _4975_/A VGND VPWR _4782_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_6521_ _6755_/CLK _6521_/D _6360_/A VGND VPWR _6521_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3733_ _6979_/Q _5427_/A _3414_/Y _3732_/X VGND VPWR _3733_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_118_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6452_ _6677_/CLK _6452_/D fanout452/X VGND VPWR _6452_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3664_ _6988_/Q _5436_/A _4139_/A _6552_/Q VGND VPWR _3664_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_134_618 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5403_ hold387/X _5526_/A1 _5408_/S VGND VPWR _5403_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6383_ _6383_/A _6401_/B VGND VPWR _6383_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3595_ input38/X _3331_/Y _4298_/A _6693_/Q _3594_/X VGND VPWR _3595_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5334_ hold417/X _5538_/A1 _5336_/S VGND VPWR _5334_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5265_ _5265_/A hold17/X VGND VPWR _5273_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_87_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7004_ _7012_/CLK _7004_/D fanout466/X VGND VPWR _7004_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4216_ _4216_/A0 _5492_/A1 _4219_/S VGND VPWR _4216_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5196_ hold858/X _5484_/A1 _5201_/S VGND VPWR _5196_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4147_ hold281/X _5534_/A1 _4150_/S VGND VPWR _4147_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4078_ hold349/X _4077_/X _4084_/S VGND VPWR _4078_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_381 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6719_ _7038_/CLK _6719_/D fanout455/X VGND VPWR _6719_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_364 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_568 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold709 _5361_/X VGND VPWR _6919_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap439 _4434_/B VGND VPWR _4591_/A VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_170_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3380_ hold65/X _3415_/B VGND VPWR hold66/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_170_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5050_ _4456_/Y _4946_/X _5049_/X _4820_/X VGND VPWR _5058_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_69_259 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1409 _6750_/Q VGND VPWR _5165_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4001_ hold263/X _5465_/A1 _4007_/S VGND VPWR _4001_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5952_ _5969_/A _5979_/A _5981_/A VGND VPWR _5952_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_46_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4903_ _4493_/B _5024_/B _4841_/X VGND VPWR _4905_/B VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5883_ _6580_/Q _5928_/A2 _5913_/B1 _6552_/Q _5882_/X VGND VPWR _5883_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4834_ _4413_/Y _4810_/B _4823_/X _4833_/X VGND VPWR _4834_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_21_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4765_ _4921_/A _4992_/B _4588_/Y VGND VPWR _4767_/B VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_193_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6504_ _6755_/CLK _6504_/D _6360_/A VGND VPWR _6504_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3716_ _6605_/Q _4202_/A _3714_/Y _6749_/Q _3715_/X VGND VPWR _3720_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4696_ _4694_/Y _4695_/Y _4482_/B VGND VPWR _4706_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_161_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6435_ _6746_/CLK _6435_/D fanout447/X VGND VPWR _6435_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3647_ _7020_/Q hold29/A _4196_/A _6601_/Q VGND VPWR _3647_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_162_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_49 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6366_ _6383_/A _6401_/B VGND VPWR _6366_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3578_ _6806_/Q _5229_/A _4102_/A _7199_/A VGND VPWR _3578_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5317_ hold918/X _5548_/A1 _5318_/S VGND VPWR _5317_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6297_ _7038_/Q _5601_/X _5959_/X _6719_/Q VGND VPWR _6297_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_88_568 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold14 hold14/A VGND VPWR hold14/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _5248_/A0 _5473_/A1 _5255_/S VGND VPWR _5248_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold25 hold25/A VGND VPWR hold25/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A VGND VPWR hold36/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_29_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold47 hold47/A VGND VPWR hold47/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_102_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold58 hold58/A VGND VPWR hold58/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A VGND VPWR hold69/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5179_ hold696/X _5469_/A1 _5181_/S VGND VPWR _5179_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_368 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_710 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4550_ _4947_/B _4553_/B VGND VPWR _4551_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_144_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3501_ _3555_/A _3546_/A VGND VPWR _4256_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold506 _4143_/X VGND VPWR _6553_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4481_ _4615_/B _4653_/C VGND VPWR _4482_/B VGND VPWR sky130_fd_sc_hd__nand2_4
Xhold517 _7068_/Q VGND VPWR hold517/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _3980_/X VGND VPWR _6425_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 _6484_/Q VGND VPWR hold539/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _6651_/Q _5973_/A _5948_/X _6696_/Q _6219_/X VGND VPWR _6220_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3432_ _6880_/Q _5310_/A _5238_/A _6816_/Q VGND VPWR _3432_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6151_ _6143_/X _6145_/X _6151_/C _6226_/B VGND VPWR _6151_/X VGND VPWR sky130_fd_sc_hd__and4bb_1
X_3363_ _3814_/A _3714_/A VGND VPWR _5505_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5102_ _4626_/Y _4663_/Y _4933_/C _5101_/X VGND VPWR _5138_/B VGND VPWR sky130_fd_sc_hd__o211a_1
X_6082_ _7083_/Q _5976_/B _5971_/C _7043_/Q VGND VPWR _6099_/B VGND VPWR sky130_fd_sc_hd__a22o_1
X_3294_ hold32/X _3975_/S hold121/X _3293_/Y VGND VPWR _3294_/X VGND VPWR sky130_fd_sc_hd__o31a_2
Xhold1206 _5455_/X VGND VPWR _7002_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1217 _6946_/Q VGND VPWR _5392_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1228 _5338_/X VGND VPWR _6898_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _5033_/A _5080_/B _5033_/C _5120_/B VGND VPWR _5034_/D VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1239 _7055_/Q VGND VPWR _5515_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6984_ _7001_/CLK _6984_/D fanout461/X VGND VPWR _6984_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_80_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5935_ _7101_/Q _7102_/Q VGND VPWR _5969_/C VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_40_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5866_ _3185_/Y _5899_/B _5651_/B VGND VPWR _5866_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_166_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4817_ _4817_/A _4972_/A VGND VPWR _5018_/A VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_178_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5797_ _5797_/A _5797_/B _5797_/C _5797_/D VGND VPWR _5797_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_31_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4748_ _4921_/A _4926_/B VGND VPWR _5074_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_135_702 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4679_ _4925_/B _4679_/B _4679_/C _4679_/D VGND VPWR _4682_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_107_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6418_ _6749_/CLK _6418_/D fanout449/X VGND VPWR _6418_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6349_ _6643_/Q _6319_/B _6348_/X VGND VPWR _6349_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_0_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_759 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput104 wb_adr_i[14] VGND VPWR _4336_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput115 wb_adr_i[24] VGND VPWR _3904_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput126 wb_adr_i[5] VGND VPWR _4739_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_76_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput137 wb_dat_i[14] VGND VPWR _6341_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_dat_i[24] VGND VPWR _6324_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VPWR _6339_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_56_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_593 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3981_ _3981_/A _6352_/B VGND VPWR _3989_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_5720_ _6941_/Q _5632_/X _5638_/X _6957_/Q VGND VPWR _5720_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5651_ _5899_/B _5651_/B VGND VPWR _5651_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
X_4602_ _4993_/B VGND VPWR _4602_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_175_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5582_ _5664_/A _5602_/A VGND VPWR _5582_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_191_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4533_ _4490_/Y _5083_/A _4912_/A _4533_/D VGND VPWR _4535_/C VGND VPWR sky130_fd_sc_hd__and4b_1
Xhold303 _6713_/Q VGND VPWR hold303/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _5522_/X VGND VPWR _7062_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _6924_/Q VGND VPWR hold325/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4464_ _5051_/B VGND VPWR _4464_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xhold336 _5508_/X VGND VPWR _7049_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _6663_/Q VGND VPWR hold347/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _5430_/X VGND VPWR _6980_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 _6836_/Q VGND VPWR hold369/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6203_/A0 _6202_/X _6303_/S VGND VPWR _6203_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3415_ hold84/X _3415_/B VGND VPWR _3571_/B VGND VPWR sky130_fd_sc_hd__nand2_8
X_7183_ _7183_/A VGND VPWR _7183_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4395_ _4642_/A _4441_/B VGND VPWR _4396_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_6134_ _7016_/Q _5940_/X _5967_/X _6856_/Q _6130_/X VGND VPWR _6134_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3346_ _3347_/A _3355_/B hold72/X VGND VPWR _5190_/B VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_85_313 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1003 _6725_/Q VGND VPWR hold1003/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 _4104_/X VGND VPWR _6519_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6065_ _6981_/Q _5945_/X _5975_/C _6837_/Q _6064_/X VGND VPWR _6066_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3277_ hold82/X _4988_/B2 _3975_/S VGND VPWR hold83/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xhold1025 _6561_/Q VGND VPWR _4153_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1036 _4141_/X VGND VPWR _6551_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 _6884_/Q VGND VPWR _5322_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 _5422_/X VGND VPWR _6973_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _4644_/Y _4975_/Y _4991_/X _5011_/X VGND VPWR _5062_/D VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_39_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1069 _6933_/Q VGND VPWR _5377_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_9 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6967_ _6967_/CLK _6967_/D fanout474/X VGND VPWR _6967_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_41_416 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_596 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5918_ _6484_/Q _5643_/X _5664_/X _6669_/Q VGND VPWR _5918_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6898_ _7083_/CLK _6898_/D fanout476/X VGND VPWR _6898_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_22_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5849_ _7035_/Q _5614_/X _5643_/X _6481_/Q VGND VPWR _5849_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_158_47 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_598 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold870 _6467_/Q VGND VPWR hold870/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_546 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold881 _5421_/X VGND VPWR _6972_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _6448_/Q VGND VPWR hold892/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_760 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1570 _7158_/Q VGND VPWR _3868_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1581 _6760_/Q VGND VPWR hold696/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1592 _7101_/Q VGND VPWR _5598_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3200_ _6973_/Q VGND VPWR _3200_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4180_ _3762_/Y _4180_/A1 _4186_/S VGND VPWR _6584_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_121_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_699 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6821_ _7076_/CLK _6821_/D fanout481/X VGND VPWR _6821_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_50_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6752_ _7011_/CLK _6752_/D fanout456/X VGND VPWR _6752_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3964_ _3964_/A _6352_/B VGND VPWR _3980_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_5703_ _6444_/Q _5614_/X _5664_/X _6924_/Q _5702_/X VGND VPWR _5706_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6683_ _6683_/CLK _6683_/D _6390_/A VGND VPWR _6683_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3895_ _7088_/Q _3886_/B _7090_/Q _7091_/Q _6509_/Q VGND VPWR _3895_/X VGND VPWR
+ sky130_fd_sc_hd__o41a_1
XFILLER_176_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5634_ _5638_/A _5667_/B _5657_/B VGND VPWR _5634_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_176_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5565_ _3176_/Y _5564_/B _5564_/A VGND VPWR _5565_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_163_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold100 _4125_/X VGND VPWR _6538_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold111 _5459_/X VGND VPWR _7006_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4531_/B _4953_/A VGND VPWR _4518_/B VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold122 _3294_/X VGND VPWR _3323_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold133 _6757_/Q VGND VPWR hold133/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ hold76/X _5541_/B VGND VPWR hold77/A VGND VPWR sky130_fd_sc_hd__and2_4
Xhold144 _5435_/X VGND VPWR _6985_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold155 _3971_/X VGND VPWR hold94/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold166 _6838_/Q VGND VPWR hold166/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _4454_/A _4611_/B VGND VPWR _4902_/A VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold177 _5531_/X VGND VPWR _7070_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold188 _6822_/Q VGND VPWR hold188/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _5494_/X VGND VPWR _7037_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7166_ net399_2/A _7166_/D _6396_/X VGND VPWR hold20/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4378_ _4360_/B _4379_/B VGND VPWR _4900_/A VGND VPWR sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_1_csclk clkbuf_3_1_0_csclk/X VGND VPWR _6677_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6117_ _6911_/Q _5973_/A _5948_/X _6951_/Q _6116_/X VGND VPWR _6117_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3329_ hold47/X hold65/X VGND VPWR _3373_/B VGND VPWR sky130_fd_sc_hd__nand2_8
X_7097_ _7113_/CLK _7097_/D fanout462/X VGND VPWR _7097_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_73_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6048_ _6812_/Q _5971_/B _5949_/X _6932_/Q _6047_/X VGND VPWR _6049_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_160_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_619 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_460 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_555 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3680_ _6812_/Q _5238_/A hold76/A _7041_/Q VGND VPWR _3680_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5350_ _5350_/A0 _5545_/A1 _5354_/S VGND VPWR _5350_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput205 _3920_/X VGND VPWR mgmt_gpio_oeb[37] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput216 _7180_/X VGND VPWR mgmt_gpio_out[12] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput227 _7189_/X VGND VPWR mgmt_gpio_out[24] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput238 _7197_/X VGND VPWR mgmt_gpio_out[34] VGND VPWR sky130_fd_sc_hd__buf_12
X_4301_ hold457/X _5544_/A1 _4303_/S VGND VPWR _4301_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput249 _3943_/X VGND VPWR pad_flash_csb VGND VPWR sky130_fd_sc_hd__buf_12
X_5281_ hold922/X _5548_/A1 _5282_/S VGND VPWR _5281_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7020_ _7051_/CLK _7020_/D fanout476/X VGND VPWR _7020_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4232_ _4232_/A _4322_/B VGND VPWR _4237_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_4163_ _6639_/Q _6307_/B VGND VPWR _4171_/S VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_68_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4094_ hold766/X _5519_/A1 _5202_/B VGND VPWR _4094_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_63_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6804_ _7067_/CLK _6804_/D fanout477/X VGND VPWR _6804_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_169_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4996_ _5021_/A _4996_/B _4996_/C _4996_/D VGND VPWR _4997_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6735_ _6735_/CLK _6735_/D _3946_/B VGND VPWR _6735_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3947_ _6404_/Q _3947_/B VGND VPWR _3948_/A VGND VPWR sky130_fd_sc_hd__nand2b_1
X_6666_ _6668_/CLK _6666_/D fanout452/X VGND VPWR _6666_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3878_ hold15/A _6402_/Q _6396_/B VGND VPWR _3961_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_136_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5617_ _6442_/Q _5614_/X _5616_/X _6842_/Q VGND VPWR _5617_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6597_ _7137_/CLK _6597_/D VGND VPWR _6597_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_164_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5548_ hold926/X _5548_/A1 _5549_/S VGND VPWR _5548_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_155_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5479_ hold315/X _5521_/A1 hold30/X VGND VPWR _5479_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xfanout410 hold156/X VGND VPWR _5518_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_120_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout421 _6353_/A1 VGND VPWR _5491_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout432 hold16/X VGND VPWR _5505_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xfanout454 fanout455/X VGND VPWR fanout454/X VGND VPWR sky130_fd_sc_hd__buf_6
X_7149_ _3937_/A1 _7149_/D fanout487/X VGND VPWR _7149_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xfanout465 fanout466/X VGND VPWR fanout465/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout476 fanout485/X VGND VPWR fanout476/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout487 _6307_/B VGND VPWR fanout487/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_58_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_176 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4850_ _4456_/A _4843_/B _4689_/Y VGND VPWR _4850_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_33_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3801_ _6978_/Q _5427_/A _3714_/Y _6748_/Q VGND VPWR _3801_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4781_ _4846_/B _4689_/B _4780_/Y _4627_/A VGND VPWR _4781_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6520_ _6777_/CLK _6520_/D fanout484/X VGND VPWR _7197_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_186_560 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3732_ _6626_/Q _4232_/A _3692_/Y _6766_/Q _3731_/X VGND VPWR _3732_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6451_ _6677_/CLK _6451_/D fanout452/X VGND VPWR _6451_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3663_ _6964_/Q _5409_/A _3381_/Y input26/X _3662_/X VGND VPWR _3670_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5402_ hold249/X _5465_/A1 _5408_/S VGND VPWR _5402_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6382_ _6401_/A _6401_/B VGND VPWR _6382_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3594_ _6612_/Q _4208_/A _4196_/A _6602_/Q VGND VPWR _3594_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_114_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5333_ hold479/X _5528_/A1 _5336_/S VGND VPWR _5333_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5264_ hold679/X _5540_/A1 _5264_/S VGND VPWR _5264_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7003_ _7012_/CLK _7003_/D fanout458/X VGND VPWR _7003_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4215_ _4215_/A0 _6353_/A1 _4219_/S VGND VPWR _4215_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5195_ hold547/X _5543_/A1 _5201_/S VGND VPWR _5195_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4146_ _4146_/A0 hold667/X _4150_/S VGND VPWR _4146_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4077_ hold158/X hold60/X _4083_/S VGND VPWR _4077_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_706 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4979_ _4626_/Y _4644_/Y _4663_/Y _4782_/Y _4978_/X VGND VPWR _4981_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6718_ _7038_/CLK _6718_/D fanout455/X VGND VPWR _6718_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_177_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6649_ _6654_/CLK _6649_/D _6383_/A VGND VPWR _6649_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_180_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VPWR _6777_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_133_630 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_376 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_csclk _7001_/CLK VGND VPWR _7033_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_74_400 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_750 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4000_ _4000_/A0 _5524_/A1 _4007_/S VGND VPWR _4000_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_488 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5951_ _5969_/A _5966_/A _5979_/A VGND VPWR _5976_/B VGND VPWR sky130_fd_sc_hd__and3_4
X_4902_ _4902_/A _4902_/B VGND VPWR _5024_/B VGND VPWR sky130_fd_sc_hd__nand2_1
X_5882_ _6467_/Q _5619_/X _5663_/X _6611_/Q VGND VPWR _5882_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4833_ _4542_/B _4810_/B _5057_/A _4832_/X VGND VPWR _4833_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_178_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4764_ _4737_/A _4608_/X _4686_/B _4738_/A _4763_/X VGND VPWR _4764_/X VGND VPWR
+ sky130_fd_sc_hd__a311o_1
XFILLER_193_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6503_ _6537_/CLK _6503_/D fanout464/X VGND VPWR _7177_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3715_ _6955_/Q _5400_/A _4157_/A _6566_/Q VGND VPWR _3715_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4695_ _4716_/A _4969_/A VGND VPWR _4695_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_119_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6434_ _6746_/CLK _6434_/D fanout447/X VGND VPWR _6434_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_162_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3646_ _6682_/Q _4286_/A _4145_/A _6557_/Q _3645_/X VGND VPWR _3651_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_736 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6365_ _6383_/A _6401_/B VGND VPWR _6365_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3577_ hold74/X _3577_/B VGND VPWR _4014_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5316_ hold515/X _5538_/A1 _5318_/S VGND VPWR _5316_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6296_ _6459_/Q _5944_/X _5975_/A _6603_/Q _6295_/X VGND VPWR _6300_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5247_ _5247_/A _5541_/B VGND VPWR _5255_/S VGND VPWR sky130_fd_sc_hd__and2_4
Xhold15 hold15/A VGND VPWR hold15/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_666 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold26 hold26/A VGND VPWR hold26/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A VGND VPWR hold37/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_603 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold48 hold48/A VGND VPWR hold48/X VGND VPWR sky130_fd_sc_hd__buf_8
Xhold59 hold59/A VGND VPWR hold59/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ hold359/X _5526_/A1 _5181_/S VGND VPWR _5178_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4129_ hold808/X _6354_/A1 _4132_/S VGND VPWR _4129_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_414 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_385 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_506 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_580 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_744 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_388 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3500_ input7/X _3365_/Y _4280_/A _6679_/Q _3498_/X VGND VPWR _3504_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4480_ _4615_/B _4653_/C VGND VPWR _4636_/A VGND VPWR sky130_fd_sc_hd__and2_2
Xhold507 _6453_/Q VGND VPWR hold507/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 _5529_/X VGND VPWR _7068_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold529 _6608_/Q VGND VPWR hold529/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3431_ _3431_/A _3431_/B VGND VPWR _3447_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_171_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6150_ _6150_/A _6150_/B _6150_/C _6150_/D VGND VPWR _6151_/C VGND VPWR sky130_fd_sc_hd__nor4_1
X_3362_ _3714_/A _3573_/A VGND VPWR _5364_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5101_ _4846_/B _4644_/Y _4997_/D _5100_/Y VGND VPWR _5101_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_112_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6081_ _7059_/Q _5954_/X _5976_/D _6878_/Q VGND VPWR _6099_/A VGND VPWR sky130_fd_sc_hd__a22o_1
X_3293_ _6726_/Q _3975_/S VGND VPWR _3293_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold1207 _6426_/Q VGND VPWR _3982_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5032_ _4662_/Y _4695_/Y _4847_/Y _4905_/B _4508_/D VGND VPWR _5120_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_85_539 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1218 _5392_/X VGND VPWR _6946_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _7039_/Q VGND VPWR _5497_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6983_ _6997_/CLK _6983_/D fanout465/X VGND VPWR _6983_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_18_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5934_ _5966_/A _5968_/A _5981_/B VGND VPWR _5934_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_288 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5865_ _5864_/Y _5863_/X _6279_/S _5865_/B2 VGND VPWR _7115_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_4816_ _4947_/B _4947_/C _4553_/B VGND VPWR _4816_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5796_ _6880_/Q _5661_/X _5663_/X _6864_/Q _5795_/X VGND VPWR _5797_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4747_ _4747_/A _4747_/B _4747_/C VGND VPWR _4926_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_135_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_500 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4678_ _4741_/A wire380/X _4660_/X _4648_/X _4942_/B VGND VPWR _4679_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_162_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6417_ _3945_/A1 _6417_/D _6373_/X VGND VPWR _6417_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3629_ _7005_/Q _3370_/Y _5490_/A _7037_/Q VGND VPWR _3629_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_162_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6348_ _6644_/Q _6320_/A _6318_/B _6642_/Q VGND VPWR _6348_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput105 wb_adr_i[15] VGND VPWR _4336_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6279_ _6279_/A0 _6278_/X _6279_/S VGND VPWR _7130_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_452 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput116 wb_adr_i[25] VGND VPWR _3906_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_88_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput127 wb_adr_i[6] VGND VPWR _4631_/D VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_102_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput138 wb_dat_i[15] VGND VPWR _6344_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VPWR _6327_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_458 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3980_ hold527/X _5513_/A1 _3980_/S VGND VPWR _3980_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5650_ _5658_/B _5667_/C VGND VPWR _5651_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_30_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4601_ _4601_/A _4601_/B VGND VPWR _4993_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_5581_ _5583_/S _5580_/X _5574_/Y VGND VPWR _7095_/D VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_7_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4810_/A _4453_/B _4530_/X _4823_/A VGND VPWR _4533_/D VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_190_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold304 _4326_/X VGND VPWR _6713_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _7024_/Q VGND VPWR hold315/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _5367_/X VGND VPWR _6924_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4463_ _4911_/A _4856_/A VGND VPWR _5051_/B VGND VPWR sky130_fd_sc_hd__and2_2
Xhold337 _6988_/Q VGND VPWR hold337/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _4266_/X VGND VPWR _6663_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6189_/Y _6201_/X _6540_/Q _6226_/B VGND VPWR _6202_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3414_ hold85/A _3511_/A VGND VPWR _3414_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
Xhold359 _6759_/Q VGND VPWR hold359/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7182_ _7182_/A VGND VPWR _7182_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_98_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4394_ _4393_/A _4393_/B _4568_/B VGND VPWR _4551_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_6133_ _7085_/Q _5976_/B _5971_/C _7045_/Q VGND VPWR _6150_/B VGND VPWR sky130_fd_sc_hd__a22o_1
X_3345_ _3355_/B hold72/X VGND VPWR _3356_/B VGND VPWR sky130_fd_sc_hd__and2_2
Xhold1004 _3297_/Y VGND VPWR _3298_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6064_ _6925_/Q _5938_/X _5952_/X _6957_/Q VGND VPWR _6064_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_85_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1015 _6461_/Q VGND VPWR _4022_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3276_ hold81/X hold24/X _6488_/Q VGND VPWR hold82/A VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1026 _4153_/X VGND VPWR _6561_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 _6716_/Q VGND VPWR _4330_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _4653_/Y _4970_/Y _5010_/Y _4645_/Y _4807_/X VGND VPWR _5064_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_100_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1048 _5322_/X VGND VPWR _6884_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 _6901_/Q VGND VPWR _5341_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6966_ _7083_/CLK _6966_/D fanout476/X VGND VPWR _6966_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_41_428 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5917_ _6564_/Q _5631_/X _5646_/X _6654_/Q VGND VPWR _5917_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6897_ _7076_/CLK _6897_/D fanout481/X VGND VPWR _6897_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_675 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5848_ _6476_/Q _5630_/X _5634_/X _6451_/Q VGND VPWR _5848_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_158_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_59 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5779_ _6960_/Q _5638_/X _5648_/X _6856_/Q VGND VPWR _5779_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_166_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_706 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold860 _6876_/Q VGND VPWR hold860/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _4029_/X VGND VPWR _6467_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _6975_/Q VGND VPWR hold882/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_558 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold893 _4006_/X VGND VPWR _6448_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1560 hold70/A VGND VPWR _3855_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 _7170_/Q VGND VPWR _3235_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1582 _6533_/Q VGND VPWR hold824/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 _6498_/Q VGND VPWR hold1593/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_189_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_458 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_511 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_406 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_572 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6820_ _6884_/CLK _6820_/D fanout475/X VGND VPWR _6820_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6751_ _7011_/CLK _6751_/D fanout459/X VGND VPWR _6751_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3963_ hold15/X _3963_/A1 _3963_/S VGND VPWR hold16/A VGND VPWR sky130_fd_sc_hd__mux2_8
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VPWR clkbuf_1_1_1_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
X_5702_ _6964_/Q _5642_/X _5667_/X _6812_/Q VGND VPWR _5702_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6682_ _6683_/CLK _6682_/D _6390_/A VGND VPWR _6682_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3894_ _5552_/B _3887_/Y _3893_/Y _6763_/Q _3894_/B2 VGND VPWR _6508_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_148_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5633_ _6818_/Q _5631_/X _5632_/X _6938_/Q VGND VPWR _5633_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_12_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5564_ _5564_/A _5564_/B _5564_/C VGND VPWR _7090_/D VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_128_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_149 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold101 _6724_/Q VGND VPWR hold101/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _4542_/A _4947_/B VGND VPWR _4515_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold112 _7000_/Q VGND VPWR hold112/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _3295_/Y VGND VPWR _3355_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5495_ hold235/X hold60/X _5495_/S VGND VPWR _5495_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold134 _5176_/X VGND VPWR _6757_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _7053_/Q VGND VPWR hold145/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4495_/A _4993_/A VGND VPWR _4531_/B VGND VPWR sky130_fd_sc_hd__nor2_2
Xhold156 hold94/X VGND VPWR hold156/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _5270_/X VGND VPWR _6838_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold178 _7059_/Q VGND VPWR hold178/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _5252_/X VGND VPWR _6822_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7165_ net399_2/A _7165_/D _6395_/X VGND VPWR hold97/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4377_ _4471_/B _4568_/B VGND VPWR _4887_/A VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_86_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6116_ _6903_/Q _5976_/C _5971_/D _6831_/Q VGND VPWR _6116_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3328_ _3571_/A hold85/X VGND VPWR _5229_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_271 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7096_ _7113_/CLK _7096_/D fanout462/X VGND VPWR _7096_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_86_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6047_ _6444_/Q _5601_/X _5959_/X _6964_/Q VGND VPWR _6047_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3259_ _3260_/A1 _3259_/A1 _3260_/S VGND VPWR _7161_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_499 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6949_ _7085_/CLK _6949_/D fanout477/X VGND VPWR _6949_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_139_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_650 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold690 _7033_/Q VGND VPWR hold690/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_472 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_61 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1390 _5214_/X VGND VPWR hold19/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_567 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput206 _3173_/Y VGND VPWR mgmt_gpio_oeb[3] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput217 _3938_/X VGND VPWR mgmt_gpio_out[13] VGND VPWR sky130_fd_sc_hd__buf_12
X_4300_ hold277/X _5534_/A1 _4303_/S VGND VPWR _4300_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput228 _7190_/X VGND VPWR mgmt_gpio_out[25] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_154_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput239 _3925_/X VGND VPWR mgmt_gpio_out[35] VGND VPWR sky130_fd_sc_hd__buf_12
X_5280_ hold780/X _5538_/A1 _5282_/S VGND VPWR _5280_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4231_ _6624_/Q _3170_/Y _4228_/Y _5006_/A _3168_/A VGND VPWR _4231_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_99_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4162_ hold233/X hold60/X _4162_/S VGND VPWR _4162_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_431 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4093_ _4093_/A0 _4092_/X _4101_/S VGND VPWR _4093_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6803_ _7067_/CLK _6803_/D fanout477/X VGND VPWR _6803_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4995_ _4995_/A _4995_/B _4995_/C VGND VPWR _5004_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_168_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6734_ _3945_/A1 _6734_/D _6386_/X VGND VPWR _6734_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_3946_ _6403_/Q _3946_/B VGND VPWR _3946_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_177_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6665_ _6755_/CLK _6665_/D _6360_/A VGND VPWR _6665_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3877_ hold15/A _6402_/Q _6396_/B VGND VPWR _3962_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_5616_ _5638_/A _5667_/B _5657_/B VGND VPWR _5616_/X VGND VPWR sky130_fd_sc_hd__and3b_4
X_6596_ _7137_/CLK _6596_/D VGND VPWR _6596_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_5547_ _5547_/A0 hold42/X _5549_/S VGND VPWR hold43/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_155_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5478_ hold56/X hold42/X hold30/X VGND VPWR hold57/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_132_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4429_ _4685_/A _4992_/A VGND VPWR _5068_/A VGND VPWR sky130_fd_sc_hd__nand2_2
Xfanout400 hold54/X VGND VPWR hold42/A VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout411 _5526_/A1 VGND VPWR _6355_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout422 hold666/X VGND VPWR _6353_/A1 VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_160_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout433 _3178_/Y VGND VPWR _6303_/S VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout444 fanout486/X VGND VPWR _3946_/B VGND VPWR sky130_fd_sc_hd__buf_8
X_7148_ _3937_/A1 _7148_/D _6307_/B VGND VPWR _7148_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xfanout455 fanout486/X VGND VPWR fanout455/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout466 fanout486/X VGND VPWR fanout466/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout477 fanout485/X VGND VPWR fanout477/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout488 input164/X VGND VPWR _6307_/B VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_7079_ _7079_/CLK _7079_/D fanout478/X VGND VPWR _7079_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_58_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_670 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3800_ _6614_/Q _4214_/A _4133_/A _6545_/Q _3799_/X VGND VPWR _3807_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4780_ _4782_/A _4707_/C _4574_/B VGND VPWR _4780_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3731_ _6803_/Q _5229_/A _4172_/A _6579_/Q VGND VPWR _3731_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6709_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6450_ _6677_/CLK _6450_/D fanout452/X VGND VPWR _6450_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3662_ _6687_/Q _4292_/A hold67/A _6467_/Q VGND VPWR _3662_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_118_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5401_ _5401_/A0 _5524_/A1 _5408_/S VGND VPWR _5401_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6381_ _6401_/A _6401_/B VGND VPWR _6381_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3593_ _6901_/Q _5337_/A _5274_/A _6845_/Q _3592_/X VGND VPWR _3593_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5332_ _5332_/A0 _5545_/A1 _5336_/S VGND VPWR _5332_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_126_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5263_ hold671/X _5521_/A1 _5264_/S VGND VPWR _5263_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7002_ _7006_/CLK _7002_/D fanout458/X VGND VPWR _7002_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4214_ _4214_/A _4322_/B VGND VPWR _4219_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_5194_ _5194_/A0 _5473_/A1 _5201_/S VGND VPWR _5194_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4145_ _4145_/A _4322_/B VGND VPWR _4150_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_4076_ _4076_/A0 hold95/X _4084_/S VGND VPWR hold96/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4978_ _4639_/Y _4692_/Y _4969_/Y _4663_/Y VGND VPWR _4978_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6717_ _7038_/CLK _6717_/D fanout455/X VGND VPWR _6717_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_20_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3929_ _6504_/Q input77/X _3956_/B VGND VPWR _3929_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_50_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6648_ _6671_/CLK _6648_/D fanout468/X VGND VPWR _6648_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_125_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6579_ _6677_/CLK _6579_/D fanout452/X VGND VPWR _6579_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_180_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_684 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_762 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_303 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5950_ _6946_/Q _5948_/X _5949_/X _6930_/Q VGND VPWR _5950_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_92_275 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4901_ _4491_/Y _4900_/Y _4707_/Y _4498_/Y VGND VPWR _5080_/A VGND VPWR sky130_fd_sc_hd__o211a_1
X_5881_ _6601_/Q _5616_/X _5880_/X VGND VPWR _5881_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_61_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4832_ _4948_/A _4810_/B _5092_/A _4831_/X VGND VPWR _4832_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XANTENNA_190 _5513_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4763_ _4921_/A _4737_/A _4668_/C _4671_/A VGND VPWR _4763_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_159_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6502_ _6539_/CLK _6502_/D fanout461/X VGND VPWR _7176_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3714_ _3714_/A _3714_/B VGND VPWR _3714_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4694_ _4716_/A _4782_/A VGND VPWR _4694_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_6433_ _6749_/CLK _6433_/D fanout449/X VGND VPWR _6433_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3645_ input37/X _3331_/Y _4202_/A _6606_/Q VGND VPWR _3645_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_20_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6364_ _6383_/A _6401_/B VGND VPWR _6364_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3576_ _6982_/Q _5427_/A _5490_/A _7038_/Q _3574_/X VGND VPWR _3580_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5315_ hold465/X _5528_/A1 _5318_/S VGND VPWR _5315_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6295_ _6469_/Q _5937_/X _5975_/D _6629_/Q VGND VPWR _6295_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_114_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5246_ hold762/X _5540_/A1 _5246_/S VGND VPWR _5246_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VPWR hold16/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A VGND VPWR hold27/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_130_678 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold38 hold38/A VGND VPWR hold38/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A VGND VPWR hold49/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ hold209/X _5494_/A1 _5181_/S VGND VPWR _5177_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4128_ _4128_/A0 _5491_/A1 _4132_/S VGND VPWR _4128_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_659 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_618 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4059_ hold997/X _4058_/X _4067_/S VGND VPWR _4059_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_426 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_736 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_61 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_80_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6755_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold508 _4012_/X VGND VPWR _6453_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold519 _6682_/Q VGND VPWR hold519/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3430_ _5182_/S _3417_/X _3426_/X _3428_/X _3429_/X VGND VPWR _3431_/B VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_109_491 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3361_ _3562_/A hold48/X VGND VPWR _5265_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_612 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5100_ _4992_/A _4737_/A _4735_/X _4588_/Y VGND VPWR _5100_/Y VGND VPWR sky130_fd_sc_hd__a31oi_1
XFILLER_32_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6080_ _7006_/Q _5958_/X _5978_/X _6998_/Q VGND VPWR _6080_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3292_ _3292_/A _6488_/Q VGND VPWR _3292_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_112_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5031_ _4542_/A _4902_/A _4695_/Y _4627_/B _4872_/D VGND VPWR _5033_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold1208 _3982_/X VGND VPWR _6426_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _7047_/Q VGND VPWR _5506_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6982_ _7065_/CLK _6982_/D fanout465/X VGND VPWR _6982_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5933_ _5966_/A _5979_/A _5981_/B VGND VPWR _5971_/A VGND VPWR sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7086_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_33_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5864_ _5552_/B _7114_/Q _6103_/B1 VGND VPWR _5864_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_4815_ _4947_/C _4553_/B _5041_/A VGND VPWR _4815_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_193_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5795_ _7024_/Q _5619_/X _5666_/X _6896_/Q VGND VPWR _5795_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_193_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_48_csclk _7001_/CLK VGND VPWR _6981_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4746_ _4948_/A _4581_/B _4611_/Y _4645_/Y VGND VPWR _4942_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_193_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_406 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4677_ _4500_/A _4902_/B _4535_/A _5021_/A VGND VPWR _4679_/C VGND VPWR sky130_fd_sc_hd__o211a_1
X_6416_ _3927_/A1 _6416_/D _6372_/X VGND VPWR _6416_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3628_ _3628_/A _3628_/B _3628_/C _3628_/D VGND VPWR _3639_/B VGND VPWR sky130_fd_sc_hd__nor4_1
X_6347_ _6347_/A1 _4228_/Y _4229_/X _3910_/A VGND VPWR _7149_/D VGND VPWR sky130_fd_sc_hd__o211a_2
X_3559_ _3714_/B _3814_/B VGND VPWR _4133_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_163_38 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6278_ _6278_/A0 _6277_/X _6303_/S VGND VPWR _6278_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput106 wb_adr_i[16] VGND VPWR _4335_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VPWR _3900_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_130_464 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput128 wb_adr_i[7] VGND VPWR _4633_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_88_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput139 wb_dat_i[16] VGND VPWR _6323_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5229_ _5229_/A _5541_/B VGND VPWR _5237_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_102_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_90 _6558_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_125_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VPWR clkbuf_3_7_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_79_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_326 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4600_ _4739_/A _4600_/B _4747_/B _4739_/B VGND VPWR _4601_/B VGND VPWR sky130_fd_sc_hd__nand4b_1
X_5580_ _7094_/Q _5576_/B _7095_/Q VGND VPWR _5580_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_30_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4531_ _4810_/A _4531_/B VGND VPWR _4823_/A VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_184_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold305 _6915_/Q VGND VPWR hold305/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold316 _5479_/X VGND VPWR _7024_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _4896_/A _4462_/B VGND VPWR _4856_/A VGND VPWR sky130_fd_sc_hd__and2_1
Xhold327 _6857_/Q VGND VPWR hold327/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _5439_/X VGND VPWR _6988_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold349 hold349/A VGND VPWR hold349/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6192_/X _6201_/B _6226_/B VGND VPWR _6201_/X VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_144_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3413_ _3412_/X _3413_/A1 _3829_/B VGND VPWR _6734_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_7181_ _7181_/A VGND VPWR _7181_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4393_ _4393_/A _4393_/B VGND VPWR _4552_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_98_632 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6132_ _7061_/Q _5954_/X _5976_/D _6880_/Q VGND VPWR _6150_/A VGND VPWR sky130_fd_sc_hd__a22o_1
X_3344_ _3374_/A hold48/X VGND VPWR _5337_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6063_ _6973_/Q _5947_/X _5965_/X _6797_/Q _6062_/X VGND VPWR _6066_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3275_ hold46/X hold26/X VGND VPWR hold47/A VGND VPWR sky130_fd_sc_hd__and2b_4
Xhold1005 _3298_/Y VGND VPWR hold72/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 _4022_/X VGND VPWR _6461_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1027 _6601_/Q VGND VPWR _4199_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 _4330_/X VGND VPWR _6716_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _4628_/Y _5010_/Y _4982_/X _4796_/A VGND VPWR _5018_/C VGND VPWR sky130_fd_sc_hd__o211a_1
Xhold1049 _6844_/Q VGND VPWR _5277_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6965_ _7080_/CLK _6965_/D fanout479/X VGND VPWR _6965_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5916_ _6719_/Q _5642_/X _5666_/X _6634_/Q VGND VPWR _5916_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_179_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6896_ _7069_/CLK _6896_/D fanout482/X VGND VPWR _6896_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5847_ _6600_/Q _5616_/X _5648_/X _6605_/Q _5846_/X VGND VPWR _5852_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5778_ _5778_/A1 _6279_/S _5776_/X _5777_/X VGND VPWR _5778_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_166_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4729_ _4964_/A _4725_/Y _4728_/X _4229_/X VGND VPWR _4729_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_108_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold850 _6804_/Q VGND VPWR hold850/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold861 _5313_/X VGND VPWR _6876_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _7020_/Q VGND VPWR hold872/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _5424_/X VGND VPWR _6975_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _7032_/Q VGND VPWR hold894/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1550 _6641_/Q VGND VPWR _3168_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 _7159_/Q VGND VPWR _3912_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1572 _7116_/Q VGND VPWR _5887_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 _6412_/Q VGND VPWR _3852_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_426 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1594 _7176_/A VGND VPWR hold349/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_698 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_372 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6750_ _7006_/CLK _6750_/D fanout457/X VGND VPWR _6750_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3962_ _3962_/A _3962_/B VGND VPWR _6639_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_5701_ _6852_/Q _5648_/X _5666_/X _6892_/Q _5700_/X VGND VPWR _5706_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6681_ _6714_/CLK _6681_/D fanout470/X VGND VPWR _6681_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3893_ _5959_/A _5966_/A VGND VPWR _3893_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_31_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5632_ _5638_/A _5667_/B _5667_/C VGND VPWR _5632_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_148_158 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5563_ _7088_/Q _7089_/Q _5562_/D _7090_/Q VGND VPWR _5564_/C VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_144_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4514_ _4514_/A _4514_/B _4514_/C VGND VPWR _4518_/D VGND VPWR sky130_fd_sc_hd__and3_1
Xhold102 _3287_/Y VGND VPWR _3356_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _5452_/X VGND VPWR _7000_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ hold198/X _5494_/A1 _5495_/S VGND VPWR _5494_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold124 _3300_/Y VGND VPWR _3571_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold135 _6840_/Q VGND VPWR hold135/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold146 _5512_/X VGND VPWR _7053_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4556_/A _4611_/B VGND VPWR _5051_/A VGND VPWR sky130_fd_sc_hd__and2_2
Xhold157 _4030_/X VGND VPWR _6468_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _6783_/Q VGND VPWR hold168/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 _5519_/X VGND VPWR _7059_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_740 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7164_ net399_2/A _7164_/D _6394_/X VGND VPWR hold40/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4376_ _4376_/A _4376_/B _4568_/B VGND VPWR _4465_/B VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_86_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6115_ _6115_/A _6115_/B _6115_/C VGND VPWR _6126_/C VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_100_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3327_ hold47/X hold84/X VGND VPWR hold85/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7095_ _7113_/CLK _7095_/D fanout462/X VGND VPWR _7095_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_112_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6046_ _7020_/Q _5937_/X _5975_/D _6884_/Q _6029_/X VGND VPWR _6049_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3258_ _3259_/A1 hold93/A _3260_/S VGND VPWR _3258_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3189_ _7058_/Q VGND VPWR _3189_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_94_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6948_ _7065_/CLK _6948_/D fanout463/X VGND VPWR _6948_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6879_ _7078_/CLK _6879_/D fanout481/X VGND VPWR _6879_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_10_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_437 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold680 _5264_/X VGND VPWR _6833_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _5489_/X VGND VPWR _7033_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_484 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_735 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1380 _6531_/Q VGND VPWR _4117_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1391 _6654_/Q VGND VPWR _4255_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_760 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3219_/Y VGND VPWR mgmt_gpio_oeb[4] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput218 _7181_/X VGND VPWR mgmt_gpio_out[16] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput229 _7191_/X VGND VPWR mgmt_gpio_out[26] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4230_ _6640_/Q _4230_/B VGND VPWR _5006_/A VGND VPWR sky130_fd_sc_hd__nand2b_2
XFILLER_4_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4161_ hold736/X _6356_/A1 _4162_/S VGND VPWR _4161_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_122_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4092_ hold904/X _5509_/A1 _5202_/B VGND VPWR _4092_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6802_ _7051_/CLK _6802_/D fanout476/X VGND VPWR _6802_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_36_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4994_ _4413_/Y _4428_/Y _4621_/X VGND VPWR _4995_/C VGND VPWR sky130_fd_sc_hd__o21a_1
X_6733_ _3927_/A1 _6733_/D _6385_/X VGND VPWR _6733_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_3945_ input83/X _3945_/A1 _6403_/Q VGND VPWR _3945_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6664_ _6712_/CLK _6664_/D _6396_/A VGND VPWR _6664_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_31_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3876_ _6485_/Q _3867_/B _3875_/X _6487_/Q VGND VPWR _6485_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_176_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5615_ _7095_/Q _7094_/Q VGND VPWR _5657_/B VGND VPWR sky130_fd_sc_hd__and2b_2
X_6595_ _7137_/CLK _6595_/D VGND VPWR _6595_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_5546_ hold816/X _5546_/A1 _5549_/S VGND VPWR _5546_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_151_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5477_ hold455/X _5528_/A1 hold30/X VGND VPWR _5477_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4428_ _4753_/A _4607_/A _4600_/B VGND VPWR _4428_/Y VGND VPWR sky130_fd_sc_hd__nand3b_4
Xfanout401 hold60/X VGND VPWR _6357_/A1 VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_99_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xfanout412 _5526_/A1 VGND VPWR _5493_/A1 VGND VPWR sky130_fd_sc_hd__buf_4
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR net399_2/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_59_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout423 hold666/X VGND VPWR _5524_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_86_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout434 _5638_/A VGND VPWR _5664_/A VGND VPWR sky130_fd_sc_hd__buf_4
X_7147_ _3937_/A1 _7147_/D _6307_/B VGND VPWR _7147_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4359_ _4382_/B _4359_/B VGND VPWR _4359_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xfanout445 _6360_/A VGND VPWR fanout445/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_86_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout456 fanout466/X VGND VPWR fanout456/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout467 fanout469/X VGND VPWR _6383_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout478 fanout480/X VGND VPWR fanout478/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout489 _4625_/A VGND VPWR _4607_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_7078_ _7078_/CLK _7078_/D fanout485/X VGND VPWR _7078_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_104_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6029_ _7028_/Q _5944_/X _5975_/A _6844_/Q VGND VPWR _6029_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_100_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_481 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3730_ _3730_/A _3730_/B _3730_/C VGND VPWR _3762_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_13_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3661_ _3661_/A _3661_/B _3661_/C _3661_/D VGND VPWR _3661_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_5400_ _5400_/A hold17/X VGND VPWR _5408_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_6380_ _6401_/A _6401_/B VGND VPWR _6380_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_173_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3592_ _6877_/Q _5310_/A _5319_/A _6885_/Q VGND VPWR _3592_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_127_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5331_ hold868/X _5484_/A1 _5336_/S VGND VPWR _5331_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5262_ hold790/X _5538_/A1 _5264_/S VGND VPWR _5262_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_142 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_687 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7001_ _7001_/CLK _7001_/D fanout464/X VGND VPWR _7001_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_114_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4213_ hold447/X _6357_/A1 _4213_/S VGND VPWR _4213_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5193_ _5193_/A _5541_/B VGND VPWR _5201_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_4144_ hold944/X _5546_/A1 _4144_/S VGND VPWR _4144_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_498 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4075_ _6535_/Q hold94/X _4083_/S VGND VPWR hold95/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_4_0_csclk clkbuf_3_5_0_csclk/A VGND VPWR _6601_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_63_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4977_ _4631_/Y _4689_/B _4970_/Y VGND VPWR _4981_/B VGND VPWR sky130_fd_sc_hd__a21o_1
X_6716_ _7038_/CLK _6716_/D fanout455/X VGND VPWR _6716_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3928_ _6510_/Q _3268_/C _6406_/Q VGND VPWR _3928_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6647_ _6671_/CLK _6647_/D _6383_/A VGND VPWR _6647_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_20_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3859_ hold44/A _6488_/Q _3851_/C hold24/A VGND VPWR _3861_/A VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_137_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6578_ _6709_/CLK _6578_/D fanout445/X VGND VPWR _6578_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_124_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5529_ hold517/X _5538_/A1 _5531_/S VGND VPWR _5529_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_182_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_741 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_287 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_90 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4900_ _4900_/A _4900_/B VGND VPWR _4900_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_5880_ _6472_/Q _5627_/X _5635_/X _6567_/Q VGND VPWR _5880_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4831_ _4542_/D _4810_/B _4824_/X _4830_/X VGND VPWR _4831_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XANTENNA_180 _6542_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_191 _5494_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4762_ _4627_/A _4627_/B _4611_/Y _4581_/B _4542_/A VGND VPWR _4769_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_6501_ _6539_/CLK hold96/X fanout459/X VGND VPWR _7175_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3713_ input62/X _4102_/A _4244_/A _6646_/Q _3712_/X VGND VPWR _3720_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_4693_ _4881_/A _4630_/X _4753_/C _4975_/B _4689_/Y VGND VPWR _4693_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6432_ _6749_/CLK _6432_/D fanout449/X VGND VPWR _6432_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3644_ _6876_/Q _5310_/A _3964_/A _6420_/Q _3643_/X VGND VPWR _3651_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6363_ _6383_/A _6401_/B VGND VPWR _6363_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3575_ hold75/X _3692_/A VGND VPWR _5490_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_5314_ hold628/X _5509_/A1 _5318_/S VGND VPWR _5314_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6294_ _6684_/Q _5934_/X _5975_/B _6618_/Q _6293_/X VGND VPWR _6300_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5245_ hold920/X _5548_/A1 _5246_/S VGND VPWR _5245_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_741 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VPWR hold17/X VGND VPWR sky130_fd_sc_hd__buf_8
Xhold28 hold28/A VGND VPWR hold28/X VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_69_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold39 hold39/A VGND VPWR hold39/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ hold133/X hold60/X _5181_/S VGND VPWR _5176_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4127_ _4127_/A _6352_/B VGND VPWR _4132_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_83_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4058_ hold692/X _5509_/A1 _4058_/S VGND VPWR _4058_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VPWR _7140_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_24_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold509 _6633_/Q VGND VPWR hold509/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3360_ hold48/X hold75/A VGND VPWR hold49/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_111_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_624 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3291_ hold34/X VGND VPWR _3295_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_151_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5030_ _4542_/A _4902_/A _4628_/Y _4691_/A _4852_/X VGND VPWR _5131_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_25_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1209 _6794_/Q VGND VPWR _5221_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_744 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6981_ _6981_/CLK _6981_/D fanout463/X VGND VPWR _6981_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_93_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5932_ _7100_/Q _7099_/Q VGND VPWR _5981_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_53_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5863_ _3184_/Y _5651_/Y _5852_/Y _5862_/Y _5552_/B VGND VPWR _5863_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4814_ _4886_/B _4958_/B VGND VPWR _5089_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_5794_ _6968_/Q _5642_/X _5905_/A2 _6800_/Q _5793_/X VGND VPWR _5797_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4745_ _4456_/Y _4672_/B _4626_/Y _4639_/Y VGND VPWR _4768_/A VGND VPWR sky130_fd_sc_hd__o22a_1
X_4676_ _4737_/A _4676_/B VGND VPWR _5021_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_107_418 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6415_ _3945_/A1 _6415_/D _6371_/X VGND VPWR _6415_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3627_ input6/X _3365_/Y _3381_/Y input29/X _3626_/X VGND VPWR _3628_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6346_ _6345_/X _6346_/A1 _6346_/S VGND VPWR _7148_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3558_ hold35/X _3573_/B VGND VPWR _4274_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_0_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_335 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6277_ _6543_/Q _6226_/B _6276_/X VGND VPWR _6277_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
X_3489_ _3554_/A _3573_/B VGND VPWR _4232_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xinput107 wb_adr_i[17] VGND VPWR _4335_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput118 wb_adr_i[27] VGND VPWR input118/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5228_ hold687/X _5513_/A1 _5228_/S VGND VPWR _5228_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VPWR _4337_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_102_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5159_ hold553/X _6357_/A1 _5160_/S VGND VPWR _5159_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_112_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_0_csclk clkbuf_2_1_0_csclk/A VGND VPWR clkbuf_3_3_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XPHY_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_80 _6869_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_91 _6558_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_343 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_338 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_714 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4530_ _4413_/Y _4453_/B _4528_/X _4529_/Y VGND VPWR _4530_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_184_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold306 _5357_/X VGND VPWR _6915_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _4690_/B _4611_/B VGND VPWR _4902_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_171_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold317 _6558_/Q VGND VPWR hold317/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _5291_/X VGND VPWR _6857_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 _7182_/A VGND VPWR hold339/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _6200_/A _6200_/B _6200_/C _6200_/D VGND VPWR _6200_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_3412_ _3410_/Y _3449_/A1 _3829_/A VGND VPWR _3412_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7180_ _7180_/A VGND VPWR _7180_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4392_ _4566_/A _4564_/A _4392_/C VGND VPWR _4393_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_6131_ _7008_/Q _5958_/X _5978_/X _7000_/Q VGND VPWR _6131_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3343_ _3573_/A hold28/X VGND VPWR _5400_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_6062_ _6893_/Q _5946_/X _5955_/X _6805_/Q VGND VPWR _6062_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3274_ hold45/X _6720_/Q _3975_/S VGND VPWR hold46/A VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_100_616 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1006 _3355_/X VGND VPWR _5171_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 _6579_/Q VGND VPWR _4174_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5013_ _4619_/Y _4970_/Y _5010_/Y _4616_/Y _4796_/C VGND VPWR _5106_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold1028 _4199_/X VGND VPWR _6601_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1039 hold1598/X VGND VPWR _4061_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7006_/CLK _6964_/D fanout458/X VGND VPWR _6964_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_22_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5915_ _6469_/Q _5619_/X _5663_/X _6613_/Q _5914_/X VGND VPWR _5915_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6895_ _7076_/CLK _6895_/D fanout481/X VGND VPWR _6895_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5846_ _6466_/Q _5619_/X _5663_/X _6610_/Q VGND VPWR _5846_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5777_ _6507_/Q _7110_/Q _6103_/B1 VGND VPWR _5777_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_4728_ _5039_/A _4964_/A _4727_/X VGND VPWR _4728_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_135_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_524 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_630 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4659_ _4846_/B _4644_/Y _4646_/Y _4657_/X _4658_/X VGND VPWR _4660_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_190_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold840 _7035_/Q VGND VPWR hold840/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _5232_/X VGND VPWR _6804_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold862 _6900_/Q VGND VPWR hold862/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _5475_/X VGND VPWR _7020_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _6736_/Q VGND VPWR hold884/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _6642_/Q _6329_/A2 _6329_/B1 _4230_/B VGND VPWR _6329_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold895 _5488_/X VGND VPWR _7032_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1540 _6351_/X VGND VPWR _7150_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 _4231_/X VGND VPWR _6624_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 _7113_/Q VGND VPWR _5821_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1573 _6761_/Q VGND VPWR hold129/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_177_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1584 _7197_/A VGND VPWR hold237/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1595 _6725_/Q VGND VPWR _5113_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_192 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7069_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_67_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_47_csclk _7001_/CLK VGND VPWR _6997_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_57_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3961_ _6644_/Q _3961_/B VGND VPWR _6636_/D VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_16_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5700_ _6900_/Q _5621_/X _5658_/X _6884_/Q VGND VPWR _5700_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_189_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6680_ _6683_/CLK _6680_/D _6390_/A VGND VPWR _6680_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3892_ _5600_/A _7102_/Q VGND VPWR _5966_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_5631_ _5664_/A _5658_/B _5657_/B VGND VPWR _5631_/X VGND VPWR sky130_fd_sc_hd__and3b_4
X_5562_ _7088_/Q _7089_/Q _7090_/Q _5562_/D VGND VPWR _5564_/B VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_191_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4513_ _4902_/A _4453_/B _4542_/A VGND VPWR _4514_/C VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_144_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold103 _3511_/A VGND VPWR _3717_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_5493_ _5493_/A0 _5493_/A1 _5495_/S VGND VPWR _5493_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold114 _6928_/Q VGND VPWR hold114/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold125 hold125/A VGND VPWR _3562_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_144_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold136 _5272_/X VGND VPWR _6840_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _4607_/A _4753_/A VGND VPWR _4993_/A VGND VPWR sky130_fd_sc_hd__nand2b_4
Xhold147 _6982_/Q VGND VPWR hold147/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A VGND VPWR hold158/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 _5208_/X VGND VPWR _6783_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ net399_2/A _7163_/D _6393_/X VGND VPWR hold58/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4375_ _4334_/B _4334_/C _4374_/A _4372_/X VGND VPWR _4568_/B VGND VPWR sky130_fd_sc_hd__a31o_2
X_6114_ _6983_/Q _5945_/X _5975_/C _6839_/Q _6113_/X VGND VPWR _6115_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3326_ _3562_/A _3714_/A VGND VPWR _3326_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
X_7094_ _7113_/CLK _7094_/D fanout462/X VGND VPWR _7094_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_86_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6045_ _7065_/Q _5934_/X _5975_/B _6868_/Q _6044_/X VGND VPWR _6045_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3257_ hold93/A _3257_/A1 _3260_/S VGND VPWR _3257_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3188_ _7066_/Q VGND VPWR _3188_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_54_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6947_ _7011_/CLK hold10/X fanout456/X VGND VPWR _6947_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_6878_ _7051_/CLK _6878_/D fanout476/X VGND VPWR _6878_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_50_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5829_ _6460_/Q _5624_/X _5654_/X _6675_/Q _5822_/Y VGND VPWR _5829_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_660 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold670 _5299_/X VGND VPWR _6864_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _6889_/Q VGND VPWR hold681/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 hold692/A VGND VPWR hold692/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1370 hold1370/A VGND VPWR wb_dat_o[3] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_18_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1381 _6526_/Q VGND VPWR _4112_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_330 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1392 _4255_/X VGND VPWR hold61/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_706 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput208 _3218_/Y VGND VPWR mgmt_gpio_oeb[5] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput219 _7182_/X VGND VPWR mgmt_gpio_out[17] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_99_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_614 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4160_ _4160_/A0 _5493_/A1 _4162_/S VGND VPWR _4160_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4091_ _4091_/A0 _4090_/X _4101_/S VGND VPWR _4091_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6801_ _7053_/CLK _6801_/D fanout459/X VGND VPWR _6801_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4993_ _4993_/A _4993_/B VGND VPWR _5069_/C VGND VPWR sky130_fd_sc_hd__nand2_1
X_6732_ _3945_/A1 _6732_/D _6384_/X VGND VPWR _6732_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_3944_ _6404_/Q _3946_/B VGND VPWR _3944_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_176_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6663_ _7058_/CLK _6663_/D _6396_/A VGND VPWR _6663_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_177_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3875_ _7167_/Q _3875_/B _3875_/C VGND VPWR _3875_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_137_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5614_ _5638_/A _5667_/B _5666_/B VGND VPWR _5614_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_6594_ _7130_/CLK _6594_/D VGND VPWR _6594_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_117_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5545_ _5545_/A0 _5545_/A1 _5549_/S VGND VPWR _5545_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_652 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_0_0_csclk clkbuf_3_1_0_csclk/A VGND VPWR clkbuf_3_0_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
X_5476_ _5476_/A0 _5545_/A1 hold30/X VGND VPWR _5476_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4427_ _4561_/B _4632_/B VGND VPWR _4992_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xfanout402 hold59/X VGND VPWR hold60/A VGND VPWR sky130_fd_sc_hd__buf_12
Xfanout413 hold6/X VGND VPWR _5526_/A1 VGND VPWR sky130_fd_sc_hd__buf_8
X_7146_ _3937_/A1 _7146_/D _6307_/B VGND VPWR hold52/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xfanout424 hold666/X VGND VPWR hold667/A VGND VPWR sky130_fd_sc_hd__buf_8
X_4358_ _4739_/A _4356_/B _4357_/B _4661_/A VGND VPWR _4359_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_1
Xfanout435 _5899_/B VGND VPWR _5638_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_101_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xfanout446 fanout486/X VGND VPWR _6360_/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_86_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout457 fanout466/X VGND VPWR fanout457/X VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout468 fanout469/X VGND VPWR fanout468/X VGND VPWR sky130_fd_sc_hd__buf_4
X_3309_ hold27/X hold65/X VGND VPWR _3370_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7077_ _7086_/CLK _7077_/D fanout483/X VGND VPWR _7077_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_86_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout479 fanout480/X VGND VPWR fanout479/X VGND VPWR sky130_fd_sc_hd__buf_8
X_4289_ hold519/X _5544_/A1 _4291_/S VGND VPWR _4289_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6028_ _6028_/A0 _6027_/X _6279_/S VGND VPWR _6028_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_73_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3660_ _7073_/Q _5532_/A _5148_/A _6739_/Q _3659_/X VGND VPWR _3661_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3591_ _6617_/Q _4214_/A _4238_/A _6633_/Q VGND VPWR _3591_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5330_ hold549/X _5543_/A1 _5336_/S VGND VPWR _5330_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_127_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5261_ hold190/X _5519_/A1 _5264_/S VGND VPWR _5261_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7000_ _7017_/CLK _7000_/D fanout461/X VGND VPWR _7000_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_141_154 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4212_ hold493/X _5518_/A1 _4213_/S VGND VPWR _4212_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5192_ hold423/X _5534_/A1 _5192_/S VGND VPWR _5192_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4143_ hold505/X _5518_/A1 _4144_/S VGND VPWR _4143_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4074_ hold170/X _4073_/X _4084_/S VGND VPWR _4074_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_64_661 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4976_ _4576_/Y _4701_/Y _4975_/Y _4613_/Y VGND VPWR _4981_/A VGND VPWR sky130_fd_sc_hd__o22a_1
X_6715_ _7038_/CLK _6715_/D fanout455/X VGND VPWR _6715_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_20_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3927_ _6511_/Q _3927_/A1 _6405_/Q VGND VPWR _3927_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_165_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_714 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6646_ _6671_/CLK _6646_/D fanout468/X VGND VPWR _6646_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3858_ _3858_/A1 _3851_/C _3857_/X VGND VPWR _6410_/D VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_109_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6577_ _7140_/CLK _6577_/D VGND VPWR _6577_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3789_ _5186_/A _3355_/X _3788_/Y hold49/A _7026_/Q VGND VPWR _3789_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_3_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5528_ hold435/X _5528_/A1 _5531_/S VGND VPWR _5528_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5459_ hold110/X hold60/X _5461_/S VGND VPWR _5459_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7129_ _7130_/CLK _7129_/D fanout486/X VGND VPWR _7129_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_19_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_474 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_385 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4830_ _4542_/A _4810_/B _4821_/X _4828_/X _4829_/X VGND VPWR _4830_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_170 _4108_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_181 _6925_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_192 _5544_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4761_ _4627_/A _4615_/Y _4626_/Y _4810_/A _4672_/B VGND VPWR _4772_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_6500_ _6539_/CLK _6500_/D fanout461/X VGND VPWR _7174_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3712_ _7019_/Q hold29/A _5256_/A _6827_/Q VGND VPWR _3712_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4692_ _4975_/B VGND VPWR _4692_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_119_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6431_ _6749_/CLK _6431_/D fanout449/X VGND VPWR _6431_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3643_ _6972_/Q _5418_/A _4058_/S input45/X VGND VPWR _3643_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_134_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6362_ _6400_/A _6400_/B VGND VPWR _6362_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3574_ _6990_/Q _5436_/A _4304_/A _6699_/Q VGND VPWR _3574_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5313_ hold860/X _5484_/A1 _5318_/S VGND VPWR _5313_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6293_ _6704_/Q _5971_/A _5979_/X _6474_/Q VGND VPWR _6293_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5244_ hold764/X _5538_/A1 _5246_/S VGND VPWR _5244_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_316 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold18 hold18/A VGND VPWR hold18/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A VGND VPWR hold29/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5182_/S hold17/X VGND VPWR _5181_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_84_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4126_ hold555/X _5513_/A1 _4126_/S VGND VPWR _4126_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_17 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4057_ hold89/X _4056_/X _4067_/S VGND VPWR hold90/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_631 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4959_ _4959_/A _4959_/B VGND VPWR _4959_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_177_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6629_ _6629_/CLK _6629_/D _6390_/A VGND VPWR _6629_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_180_503 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3290_ _3975_/S hold33/X VGND VPWR hold34/A VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_111_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6980_ _7065_/CLK _6980_/D fanout465/X VGND VPWR _6980_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_53_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5931_ _7118_/Q _6279_/S _5929_/X _5930_/X VGND VPWR _7118_/D VGND VPWR sky130_fd_sc_hd__o22a_1
X_5862_ _5862_/A _5862_/B _5862_/C _5862_/D VGND VPWR _5862_/Y VGND VPWR sky130_fd_sc_hd__nor4_2
XFILLER_33_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4813_ _4813_/A _4959_/B VGND VPWR _4958_/B VGND VPWR sky130_fd_sc_hd__and2_1
X_5793_ _6872_/Q _5628_/X _5643_/X _7000_/Q VGND VPWR _5793_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_21_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4744_ _4542_/B _4581_/B _4611_/Y _4619_/Y VGND VPWR _4771_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_159_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4675_ _4565_/X _4741_/A _4609_/Y _4663_/Y _5002_/A VGND VPWR _4682_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6414_ _3568_/A1 _6414_/D _6370_/X VGND VPWR _6414_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3626_ _6688_/Q _4292_/A _4032_/A _6473_/Q VGND VPWR _3626_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6345_ _6642_/Q _6345_/A2 _6345_/B1 _6350_/A2 _6344_/X VGND VPWR _6345_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3557_ _6694_/Q _4298_/A _4268_/A _6669_/Q _3556_/X VGND VPWR _3565_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6276_ _6267_/X _6301_/C _6276_/C _6276_/D VGND VPWR _6276_/X VGND VPWR sky130_fd_sc_hd__and4b_2
XFILLER_142_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3488_ _3487_/X _3488_/A1 _3829_/B VGND VPWR _3488_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput108 wb_adr_i[18] VGND VPWR _4335_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5227_ hold722/X _5521_/A1 _5227_/S VGND VPWR _5227_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput119 wb_adr_i[28] VGND VPWR input119/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5158_ hold754/X _6356_/A1 _5160_/S VGND VPWR _5158_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4109_ _6396_/B hold37/X _5505_/B VGND VPWR hold38/A VGND VPWR sky130_fd_sc_hd__and3b_4
X_5089_ _5089_/A _5089_/B _5089_/C _5089_/D VGND VPWR _5122_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_71_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_491 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_511 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_70 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_81 _6619_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_92 _6558_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_369 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_73 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4460_ _4460_/A _4993_/A VGND VPWR _4782_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold307 _6937_/Q VGND VPWR hold307/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold318 _4149_/X VGND VPWR _6558_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 _6897_/Q VGND VPWR hold329/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _7170_/Q _6487_/Q VGND VPWR _3829_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_4391_ _4564_/A _4392_/C _4566_/A VGND VPWR _4393_/A VGND VPWR sky130_fd_sc_hd__a21oi_1
X_6130_ _6864_/Q _5943_/X _5981_/X _6920_/Q VGND VPWR _6130_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3342_ hold27/X _3454_/B VGND VPWR hold28/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_98_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_590 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6061_ _6941_/Q _5961_/X _6055_/X _6060_/X VGND VPWR _6066_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_97_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3273_ hold44/X _3251_/A _6488_/Q VGND VPWR hold45/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_112_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_628 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1007 _5164_/X VGND VPWR _5165_/S VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5012_ _4689_/B _4970_/Y _5010_/Y _4628_/Y _4796_/A VGND VPWR _5134_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold1018 _4174_/X VGND VPWR _6579_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 _6466_/Q VGND VPWR _4028_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6963_ _6963_/CLK hold14/X fanout458/X VGND VPWR _6963_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5914_ _6549_/Q _5655_/X _5912_/X _5913_/X VGND VPWR _5914_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_6894_ _7051_/CLK _6894_/D fanout476/X VGND VPWR _6894_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5845_ _6646_/Q _5621_/X _5628_/X _6615_/Q _5844_/X VGND VPWR _5852_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5776_ _6791_/Q _5652_/Y _5769_/X _5775_/X _6303_/S VGND VPWR _5776_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_175_650 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4727_ _4500_/A _4611_/Y _4964_/B _5039_/B VGND VPWR _4727_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_175_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4658_ _5088_/A _5099_/B _4658_/C VGND VPWR _4658_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_174_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput90 spimemio_flash_io2_oeb VGND VPWR input90/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold830 _6664_/Q VGND VPWR hold830/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3609_ _6622_/Q _4220_/A _4151_/A _6563_/Q VGND VPWR _3609_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold841 _5492_/X VGND VPWR _7035_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold852 _6749_/Q VGND VPWR hold852/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4589_ _4589_/A _4589_/B _4589_/C _4589_/D VGND VPWR _4589_/Y VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_103_400 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold863 _5340_/X VGND VPWR _6900_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _6916_/Q VGND VPWR hold874/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _6327_/X _6328_/A1 _6346_/S VGND VPWR _7142_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold885 _5147_/X VGND VPWR _6736_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _6885_/Q VGND VPWR hold896/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6259_ _6688_/Q _5961_/X _6257_/X _6258_/X VGND VPWR _6264_/A VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_67_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1530 _7104_/Q VGND VPWR _5607_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1541 _6723_/Q VGND VPWR _5061_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _7117_/Q VGND VPWR _5909_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 _7091_/Q VGND VPWR _3176_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_715 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1574 _7168_/Q VGND VPWR _3249_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1585 _6527_/Q VGND VPWR hold692/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1596 _6536_/Q VGND VPWR hold158/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_672 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_355 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3960_ _6769_/Q _3960_/B VGND VPWR _3960_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3891_ _5978_/A _5969_/A VGND VPWR _5959_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_149_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5630_ _5664_/A _5658_/B _5666_/B VGND VPWR _5630_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_31_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5561_ _5561_/A1 _5554_/Y _5604_/B _5560_/X VGND VPWR _7089_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4512_ _4947_/B _4947_/C _4456_/Y VGND VPWR _4514_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_156_171 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5492_ hold840/X _5492_/A1 _5495_/S VGND VPWR _5492_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_156_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold104 _3372_/Y VGND VPWR _3990_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _5371_/X VGND VPWR _6928_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold126 _3326_/Y VGND VPWR _5220_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4607_/A _4753_/A VGND VPWR _4611_/B VGND VPWR sky130_fd_sc_hd__and2b_4
Xhold137 _6960_/Q VGND VPWR hold137/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold148 _5432_/X VGND VPWR _6982_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _4123_/X VGND VPWR _6536_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ net399_2/A _7162_/D _6392_/X VGND VPWR hold93/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4374_ _4374_/A _4374_/B VGND VPWR _4471_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_6113_ _6927_/Q _5938_/X _5952_/X _6959_/Q VGND VPWR _6113_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3325_ _3379_/A _3543_/A VGND VPWR _5418_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_7093_ _7113_/CLK _7093_/D fanout462/X VGND VPWR _7093_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_86_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6044_ _7049_/Q _5971_/A _5979_/X _6988_/Q VGND VPWR _6044_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3256_ _3257_/A1 _3256_/A1 _3260_/S VGND VPWR _7164_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_447 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3187_ _7074_/Q VGND VPWR _3187_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_54_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6946_ _7049_/CLK _6946_/D fanout457/X VGND VPWR _6946_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_81_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6877_ _7076_/CLK _6877_/D fanout481/X VGND VPWR _6877_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5828_ _6475_/Q _5630_/X _5824_/X _5825_/X _5827_/X VGND VPWR _5828_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
X_5759_ _7007_/Q _5625_/X _5661_/X _6879_/Q VGND VPWR _5759_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_185_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_420 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold660 _6793_/Q VGND VPWR hold660/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 _6832_/Q VGND VPWR hold671/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold682 _5327_/X VGND VPWR _6889_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _4113_/X VGND VPWR _6527_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1360 hold1360/A VGND VPWR wb_dat_o[20] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_94_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1371 _4188_/A1 VGND VPWR hold1371/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_139 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1382 _4112_/X VGND VPWR hold7/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _7041_/Q VGND VPWR _5499_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput209 _3217_/Y VGND VPWR mgmt_gpio_oeb[6] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_5_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_696 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_185 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4090_ _5205_/A0 _5484_/A1 _5202_/B VGND VPWR _4090_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_128 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6800_ _6920_/CLK _6800_/D fanout474/X VGND VPWR _6800_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_91_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4992_ _4992_/A _4992_/B VGND VPWR _4996_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_6731_ _3945_/A1 _6731_/D _6383_/X VGND VPWR _6731_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_3943_ input84/X _3268_/C _6404_/Q VGND VPWR _3943_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_149_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6662_ _7058_/CLK _6662_/D _6396_/A VGND VPWR _6662_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3874_ _7104_/Q _6757_/Q _6762_/Q VGND VPWR _5606_/A VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_177_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5613_ _7095_/Q _7094_/Q VGND VPWR _5666_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_6593_ _7130_/CLK _6593_/D VGND VPWR _6593_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_191_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5544_ hold215/X _5544_/A1 _5549_/S VGND VPWR _5544_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5475_ hold872/X _5484_/A1 hold30/X VGND VPWR _5475_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_144_163 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4426_ _4753_/A _4607_/A VGND VPWR _4632_/B VGND VPWR sky130_fd_sc_hd__nand2b_4
Xfanout403 _5519_/A1 VGND VPWR _5546_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_160_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout414 _5544_/A1 VGND VPWR _5484_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_7145_ _3937_/A1 _7145_/D _6307_/B VGND VPWR _7145_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_113_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout425 hold666/X VGND VPWR _5473_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_4357_ _4642_/A _4357_/B VGND VPWR _4382_/B VGND VPWR sky130_fd_sc_hd__xnor2_1
Xfanout436 _7096_/Q VGND VPWR _5899_/B VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout447 fanout450/X VGND VPWR fanout447/X VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout458 fanout466/X VGND VPWR fanout458/X VGND VPWR sky130_fd_sc_hd__buf_8
X_3308_ _3453_/A hold64/X VGND VPWR hold65/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_100_222 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout469 fanout486/X VGND VPWR fanout469/X VGND VPWR sky130_fd_sc_hd__buf_6
X_7076_ _7076_/CLK _7076_/D fanout481/X VGND VPWR _7076_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4288_ hold269/X _5534_/A1 _4291_/S VGND VPWR _4288_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3239_ _3837_/A _3239_/B VGND VPWR _3875_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_46_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6027_ _7119_/Q _6026_/X _6303_/S VGND VPWR _6027_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6929_ _7054_/CLK _6929_/D fanout461/X VGND VPWR _6929_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7085_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_168_723 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_csclk _7001_/CLK VGND VPWR _7065_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_182_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_664 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold490 _5363_/X VGND VPWR _6921_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VPWR clkbuf_1_0_1_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_104_594 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1190 _6353_/X VGND VPWR _7151_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3590_ _6837_/Q _5265_/A _4172_/A _6581_/Q VGND VPWR _3590_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_127_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5260_ hold652/X _5509_/A1 _5264_/S VGND VPWR _5260_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_48_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4211_ _4211_/A0 _5493_/A1 _4213_/S VGND VPWR _4211_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5191_ _5191_/A0 hold667/X _5192_/S VGND VPWR _5191_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_710 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4142_ _4142_/A0 _5493_/A1 _4144_/S VGND VPWR _4142_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4073_ hold401/X hold6/X _4083_/S VGND VPWR _4073_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4975_ _4975_/A _4975_/B VGND VPWR _4975_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_149_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6714_ _6714_/CLK _6714_/D fanout470/X VGND VPWR _6714_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3926_ _6512_/Q _3251_/A _6406_/Q VGND VPWR _3926_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6645_ _6671_/CLK _6645_/D fanout468/X VGND VPWR _6645_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3857_ hold81/A _6488_/Q _3850_/Y _3856_/X _3866_/S VGND VPWR _3857_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_428 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6576_ _7140_/CLK _6576_/D VGND VPWR _6576_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3788_ _3788_/A VGND VPWR _3788_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_117_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5527_ _5527_/A0 _5545_/A1 _5531_/S VGND VPWR _5527_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_133_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5458_ _5458_/A0 _5494_/A1 _5462_/S VGND VPWR _5458_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4409_ _4551_/A _4570_/A _4459_/B VGND VPWR _4584_/A VGND VPWR sky130_fd_sc_hd__and3_1
X_5389_ hold149/X hold99/X _5390_/S VGND VPWR _5389_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7128_ _7130_/CLK _7128_/D fanout486/X VGND VPWR _7128_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7083_/CLK _7059_/D _6396_/A VGND VPWR _7059_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_131_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_486 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_160 hold666/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_171 _5291_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_182 _7066_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_687 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_193 _5465_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4760_ _4948_/A _4672_/B _4626_/Y _4653_/Y VGND VPWR _5003_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_193_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3711_ _6435_/Q _3372_/Y _5319_/A _6883_/Q _3710_/X VGND VPWR _3720_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4691_ _4691_/A _4902_/B VGND VPWR _4975_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_6430_ _6749_/CLK _6430_/D fanout449/X VGND VPWR _6430_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3642_ _3641_/X _3642_/A1 _3829_/B VGND VPWR _3642_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_174_556 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6361_ _6400_/A _6400_/B VGND VPWR _6361_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3573_ _3573_/A _3573_/B VGND VPWR _4304_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_114_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5312_ hold541/X _5543_/A1 _5318_/S VGND VPWR _5312_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6292_ _6564_/Q _5953_/X _5960_/X _6674_/Q _6291_/X VGND VPWR _6292_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5243_ hold196/X _5519_/A1 _5246_/S VGND VPWR _5243_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_328 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold19 hold19/A VGND VPWR hold19/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ hold48/X _3717_/B hold667/X _5173_/X hold16/X VGND VPWR _5174_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_68_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4125_ _4125_/A0 hold99/X _4126_/S VGND VPWR _4125_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4056_ _4112_/A0 hold6/X _4058_/S VGND VPWR _4056_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4958_ _5042_/B _4958_/B VGND VPWR _5046_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_184_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3909_ _3909_/A _3909_/B VGND VPWR _3910_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_177_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4889_ _4689_/A _4645_/Y _4892_/B _4491_/Y _4523_/Y VGND VPWR _5084_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_137_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6628_ _6683_/CLK _6628_/D _6390_/A VGND VPWR _6628_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_137_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_450 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6559_ _6629_/CLK _6559_/D _6390_/A VGND VPWR _6559_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5930_ _5552_/B _7117_/Q _6103_/B1 VGND VPWR _5930_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_5861_ _6471_/Q _5627_/X _5655_/X _6546_/Q _5860_/X VGND VPWR _5862_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4812_ _4562_/Y _4810_/B _4948_/D VGND VPWR _4812_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_5792_ _6984_/Q _5624_/X _5818_/A2 _6824_/Q _5791_/X VGND VPWR _5797_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4743_ _4810_/A _4581_/B _4611_/Y _4613_/Y VGND VPWR _4772_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_187_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4674_ _4608_/X _4644_/B _4984_/B _4673_/Y _4472_/A VGND VPWR _4674_/Y VGND VPWR
+ sky130_fd_sc_hd__a2111oi_1
X_6413_ _3568_/A1 _6413_/D _6369_/X VGND VPWR hold32/A VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_135_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3625_ _6437_/Q _3372_/Y _3964_/A _6421_/Q _3624_/X VGND VPWR _3628_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_431 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6344_ _6644_/Q _6344_/A2 _6344_/B1 _6643_/Q VGND VPWR _6344_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3556_ _7022_/Q hold29/A _4238_/A _6634_/Q VGND VPWR _3556_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_88_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6275_ _6275_/A _6275_/B _6275_/C _6275_/D VGND VPWR _6276_/D VGND VPWR sky130_fd_sc_hd__nor4_1
X_3487_ _3486_/Y _6731_/Q _3829_/A VGND VPWR _3487_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput109 wb_adr_i[19] VGND VPWR _4335_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5226_ _5226_/A0 _5538_/A1 _5227_/S VGND VPWR _5226_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_69_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5157_ hold950/X _6355_/A1 _5160_/S VGND VPWR _5157_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4108_ hold383/X _5538_/A1 _4108_/S VGND VPWR _4108_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5088_ _5088_/A _5088_/B _5088_/C _5088_/D VGND VPWR _5089_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_56_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_278 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4039_ _4039_/A0 _5491_/A1 _4043_/S VGND VPWR _4039_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_440 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_60 _6025_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_71 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_82 _6898_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_126_718 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_93 _6568_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold308 _5381_/X VGND VPWR _6937_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold319 _7061_/Q VGND VPWR hold319/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_559 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3410_ _3410_/A _3410_/B VGND VPWR _3410_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4390_ _4631_/D _4633_/B _4661_/A _4441_/B VGND VPWR _4392_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_125_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3341_ hold36/X hold85/X VGND VPWR hold86/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_98_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6060_ _7013_/Q _5940_/X _5967_/X _6853_/Q _6054_/X VGND VPWR _6060_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3272_ hold25/X _4885_/B2 _3975_/S VGND VPWR hold26/A VGND VPWR sky130_fd_sc_hd__mux2_2
Xhold1008 _5165_/X VGND VPWR _6750_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _4689_/A _4644_/Y _5010_/Y _4639_/Y VGND VPWR _5011_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_112_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1019 _6546_/Q VGND VPWR _4135_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_278 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6962_ _7006_/CLK _6962_/D fanout457/X VGND VPWR _6962_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_53_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5913_ _6603_/Q _5616_/X _5913_/B1 _6554_/Q VGND VPWR _5913_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6893_ _7076_/CLK _6893_/D fanout481/X VGND VPWR _6893_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_34_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5844_ _6456_/Q _5645_/X _5910_/B1 _6626_/Q VGND VPWR _5844_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5775_ _6935_/Q _5654_/X _5770_/X _5772_/X _5774_/X VGND VPWR _5775_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_4726_ _4984_/A _4965_/B _4975_/A VGND VPWR _5039_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_175_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4657_ _4611_/Y _4639_/Y _4652_/Y _4620_/Y VGND VPWR _4657_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xinput80 spi_sck VGND VPWR input80/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold820 _6623_/Q VGND VPWR hold820/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3608_ input55/X _5193_/A _4256_/A _6658_/Q _3589_/X VGND VPWR _3611_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput91 spimemio_flash_io3_do VGND VPWR input91/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold831 _4267_/X VGND VPWR _6664_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _4948_/B _4672_/B VGND VPWR _4588_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold842 _6629_/Q VGND VPWR hold842/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold853 _5163_/X VGND VPWR _6749_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _6932_/Q VGND VPWR hold864/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6327_ _6644_/Q _6327_/A2 _6327_/B1 _6350_/A2 _6326_/X VGND VPWR _6327_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xmgmt_gpio_15_buff_inst _3936_/X VGND VPWR mgmt_gpio_out[15] VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold875 _5358_/X VGND VPWR _6916_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ hold74/X _3571_/B VGND VPWR _6352_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_412 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold886 _6444_/Q VGND VPWR hold886/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _5323_/X VGND VPWR _6885_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6258_ _6478_/Q _5940_/X _5967_/X _6607_/Q _6256_/X VGND VPWR _6258_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5209_ hold291/X _5521_/A1 _5210_/S VGND VPWR _5209_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_190_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6189_ _6189_/A _6189_/B _6189_/C VGND VPWR _6189_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
Xhold1520 _7110_/Q VGND VPWR _5757_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 hold52/A VGND VPWR _6340_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _6640_/Q VGND VPWR _3954_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 _7114_/Q VGND VPWR _5843_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1564 _7126_/Q VGND VPWR _6179_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 _7087_/Q VGND VPWR _5551_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 _7098_/Q VGND VPWR _5590_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 _6784_/Q VGND VPWR hold291/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_646 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3890_ _7100_/Q _7099_/Q VGND VPWR _5969_/A VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_149_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5560_ _7088_/Q _7089_/Q _6509_/Q _5552_/B _3885_/Y VGND VPWR _5560_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_163_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4511_ _4453_/B _4948_/C _4508_/X _4510_/X VGND VPWR _4514_/A VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_157_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5491_ _5491_/A0 _5491_/A1 _5495_/S VGND VPWR _5491_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold105 _3997_/X VGND VPWR _6440_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 _6942_/Q VGND VPWR hold116/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _4465_/B _4900_/A _4896_/B _4724_/A VGND VPWR _4442_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
Xhold127 _5227_/S VGND VPWR _5228_/S VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _5407_/X VGND VPWR _6960_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _6944_/Q VGND VPWR hold149/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7161_ net399_2/A _7161_/D _6391_/X VGND VPWR _7161_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_113_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4373_ _4702_/B _4434_/B VGND VPWR _4627_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_171_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6112_ _6975_/Q _5947_/X _5965_/X _6799_/Q _6111_/X VGND VPWR _6115_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3324_ _3356_/A hold73/X VGND VPWR _3543_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7092_ _7113_/CLK _7092_/D fanout462/X VGND VPWR _7092_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6043_ _6820_/Q _5953_/X _5960_/X _7073_/Q _6042_/X VGND VPWR _6043_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3255_ _3256_/A1 _3255_/A1 _3260_/S VGND VPWR _7165_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3186_ _7082_/Q VGND VPWR _3186_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6945_ _7054_/CLK _6945_/D fanout461/X VGND VPWR _6945_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_35_760 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A VGND VPWR clkbuf_3_5_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6876_ _7067_/CLK _6876_/D fanout476/X VGND VPWR _6876_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_167_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5827_ _6578_/Q _5928_/A2 _5913_/B1 _6550_/Q _5826_/X VGND VPWR _5827_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5758_ _3226_/Y _5899_/B _5651_/B VGND VPWR _5758_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_147_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4709_ _4691_/A _4902_/B _4619_/Y VGND VPWR _5084_/C VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_135_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5689_ _6939_/Q _5632_/X _5663_/X _6859_/Q _5688_/X VGND VPWR _5690_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold650 _7054_/Q VGND VPWR hold650/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _5219_/X VGND VPWR _6793_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold672 _5263_/X VGND VPWR _6832_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xmax_cap391 _4230_/B VGND VPWR _6350_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold683 _6791_/Q VGND VPWR hold683/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _6935_/Q VGND VPWR hold694/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_242 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_159 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1350 hold1350/A VGND VPWR wb_dat_o[27] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1361 _6313_/A1 VGND VPWR hold1361/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1372 hold1372/A VGND VPWR wb_dat_o[0] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_85_693 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1383 hold1578/X VGND VPWR _4125_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 _5499_/X VGND VPWR hold3/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_107 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4991_ _4626_/Y _4644_/Y _4646_/Y VGND VPWR _4991_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_91_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6730_ _3945_/A1 _6730_/D _6382_/X VGND VPWR _6730_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_189_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3942_ _3975_/S _3942_/A2 _6396_/B _3941_/Y VGND VPWR _3942_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_149_415 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6661_ _6712_/CLK _6661_/D _6396_/A VGND VPWR _6661_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3873_ _3264_/B _3838_/A _3872_/X _3832_/B _6402_/Q VGND VPWR _6402_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5612_ _5552_/B _5606_/A _5610_/Y VGND VPWR _6304_/S VGND VPWR sky130_fd_sc_hd__a21o_2
X_6592_ _7130_/CLK _6592_/D VGND VPWR _6592_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_191_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5543_ hold644/X _5543_/A1 _5549_/S VGND VPWR _5543_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5474_ hold594/X _5543_/A1 hold30/X VGND VPWR _5474_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4425_ _4685_/A _4921_/A VGND VPWR _5023_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_144_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_668 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout404 _5519_/A1 VGND VPWR _5528_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_7144_ _3937_/A1 _7144_/D fanout487/X VGND VPWR _7144_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4356_ _4356_/A _4356_/B VGND VPWR _4492_/D VGND VPWR sky130_fd_sc_hd__nor2_2
Xfanout415 hold6/X VGND VPWR _5544_/A1 VGND VPWR sky130_fd_sc_hd__buf_8
Xfanout426 hold665/X VGND VPWR hold666/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_48_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout437 _3963_/S VGND VPWR _3975_/S VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xfanout448 fanout450/X VGND VPWR fanout448/X VGND VPWR sky130_fd_sc_hd__buf_4
X_3307_ _3586_/A _3374_/A VGND VPWR _5355_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_113_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout459 fanout462/X VGND VPWR fanout459/X VGND VPWR sky130_fd_sc_hd__buf_8
X_7075_ _7083_/CLK _7075_/D _6396_/A VGND VPWR _7075_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4287_ _4287_/A0 hold667/X _4291_/S VGND VPWR _4287_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6026_ _6014_/Y _6025_/X _6787_/Q _6226_/B VGND VPWR _6026_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3238_ _6416_/Q _3837_/A _6485_/Q _3829_/A _3239_/B VGND VPWR _3249_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_100_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3169_ _6642_/Q VGND VPWR _3962_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_64_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_376 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6928_ _7017_/CLK _6928_/D fanout461/X VGND VPWR _6928_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_23_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_735 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6859_ _7011_/CLK _6859_/D fanout456/X VGND VPWR _6859_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_168_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_676 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold480 _5333_/X VGND VPWR _6894_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _6648_/Q VGND VPWR hold491/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1180 _5293_/X VGND VPWR _6858_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 _6922_/Q VGND VPWR _5365_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_200 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4210_ _4210_/A0 _5492_/A1 _4213_/S VGND VPWR _4210_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5190_ _5190_/A _5190_/B hold16/X VGND VPWR _5192_/S VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_68_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4141_ _4141_/A0 _5492_/A1 _4144_/S VGND VPWR _4141_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4072_ _4072_/A0 _4071_/X _4084_/S VGND VPWR _4072_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4974_ _5021_/B _4974_/B _5008_/C _4974_/D VGND VPWR _4983_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_51_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6713_ _7083_/CLK _6713_/D _6396_/A VGND VPWR _6713_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3925_ _6521_/Q input81/X _3957_/B VGND VPWR _3925_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_20_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6644_ _3937_/A1 _6644_/D fanout487/X VGND VPWR _6644_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3856_ hold81/A hold24/A hold44/A hold62/A VGND VPWR _3856_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_177_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6575_ _7140_/CLK _6575_/D VGND VPWR _6575_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3787_ _7159_/Q _6404_/Q _6755_/Q VGND VPWR _3788_/A VGND VPWR sky130_fd_sc_hd__nor3_1
X_5526_ hold371/X _5526_/A1 _5531_/S VGND VPWR _5526_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5457_ hold343/X _5526_/A1 _5462_/S VGND VPWR _5457_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4408_ _4633_/B _4408_/B VGND VPWR _4459_/B VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_132_156 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5388_ hold712/X _5469_/A1 _5390_/S VGND VPWR _5388_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7127_ _7130_/CLK _7127_/D fanout486/X VGND VPWR _7127_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4339_ _4739_/A _4642_/A VGND VPWR _4661_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7058_ _7058_/CLK _7058_/D _6396_/A VGND VPWR _7058_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_115_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6009_ _6939_/Q _5961_/X _6006_/X _6008_/X VGND VPWR _6014_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_27_310 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_696 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_708 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_451 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_150 _5534_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_161 hold666/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_172 _5948_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_183 _6558_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_194 _5473_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3710_ _6923_/Q _5364_/A _4044_/A _6481_/Q VGND VPWR _3710_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_81_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_716 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4690_ _4690_/A _4690_/B VGND VPWR _4690_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_119_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3641_ _3640_/Y _6729_/Q _3829_/A VGND VPWR _3641_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_146_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6360_ _6360_/A _6400_/B VGND VPWR _6360_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3572_ _6950_/Q _3781_/A2 _4145_/A _6559_/Q _3570_/X VGND VPWR _3580_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5311_ _5311_/A0 _5473_/A1 _5318_/S VGND VPWR _5311_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6291_ _6654_/Q _5973_/A _5948_/X _6699_/Q _6290_/X VGND VPWR _6291_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_605 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5242_ _5242_/A0 _5545_/A1 _5246_/S VGND VPWR _5242_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7082_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5173_ _3320_/X _3355_/X _5173_/B1 VGND VPWR _5173_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_69_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4124_ hold742/X _5469_/A1 _4126_/S VGND VPWR _4124_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput1 debug_mode VGND VPWR input1/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4055_ hold339/X _4054_/X _4067_/S VGND VPWR _4055_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk clkbuf_opt_4_0_csclk/X VGND VPWR _6908_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_37_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4957_ _4574_/Y _4956_/Y _4575_/Y VGND VPWR _4957_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3908_ _3909_/B VGND VPWR _3908_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_138_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4888_ _4469_/A _4947_/C _4887_/A _4633_/B _4379_/B VGND VPWR _4892_/B VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
X_3839_ _6488_/Q _3867_/A VGND VPWR _3860_/B VGND VPWR sky130_fd_sc_hd__nand2_2
X_6627_ _6629_/CLK _6627_/D _6390_/A VGND VPWR _6627_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_192_343 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6558_ _6712_/CLK _6558_/D _6390_/A VGND VPWR _6558_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_118_462 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5509_ hold598/X _5509_/A1 _5513_/S VGND VPWR _5509_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6489_ _3927_/A1 _6489_/D _6378_/X VGND VPWR _6489_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_106_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xwire443 _3268_/Y VGND VPWR _6367_/B VGND VPWR sky130_fd_sc_hd__buf_4
XFILLER_124_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5860_ _6461_/Q _5624_/X _5664_/X _6666_/Q VGND VPWR _5860_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_463 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4811_ _4581_/B _4947_/C _4500_/A VGND VPWR _5039_/C VGND VPWR sky130_fd_sc_hd__a21o_1
X_5791_ _6976_/Q _5634_/X _5652_/B _5790_/Y VGND VPWR _5791_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4742_ _4472_/A _4574_/B _4737_/A VGND VPWR _4996_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_193_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A _4673_/B VGND VPWR _4673_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_119_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6412_ _3568_/A1 _6412_/D _6368_/X VGND VPWR _6412_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3624_ _6933_/Q _5373_/A _4316_/A _6708_/Q VGND VPWR _3624_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_174_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6343_ _6342_/X _6343_/A1 _6346_/S VGND VPWR _7147_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_127_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3555_ _3555_/A hold66/X VGND VPWR _4238_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6274_ _6693_/Q _5954_/X _5976_/D _6622_/Q _6255_/X VGND VPWR _6275_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3486_ _3486_/A _3486_/B VGND VPWR _3486_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_102_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5225_ _5225_/A0 hold60/X _5228_/S VGND VPWR _5225_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5156_ hold832/X _6354_/A1 _5160_/S VGND VPWR _5156_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_57_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4107_ hold433/X _5528_/A1 _4108_/S VGND VPWR _4107_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5087_ _5087_/A _5087_/B _5115_/C _5087_/D VGND VPWR _5087_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_110_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_555 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4038_ _4038_/A _6352_/B VGND VPWR _4043_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_71_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_452 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A _5989_/B _5989_/C VGND VPWR _6001_/C VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_8_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _5654_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_61 _6025_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_72 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_138_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 _6949_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_94 _6837_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_180_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput190 _3200_/Y VGND VPWR mgmt_gpio_oeb[23] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_121_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_688 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_67 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold309 _6622_/Q VGND VPWR hold309/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_109_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/A VGND VPWR _7137_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_3340_ _3370_/A _3455_/A VGND VPWR _5523_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3271_ hold24/X hold44/A _6488_/Q VGND VPWR hold25/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5010_ _5010_/A _5010_/B VGND VPWR _5010_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_87_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1009 _6651_/Q VGND VPWR _4252_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7103__490 VGND VGND VPWR VPWR _7103_/D _7103__490/LO sky130_fd_sc_hd__conb_1
XFILLER_93_352 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6961_ _7017_/CLK _6961_/D fanout461/X VGND VPWR _6961_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_53_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5912_ _6474_/Q _5627_/X _5635_/X _6569_/Q VGND VPWR _5912_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6892_ _7067_/CLK _6892_/D fanout477/X VGND VPWR _6892_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5843_ _5843_/A1 _6279_/S _5842_/X VGND VPWR _7114_/D VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_21_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_468 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5774_ _6839_/Q _5657_/X _5660_/X _6807_/Q _5773_/X VGND VPWR _5774_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4725_ _5114_/A _4725_/B VGND VPWR _4725_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_30_680 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4656_ _4632_/Y _4645_/Y _4654_/X _4655_/X VGND VPWR _4660_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_174_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput70 mgmt_gpio_in[7] VGND VPWR _3959_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_3607_ _6853_/Q _5283_/A _5256_/A _6829_/Q _3590_/X VGND VPWR _3611_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xinput81 spi_sdo VGND VPWR input81/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold810 _6566_/Q VGND VPWR hold810/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold821 _4225_/X VGND VPWR _6623_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _4690_/A _4495_/A _4570_/Y _4580_/X _4586_/X VGND VPWR _4589_/D VGND VPWR
+ sky130_fd_sc_hd__o311a_1
Xinput92 spimemio_flash_io3_oeb VGND VPWR input92/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold832 _6743_/Q VGND VPWR hold832/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 _4237_/X VGND VPWR _6629_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 _6812_/Q VGND VPWR hold854/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ _6642_/Q _6326_/A2 _6326_/B1 _6643_/Q VGND VPWR _6326_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3538_ _3538_/A _3538_/B _3538_/C _3538_/D VGND VPWR _3538_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
Xhold865 _5376_/X VGND VPWR _6932_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _6471_/Q VGND VPWR hold876/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_424 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold887 _4002_/X VGND VPWR _6444_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _7077_/Q VGND VPWR hold898/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6257_ _7154_/Q _5958_/X _5978_/X _6483_/Q VGND VPWR _6257_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3469_ _3956_/A _4083_/S _5337_/A _6903_/Q _3468_/X VGND VPWR _3472_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5208_ hold168/X hold42/X _5210_/S VGND VPWR _5208_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6188_ _6665_/Q _5938_/X _5952_/X _6705_/Q _6187_/X VGND VPWR _6189_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1510 hold20/A VGND VPWR _3254_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_691 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1521 _5757_/X VGND VPWR _7110_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1532 _7160_/Q VGND VPWR _3260_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5139_ _5001_/B _5077_/C _5138_/X _5103_/Y VGND VPWR _5143_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_123_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1543 _7169_/Q VGND VPWR _3248_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _6720_/Q VGND VPWR _4731_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 hold44/A VGND VPWR _3866_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1576 _6524_/Q VGND VPWR hold1576/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1587 _6525_/Q VGND VPWR hold622/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 _7185_/A VGND VPWR hold1598/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_590 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_51 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4510_ _4902_/A _4456_/Y _4509_/X VGND VPWR _4510_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_117_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5490_ _5490_/A _5490_/B VGND VPWR _5495_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_117_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold106 _7147_/Q VGND VPWR hold106/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _4441_/A _4441_/B VGND VPWR _4947_/B VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold117 _5387_/X VGND VPWR _6942_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _5225_/X VGND VPWR _6798_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold139 _6792_/Q VGND VPWR hold139/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_7160_ net399_2/A _7160_/D _6390_/X VGND VPWR _7160_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4372_ _4702_/B _4591_/A VGND VPWR _4372_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_6111_ _6895_/Q _5946_/X _5955_/X _6807_/Q VGND VPWR _6111_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_98_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3323_ hold34/X _3323_/B hold72/X VGND VPWR hold73/A VGND VPWR sky130_fd_sc_hd__and3_4
X_7091_ _7113_/CLK _7091_/D fanout460/X VGND VPWR _7091_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_112_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6042_ _6908_/Q _5973_/A _5948_/X _6948_/Q _6041_/X VGND VPWR _6042_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3254_ hold97/A _3254_/A1 _3260_/S VGND VPWR _3254_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3185_ _6657_/Q VGND VPWR _3185_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_54_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6944_ _6981_/CLK _6944_/D fanout463/X VGND VPWR _6944_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6875_ _7067_/CLK _6875_/D fanout477/X VGND VPWR _6875_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_179_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5826_ _6465_/Q _5619_/X _5663_/X _6609_/Q VGND VPWR _5826_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_22_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5757_ _5757_/A0 _5756_/X _6279_/S VGND VPWR _5757_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_148_674 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4708_ _4469_/A _4689_/B _4639_/Y _4690_/Y VGND VPWR _5062_/B VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_175_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5688_ _6987_/Q _5627_/X _5661_/X _6875_/Q VGND VPWR _5688_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4639_ _4716_/A _4707_/C VGND VPWR _4639_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold640 _6422_/Q VGND VPWR hold640/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold651 _5513_/X VGND VPWR _7054_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap370 hold36/X VGND VPWR _3814_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold662 _6616_/Q VGND VPWR hold662/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 _6912_/Q VGND VPWR hold673/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold684 _5217_/X VGND VPWR _6791_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6309_ _3762_/Y _6309_/A1 _6315_/S VGND VPWR _7134_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold695 _5379_/X VGND VPWR _6935_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_254 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1340 hold1340/A VGND VPWR wb_dat_o[15] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1351 _4164_/A1 VGND VPWR hold1351/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 hold1362/A VGND VPWR wb_dat_o[29] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1373 _6308_/A1 VGND VPWR hold1373/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_175_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1384 _7175_/A VGND VPWR _4076_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1395 _7025_/Q VGND VPWR _5480_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_138 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4990_ _4948_/A _4428_/Y _4846_/B _4645_/Y VGND VPWR _5003_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_63_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3941_ _3975_/S _3941_/B VGND VPWR _3941_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
X_6660_ _7058_/CLK _6660_/D _6396_/A VGND VPWR _6660_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3872_ _7170_/Q _6402_/Q _3867_/A VGND VPWR _3872_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_149_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5611_ _5552_/B _5606_/A _5610_/Y VGND VPWR _5611_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_6591_ _7130_/CLK _6591_/D VGND VPWR _6591_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_192_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5542_ _5542_/A0 hold667/X _5549_/S VGND VPWR _5542_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_157_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5473_ _5473_/A0 _5473_/A1 hold30/X VGND VPWR _5473_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4424_ _4500_/A _4581_/B VGND VPWR _4424_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_160_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7143_ _7150_/CLK _7143_/D fanout487/X VGND VPWR hold4/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4355_ _4556_/A _4563_/A _4753_/A _4607_/A _4642_/A VGND VPWR _4356_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_113_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout405 hold59/X VGND VPWR _5519_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout416 _5465_/A1 VGND VPWR _6354_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout427 _5490_/B VGND VPWR _6352_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_3306_ _3554_/A _3379_/A VGND VPWR _5346_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_140_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xfanout438 _6507_/Q VGND VPWR _5552_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_7074_ _7085_/CLK _7074_/D fanout479/X VGND VPWR _7074_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout449 fanout450/X VGND VPWR fanout449/X VGND VPWR sky130_fd_sc_hd__buf_6
X_4286_ _4286_/A _4322_/B VGND VPWR _4291_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_6025_ _6017_/X _6025_/B _6226_/B VGND VPWR _6025_/X VGND VPWR sky130_fd_sc_hd__and3b_2
X_3237_ _6417_/Q _6416_/Q VGND VPWR _3239_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_100_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3168_ _3168_/A VGND VPWR _3910_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_54_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_388 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6927_ _7054_/CLK _6927_/D fanout460/X VGND VPWR _6927_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6858_ _6926_/CLK _6858_/D fanout457/X VGND VPWR _6858_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_168_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5809_ _6985_/Q _5624_/X _5634_/X _6977_/Q _5802_/Y VGND VPWR _5809_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6789_ _6963_/CLK _6789_/D fanout456/X VGND VPWR _6789_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_129_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_688 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold470 _5415_/X VGND VPWR _6967_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold481 _6673_/Q VGND VPWR hold481/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _4248_/X VGND VPWR _6648_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1170 _4070_/X VGND VPWR _6498_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_642 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1181 _6764_/Q VGND VPWR _5185_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _5365_/X VGND VPWR _6922_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_163 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_460 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4140_ _4140_/A0 _6353_/A1 _4144_/S VGND VPWR _4140_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_609 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4071_ hold824/X _6354_/A1 _4118_/B VGND VPWR _4071_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4973_ _4616_/Y _4628_/Y _4970_/Y VGND VPWR _4974_/D VGND VPWR sky130_fd_sc_hd__a21o_1
X_6712_ _6712_/CLK _6712_/D fanout470/X VGND VPWR _6712_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3924_ _6519_/Q input78/X _3957_/B VGND VPWR _3924_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_189_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6643_ _7150_/CLK _6643_/D fanout487/X VGND VPWR _6643_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3855_ _3854_/X _3855_/A1 _3866_/S VGND VPWR _6411_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_6574_ _7137_/CLK _6574_/D VGND VPWR _6574_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3786_ _6866_/Q _5301_/A _4038_/A _6475_/Q _3785_/X VGND VPWR _3793_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5525_ hold543/X _5543_/A1 _5531_/S VGND VPWR _5525_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5456_ hold253/X _5465_/A1 _5462_/S VGND VPWR _5456_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4407_ _4551_/A _4570_/A VGND VPWR _4498_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_5387_ hold116/X hold60/X _5390_/S VGND VPWR _5387_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_132_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7126_ _7126_/CLK _7126_/D fanout459/X VGND VPWR _7126_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4338_ _4338_/A _4338_/B _4338_/C VGND VPWR _4564_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_115_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7057_ _7079_/CLK _7057_/D fanout478/X VGND VPWR _7057_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4269_ _4269_/A0 _6353_/A1 _4273_/S VGND VPWR _4269_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6008_ _7011_/Q _5940_/X _5967_/X _6851_/Q _6005_/X VGND VPWR _6008_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_322 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_566 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_712 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_140 _6226_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_151 _5473_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_162 _5193_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_173 _5953_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_184 _6853_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_195 _5490_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3640_ _3597_/X _3640_/B _3640_/C _3640_/D VGND VPWR _3640_/Y VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_127_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3571_ _3571_/A _3571_/B VGND VPWR _4145_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_155_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5310_ _5310_/A _5541_/B VGND VPWR _5318_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6290_ _6649_/Q _5976_/C _5971_/D _6569_/Q VGND VPWR _6290_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5241_ hold854/X _5484_/A1 _5246_/S VGND VPWR _5241_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5172_ _5172_/A0 _5491_/A1 _5172_/S VGND VPWR _5172_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4123_ hold158/X hold60/X _4126_/S VGND VPWR _4123_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_575 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput2 debug_oeb VGND VPWR input2/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4054_ hold622/X _5534_/A1 _4058_/S VGND VPWR _4054_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_opt_1_0_csclk clkbuf_3_1_0_csclk/X VGND VPWR clkbuf_leaf_4_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4956_ _4965_/B _5051_/A _4554_/B VGND VPWR _4956_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3907_ _3907_/A _3907_/B _3907_/C _3907_/D VGND VPWR _3909_/B VGND VPWR sky130_fd_sc_hd__nand4_2
X_4887_ _4887_/A _4887_/B VGND VPWR _4900_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_6626_ _6769_/CLK _6626_/D fanout469/X VGND VPWR _6626_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3838_ _3838_/A _3838_/B VGND VPWR _6415_/D VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_192_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6557_ _6629_/CLK _6557_/D _6390_/A VGND VPWR _6557_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3769_ _6786_/Q _5211_/A _4280_/A _6675_/Q VGND VPWR _3769_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_3_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5508_ hold335/X _5526_/A1 _5513_/S VGND VPWR _5508_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6488_ _3927_/A1 _6488_/D _6377_/X VGND VPWR _6488_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5439_ hold337/X _5526_/A1 _5444_/S VGND VPWR _5439_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7109_ _7126_/CLK _7109_/D fanout456/X VGND VPWR _7109_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_47_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_214 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_741 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4810_ _4810_/A _4810_/B VGND VPWR _4810_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_92_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5790_ _6920_/Q _5899_/B VGND VPWR _5790_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_33_199 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4741_ _4741_/A _4741_/B VGND VPWR _4992_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_4672_ _4672_/A _4672_/B VGND VPWR _4984_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_6411_ _3568_/A1 _6411_/D _6367_/X VGND VPWR hold70/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3623_ _7021_/Q hold29/A _4127_/A _6543_/Q _3587_/X VGND VPWR _3628_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6342_ _6642_/Q _6342_/A2 _6342_/B1 _6350_/A2 _6341_/X VGND VPWR _6342_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3554_ _3554_/A _3814_/B VGND VPWR _4268_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_6273_ _6558_/Q _5971_/B _5949_/X _6678_/Q _6272_/X VGND VPWR _6275_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_3485_ _3485_/A _3485_/B _3485_/C VGND VPWR _3486_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_103_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5224_ hold200/X _5494_/A1 _5228_/S VGND VPWR _5224_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5155_ _5155_/A0 _5491_/A1 _5160_/S VGND VPWR _5155_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4106_ hold752/X _6356_/A1 _4108_/S VGND VPWR _4106_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5086_ _5088_/A _5086_/B _5086_/C VGND VPWR _5114_/D VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_56_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_567 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4037_ hold582/X _6357_/A1 _4037_/S VGND VPWR _4037_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5988_ _7047_/Q _5971_/A _5938_/X _6922_/Q _5980_/X VGND VPWR _5989_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4939_ _4460_/A _4484_/Y _4967_/A _4563_/A _4923_/Y VGND VPWR _5073_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_40 _5300_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_51 _5940_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_62 _6025_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA_73 _6100_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_138_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6609_ _6653_/CLK _6609_/D fanout454/X VGND VPWR _6609_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA_84 _7152_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_33 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_95 _6405_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_137_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_306 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput180 _3209_/Y VGND VPWR mgmt_gpio_oeb[14] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput191 _3199_/Y VGND VPWR mgmt_gpio_oeb[24] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_94_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_44_csclk _6888_/CLK VGND VPWR _7016_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_109_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_369 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_274 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3270_ _7171_/Q hold15/A _6487_/Q _3875_/B VGND VPWR _7156_/D VGND VPWR sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_59_csclk _6447_/CLK VGND VPWR _7053_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_112_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6960_ _6997_/CLK _6960_/D fanout465/X VGND VPWR _6960_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_19_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5911_ _3225_/Y _5899_/B _5651_/B VGND VPWR _5911_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_6891_ _7067_/CLK _6891_/D fanout477/X VGND VPWR _6891_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5842_ _5552_/B _7113_/Q _6103_/B1 _5841_/X VGND VPWR _5842_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_22_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5773_ hold56/A _5619_/X _5663_/X _6863_/Q VGND VPWR _5773_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4724_ _4724_/A _4972_/A VGND VPWR _4775_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_147_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4655_ _4626_/Y _4628_/Y _4653_/Y _4609_/Y VGND VPWR _4655_/X VGND VPWR sky130_fd_sc_hd__o22a_1
Xinput60 mgmt_gpio_in[31] VGND VPWR input60/X VGND VPWR sky130_fd_sc_hd__buf_2
Xhold800 _6823_/Q VGND VPWR hold800/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3606_ _6797_/Q _3326_/Y _4139_/A _6553_/Q _3605_/X VGND VPWR _3611_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xinput71 mgmt_gpio_in[8] VGND VPWR input71/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold811 _4159_/X VGND VPWR _6566_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput82 spi_sdoenb VGND VPWR input82/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4563_/A _4951_/B _4942_/A _4583_/X VGND VPWR _4586_/X VGND VPWR sky130_fd_sc_hd__o211a_1
Xinput93 trap VGND VPWR input93/X VGND VPWR sky130_fd_sc_hd__buf_4
Xhold822 _6605_/Q VGND VPWR hold822/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _5156_/X VGND VPWR _6743_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _6828_/Q VGND VPWR hold844/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _6324_/X _6325_/A1 _6346_/S VGND VPWR _7141_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold855 _5241_/X VGND VPWR _6812_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3537_ _6926_/Q _5364_/A _3964_/A _6422_/Q _3536_/X VGND VPWR _3538_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold866 _6547_/Q VGND VPWR hold866/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _4034_/X VGND VPWR _6471_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _6652_/Q VGND VPWR hold888/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold899 _5539_/X VGND VPWR _7077_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _6612_/Q _5943_/X _5981_/X _6658_/Q VGND VPWR _6256_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_170_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3468_ _7076_/Q _5532_/A _5319_/A _6887_/Q VGND VPWR _3468_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_76_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5207_ hold766/X _5528_/A1 _5210_/S VGND VPWR _5207_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6187_ _6460_/Q _5945_/X _5975_/C _6578_/Q VGND VPWR _6187_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_191_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1500 hold4/A VGND VPWR _6331_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3399_ _6841_/Q _5265_/A hold76/A _7046_/Q _3398_/X VGND VPWR _3409_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1511 _3254_/X VGND VPWR _7166_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1522 hold11/A VGND VPWR _6328_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1533 _7148_/Q VGND VPWR _6346_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5138_ _5138_/A _5138_/B _5138_/C VGND VPWR _5138_/X VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1544 _3248_/X VGND VPWR _7169_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1555 hold62/A VGND VPWR _3858_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 _6637_/Q VGND VPWR _3879_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 _6755_/Q VGND VPWR hold1577/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1588 _7177_/A VGND VPWR hold405/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5069_ _5069_/A _5069_/B _5069_/C _5069_/D VGND VPWR _5103_/B VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1599 _7089_/Q VGND VPWR _5561_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_764 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_770 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4440_ _4690_/A _4495_/A VGND VPWR _4724_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_172_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold107 _3977_/X VGND VPWR hold98/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_133 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold118 _6790_/Q VGND VPWR hold118/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A VGND VPWR hold129/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4371_ _4702_/A _4566_/A VGND VPWR _4374_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_98_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6110_ _6943_/Q _5961_/X _6108_/X _6109_/X VGND VPWR _6115_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3322_ _3455_/A hold48/X VGND VPWR _5193_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_152_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7090_ _7113_/CLK _7090_/D fanout460/X VGND VPWR _7090_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_58_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6041_ _6900_/Q _5976_/C _5971_/D _6828_/Q VGND VPWR _6041_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3253_ _3252_/Y _3253_/A1 _3253_/S VGND VPWR _7167_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3184_ _6541_/Q VGND VPWR _3184_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6943_ _6999_/CLK _6943_/D fanout464/X VGND VPWR _6943_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_19_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6874_ _7051_/CLK _6874_/D fanout476/X VGND VPWR _6874_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_5825_ _6695_/Q _5637_/X _5645_/X _6455_/Q VGND VPWR _5825_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_179_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5756_ _7109_/Q _5755_/X _6303_/S VGND VPWR _5756_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4707_ _4716_/A _4911_/B _4707_/C VGND VPWR _4707_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
X_5687_ _7011_/Q _5630_/X _5635_/X _6827_/Q _5686_/X VGND VPWR _5690_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4638_ _4638_/A _4661_/B VGND VPWR _4638_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
Xhold630 _6431_/Q VGND VPWR hold630/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold641 _3974_/X VGND VPWR _6422_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _4636_/A _5043_/A _4737_/A VGND VPWR _5099_/A VGND VPWR sky130_fd_sc_hd__nand3_2
Xhold652 _6829_/Q VGND VPWR hold652/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmax_cap371 hold35/X VGND VPWR hold36/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold663 _4217_/X VGND VPWR _6616_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap382 _5660_/X VGND VPWR _5913_/B1 VGND VPWR sky130_fd_sc_hd__buf_6
Xhold674 _5353_/X VGND VPWR _6912_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ _3828_/Y _6308_/A1 _6315_/S VGND VPWR _7133_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold685 _6993_/Q VGND VPWR hold685/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/A VGND VPWR hold696/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6239_ _6462_/Q _5945_/X _5975_/C _6580_/Q _6238_/X VGND VPWR _6240_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1330 hold1330/A VGND VPWR wb_dat_o[8] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1341 hold1426/X VGND VPWR hold1341/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1352 hold1352/A VGND VPWR wb_dat_o[16] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_85_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1363 _6309_/A1 VGND VPWR hold1363/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1374 hold1374/A VGND VPWR wb_dat_o[24] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1385 _6529_/Q VGND VPWR _4115_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 _7161_/Q VGND VPWR hold1/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_75 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3940_ _7105_/Q _6758_/Q _6762_/Q VGND VPWR _3940_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3871_ _3837_/B _3912_/B1 _3837_/C _6403_/Q VGND VPWR _6403_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_5610_ _6507_/Q _5610_/B VGND VPWR _5610_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_83_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6590_ _7137_/CLK _6590_/D VGND VPWR _6590_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_5541_ _5541_/A _5541_/B VGND VPWR _5549_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_157_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5472_ hold29/X _5541_/B VGND VPWR hold30/A VGND VPWR sky130_fd_sc_hd__and2_4
X_4423_ _4600_/B _4626_/B VGND VPWR _4581_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_160_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7142_ _3937_/A1 _7142_/D fanout487/X VGND VPWR hold11/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4354_ _4642_/A _4357_/B VGND VPWR _4356_/A VGND VPWR sky130_fd_sc_hd__nor2_1
Xfanout406 _5494_/A1 VGND VPWR _6356_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_113_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout417 _5465_/A1 VGND VPWR _5492_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
Xfanout428 hold17/X VGND VPWR _5490_/B VGND VPWR sky130_fd_sc_hd__buf_4
X_3305_ _3313_/A hold27/X VGND VPWR _3379_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7073_ _7083_/CLK _7073_/D _6390_/A VGND VPWR _7073_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4285_ hold229/X hold60/X _4285_/S VGND VPWR _4285_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6024_ _6024_/A _6024_/B _6024_/C _6024_/D VGND VPWR _6025_/B VGND VPWR sky130_fd_sc_hd__nor4_1
X_3236_ _6417_/Q _6416_/Q VGND VPWR _3264_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_73_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3167_ hold44/A VGND VPWR _3167_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_27_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6926_ _6926_/CLK _6926_/D fanout457/X VGND VPWR _6926_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_6857_ _7086_/CLK _6857_/D fanout482/X VGND VPWR _6857_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_167_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5808_ _6945_/Q _5632_/X _5804_/X _5805_/X _5807_/X VGND VPWR _5808_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6788_ _7012_/CLK hold19/X fanout458/X VGND VPWR _6788_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_148_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5739_ _7022_/Q _5619_/X _5663_/X _6862_/Q VGND VPWR _5739_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_129_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold460 _5288_/X VGND VPWR _6854_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_391 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold471 _6662_/Q VGND VPWR hold471/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _4278_/X VGND VPWR _6673_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold493 _6612_/Q VGND VPWR hold493/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _5194_/X VGND VPWR _6770_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _6810_/Q VGND VPWR _5239_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _5185_/X VGND VPWR _6764_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1193 _6700_/Q VGND VPWR _4311_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_472 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR _3568_/A1 VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_5_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4070_ _4070_/A0 _4069_/X _4084_/S VGND VPWR _4070_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4972_ _4972_/A _5010_/B VGND VPWR _5008_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_51_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6711_ _6714_/CLK _6711_/D fanout470/X VGND VPWR _6711_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3923_ _6518_/Q input80/X _3957_/B VGND VPWR _3923_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_189_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6642_ _7150_/CLK _6642_/D fanout487/X VGND VPWR _6642_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3854_ _3284_/X _3283_/Y _3854_/S VGND VPWR _3854_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6573_ _7140_/CLK _6573_/D VGND VPWR _6573_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3785_ _7039_/Q hold76/A _4322_/A _6710_/Q VGND VPWR _3785_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_164_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5524_ _5524_/A0 _5524_/A1 _5531_/S VGND VPWR _5524_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5455_ _5455_/A0 _5524_/A1 _5462_/S VGND VPWR _5455_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4406_ _4739_/A _4415_/A VGND VPWR _4570_/A VGND VPWR sky130_fd_sc_hd__and2b_1
X_5386_ hold217/X _5494_/A1 _5390_/S VGND VPWR _5386_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7125_ _7126_/CLK _7125_/D fanout459/X VGND VPWR _7125_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4337_ _4337_/A _4337_/B _4337_/C _4337_/D VGND VPWR _4338_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_59_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7056_ _7085_/CLK _7056_/D fanout485/X VGND VPWR _7056_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4268_ _4268_/A _5490_/B VGND VPWR _4273_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_6007_ _7080_/Q _5976_/B _5954_/X _7056_/Q _6004_/X VGND VPWR _6024_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3219_ _6821_/Q VGND VPWR _3219_/Y VGND VPWR sky130_fd_sc_hd__clkinv_2
X_4199_ _4199_/A0 _5544_/A1 _4201_/S VGND VPWR _4199_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6909_ _7076_/CLK _6909_/D fanout481/X VGND VPWR _6909_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_24_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_381 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold290 _5222_/X VGND VPWR _6795_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_130 _3923_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_141 _6226_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 _5552_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_163 _5532_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_174 _5976_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_185 _7173_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_196 hold94/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3570_ _7059_/Q hold86/A _4008_/A _6454_/Q VGND VPWR _3570_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5240_ hold604/X _5543_/A1 _5246_/S VGND VPWR _5240_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_510 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5171_ _5186_/A _5171_/B _6352_/B VGND VPWR _5172_/S VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_68_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4122_ hold243/X _5494_/A1 _4126_/S VGND VPWR _4122_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4053_ _4053_/A0 _4052_/X _4067_/S VGND VPWR _4053_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput3 debug_out VGND VPWR input3/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4955_ _5068_/A _4964_/B _5068_/B VGND VPWR _5039_/D VGND VPWR sky130_fd_sc_hd__and3_1
X_3906_ _3906_/A _3906_/B _3906_/C VGND VPWR _3907_/D VGND VPWR sky130_fd_sc_hd__and3_1
X_4886_ _5010_/A _4886_/B VGND VPWR _4887_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_177_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6625_ _6629_/CLK _6625_/D _6390_/A VGND VPWR _6625_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3837_ _3837_/A _3837_/B _3837_/C VGND VPWR _3838_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_6556_ _6629_/CLK _6556_/D _6390_/A VGND VPWR _6556_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3768_ _6418_/Q _3964_/A _4014_/A _6455_/Q _3767_/X VGND VPWR _3773_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5507_ hold558/X _5543_/A1 _5513_/S VGND VPWR _5507_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6487_ _3945_/A1 _6487_/D _6376_/X VGND VPWR _6487_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3699_ _3699_/A _3699_/B _3699_/C _3699_/D VGND VPWR _3700_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_5438_ hold570/X _5543_/A1 _5444_/S VGND VPWR _5438_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput340 hold1375/X VGND VPWR hold1376/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5369_ hold568/X _6357_/A1 _5372_/S VGND VPWR _5369_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7108_ _7126_/CLK _7108_/D fanout456/X VGND VPWR _7108_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_47_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7039_ _7083_/CLK _7039_/D fanout470/X VGND VPWR _7039_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_75_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_226 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_353 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_547 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_407 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4740_ _4740_/A _4740_/B VGND VPWR _4741_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_187_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_364 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4671_ _4671_/A VGND VPWR _4679_/B VGND VPWR sky130_fd_sc_hd__clkinv_2
X_6410_ _3568_/A1 _6410_/D _6366_/X VGND VPWR hold62/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3622_ _6429_/Q _3981_/A _4304_/A _6698_/Q _3621_/X VGND VPWR _3628_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6341_ _6644_/Q _6341_/A2 _6341_/B1 _6643_/Q VGND VPWR _6341_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3553_ hold36/X _3562_/B VGND VPWR _4298_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_6272_ _7037_/Q _5601_/X _5959_/X _6718_/Q VGND VPWR _6272_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3484_ _3484_/A _3484_/B _3484_/C _3484_/D VGND VPWR _3485_/C VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_142_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5223_ hold381/X _5526_/A1 _5228_/S VGND VPWR _5223_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5154_ _5154_/A _6352_/B VGND VPWR _5160_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_111_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4105_ hold237/X _5544_/A1 _4108_/S VGND VPWR _4105_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5085_ _5085_/A _5085_/B _5085_/C VGND VPWR _5087_/D VGND VPWR sky130_fd_sc_hd__and3_1
X_4036_ hold778/X _6356_/A1 _4037_/S VGND VPWR _4036_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_646 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5987_ _6442_/Q _5601_/X _5981_/X _6914_/Q _5950_/X VGND VPWR _5989_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XPHY_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4938_ _5068_/A _5046_/A _5068_/B _5103_/A VGND VPWR _4941_/B VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_30 _3612_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_41 _5300_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4869_ _4841_/X _4869_/B _4869_/C _4869_/D VGND VPWR _4870_/C VGND VPWR sky130_fd_sc_hd__and4b_1
XANTENNA_52 _5973_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_63 _6025_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_74 _6268_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6608_ _6746_/CLK _6608_/D fanout448/X VGND VPWR _6608_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XANTENNA_85 _6467_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_96 _6406_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_21_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6539_ _6539_/CLK _6539_/D fanout461/X VGND VPWR _6539_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_137_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_318 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput181 _3208_/Y VGND VPWR mgmt_gpio_oeb[15] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput192 _3198_/Y VGND VPWR mgmt_gpio_oeb[25] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_47_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_259 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_624 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1177_ clkbuf_0__1177_/X VGND VPWR _6312_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_171_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5910_ _6618_/Q _5628_/X _5910_/B1 _6629_/Q VGND VPWR _5910_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6890_ _6890_/CLK _6890_/D fanout476/X VGND VPWR _6890_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_34_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5841_ _6540_/Q _5652_/Y _5828_/X _5840_/X _6303_/S VGND VPWR _5841_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5772_ _6903_/Q _5621_/X _5648_/X _6855_/Q _5771_/X VGND VPWR _5772_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4723_ _4984_/A _4723_/B VGND VPWR _5046_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_4654_ _4619_/Y _4653_/Y _4846_/B VGND VPWR _4654_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_147_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput50 mgmt_gpio_in[22] VGND VPWR input50/X VGND VPWR sky130_fd_sc_hd__buf_2
X_3605_ _6628_/Q _4232_/A _4244_/A _6648_/Q VGND VPWR _3605_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xinput61 mgmt_gpio_in[32] VGND VPWR input61/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput72 mgmt_gpio_in[9] VGND VPWR input72/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold801 _5253_/X VGND VPWR _6823_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4585_ _5051_/A _4881_/B VGND VPWR _4951_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_174_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold812 hold812/A VGND VPWR hold812/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VPWR input83/X VGND VPWR sky130_fd_sc_hd__buf_2
Xhold823 _4204_/X VGND VPWR _6605_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput94 uart_enabled VGND VPWR _3956_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xhold834 _6701_/Q VGND VPWR hold834/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ _6644_/Q _6324_/A2 _6324_/B1 _6643_/Q _6323_/X VGND VPWR _6324_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3536_ _7075_/Q _5532_/A _4286_/A _6684_/Q VGND VPWR _3536_/X VGND VPWR sky130_fd_sc_hd__a22o_2
Xhold845 _5259_/X VGND VPWR _6828_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _6908_/Q VGND VPWR hold856/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold867 _4136_/X VGND VPWR _6547_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _7028_/Q VGND VPWR hold878/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _4253_/X VGND VPWR _6652_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _6663_/Q _5976_/B _5971_/C _6713_/Q VGND VPWR _6255_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3467_ _3467_/A _3467_/B _3467_/C _3467_/D VGND VPWR _3467_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_5206_ hold904/X _5509_/A1 _5210_/S VGND VPWR _5206_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6186_ _6450_/Q _5947_/X _5965_/X _6545_/Q _6185_/X VGND VPWR _6189_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3398_ input28/X _3367_/Y _3964_/A _6425_/Q _3384_/X VGND VPWR _3398_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1501 _7120_/Q VGND VPWR _6028_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _6598_/Q VGND VPWR _4195_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _4428_/Y _4542_/D _4846_/B _4653_/Y _4769_/A VGND VPWR _5138_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold1523 _7144_/Q VGND VPWR _6334_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1534 _7123_/Q VGND VPWR _6104_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1545 _7183_/A VGND VPWR hold89/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 _6506_/Q VGND VPWR _3894_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1567 _6417_/Q VGND VPWR _3834_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _5068_/A _5068_/B _5068_/C VGND VPWR _5069_/D VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1578 _6538_/Q VGND VPWR hold1578/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1589 _6532_/Q VGND VPWR hold1589/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4019_ hold616/X _6357_/A1 _4019_/S VGND VPWR _4019_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_443 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold108 hold98/X VGND VPWR hold108/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold119 _5216_/X VGND VPWR _6790_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_145 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4370_ _4556_/A _4441_/A VGND VPWR _4495_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_125_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3321_ hold47/X _3454_/B VGND VPWR hold48/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_98_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6040_ _6040_/A _6040_/B _6040_/C VGND VPWR _6040_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_3252_ _7167_/Q _6485_/Q _3262_/C VGND VPWR _3252_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_79_660 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3183_ _6655_/Q VGND VPWR _3183_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_94_652 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_302 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6942_ _7006_/CLK _6942_/D fanout457/X VGND VPWR _6942_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6873_ _7070_/CLK _6873_/D fanout473/X VGND VPWR _6873_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_744 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5824_ _6599_/Q _5616_/X _5655_/X _6545_/Q _5823_/X VGND VPWR _5824_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5755_ wire367/X _5754_/Y _6790_/Q _5652_/Y VGND VPWR _5755_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4706_ _4693_/X _4706_/B _4706_/C _4706_/D VGND VPWR _4722_/B VGND VPWR sky130_fd_sc_hd__and4b_1
X_5686_ _6851_/Q _5648_/X _5910_/B1 _6883_/Q VGND VPWR _5686_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4637_ _4638_/A _4661_/B VGND VPWR _4707_/C VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_175_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_186 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_443 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold620 _6430_/Q VGND VPWR hold620/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _3987_/X VGND VPWR _6431_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _4664_/B _4568_/B VGND VPWR _4741_/A VGND VPWR sky130_fd_sc_hd__nand2b_2
Xhold642 _6657_/Q VGND VPWR hold642/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap361 hold37/X VGND VPWR _4058_/S VGND VPWR sky130_fd_sc_hd__buf_6
Xhold653 _5260_/X VGND VPWR _6829_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _7141_/Q VGND VPWR hold664/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6307_ _6636_/Q _6307_/B VGND VPWR _6315_/S VGND VPWR sky130_fd_sc_hd__nand2_4
X_3519_ _6910_/Q _5346_/A _4214_/A _6618_/Q _3518_/X VGND VPWR _3523_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xmax_cap383 _5658_/X VGND VPWR _5910_/B1 VGND VPWR sky130_fd_sc_hd__buf_8
Xhold675 _6913_/Q VGND VPWR hold675/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _5444_/X VGND VPWR _6993_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _5051_/B _4582_/B VGND VPWR _4535_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold697 _5179_/X VGND VPWR _6760_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6238_ _6667_/Q _5938_/X _5952_/X _6707_/Q VGND VPWR _6238_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_57_310 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6169_ _7054_/Q _5971_/A _5979_/X _6993_/Q VGND VPWR _6169_/X VGND VPWR sky130_fd_sc_hd__a22o_2
Xhold1320 hold1320/A VGND VPWR wb_dat_o[18] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_85_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1331 hold1420/X VGND VPWR hold1331/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 hold1342/A VGND VPWR wb_dat_o[9] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1353 _4183_/A1 VGND VPWR hold1353/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 hold1364/A VGND VPWR wb_dat_o[25] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_45_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1375 _4192_/A1 VGND VPWR hold1375/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 _7044_/Q VGND VPWR _5502_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1397 _7086_/Q VGND VPWR _5549_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_43_csclk _6888_/CLK VGND VPWR _6920_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_25_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_csclk _6447_/CLK VGND VPWR _6953_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_43_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_595 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_376 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3870_ _6404_/Q _3912_/A1 _3870_/S VGND VPWR _6404_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XPHY_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5540_ hold397/X _5540_/A1 _5540_/S VGND VPWR _5540_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_192_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5471_ hold626/X _5513_/A1 _5471_/S VGND VPWR _5471_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4422_ _4607_/A _4947_/A VGND VPWR _4921_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_7141_ _7150_/CLK _7141_/D fanout487/X VGND VPWR _7141_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_125_370 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4353_ _4379_/B _4360_/B VGND VPWR _4896_/A VGND VPWR sky130_fd_sc_hd__and2_1
Xfanout407 hold156/X VGND VPWR _5494_/A1 VGND VPWR sky130_fd_sc_hd__buf_12
Xfanout418 hold13/X VGND VPWR _5465_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_3304_ _3313_/A hold27/X VGND VPWR _5190_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_7072_ _7083_/CLK _7072_/D fanout470/X VGND VPWR _7072_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_98_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout429 hold16/X VGND VPWR hold17/A VGND VPWR sky130_fd_sc_hd__buf_8
X_4284_ hold194/X _5494_/A1 _4285_/S VGND VPWR _4284_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6023_ _6811_/Q _5971_/B _5949_/X _6931_/Q _6022_/X VGND VPWR _6024_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_3235_ _3235_/A0 _3251_/A _3235_/S VGND VPWR _7170_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3166_ _6415_/Q VGND VPWR _3837_/A VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_27_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6925_ _6925_/CLK _6925_/D fanout461/X VGND VPWR _6925_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_35_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6856_ _6981_/CLK _6856_/D fanout464/X VGND VPWR _6856_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5807_ _7017_/Q _5630_/X _5638_/X _6961_/Q _5806_/X VGND VPWR _5807_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6787_ _7012_/CLK _6787_/D fanout458/X VGND VPWR _6787_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3999_ _3999_/A _5541_/B VGND VPWR _4007_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_13_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5738_ _6966_/Q _5642_/X _5667_/X _6814_/Q VGND VPWR _5738_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_129_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5669_ _5669_/A _5669_/B _5669_/C _5669_/D VGND VPWR _5670_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_191_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold450 _5352_/X VGND VPWR _6911_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 _6627_/Q VGND VPWR hold461/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 _4265_/X VGND VPWR _6662_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _7051_/Q VGND VPWR hold483/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _4212_/X VGND VPWR _6612_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_600 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1150 _5347_/X VGND VPWR _6906_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1161 _7018_/Q VGND VPWR _5473_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _5239_/X VGND VPWR _6810_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 _6455_/Q VGND VPWR _4015_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 _4311_/X VGND VPWR _6700_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_338 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VPWR clkbuf_3_3_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_1_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4971_ _4691_/A _4902_/B _4625_/B _4645_/Y VGND VPWR _4974_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_91_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6710_ _6714_/CLK _6710_/D fanout470/X VGND VPWR _6710_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_51_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3922_ _3188_/Y input82/X _3957_/B VGND VPWR _3922_/X VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_189_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_535 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6641_ _7150_/CLK _6641_/D fanout487/X VGND VPWR _6641_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3853_ _3853_/A _3853_/B VGND VPWR _6412_/D VGND VPWR sky130_fd_sc_hd__xnor2_1
X_6572_ _7140_/CLK _6572_/D VGND VPWR _6572_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3784_ _6954_/Q _5400_/A _5154_/A _6742_/Q _3783_/X VGND VPWR _3793_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5523_ _5523_/A _5541_/B VGND VPWR _5531_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_157_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5454_ _5454_/A hold17/X VGND VPWR _5461_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_105_307 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4405_ _4459_/A _4549_/A VGND VPWR _4810_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_132_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5385_ hold399/X _5526_/A1 _5390_/S VGND VPWR _5385_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_703 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7124_ _7131_/CLK _7124_/D fanout459/X VGND VPWR _7124_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4336_ _4336_/A _4336_/B _4336_/C _4336_/D VGND VPWR _4338_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_113_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7055_ _7079_/CLK _7055_/D _6396_/A VGND VPWR _7055_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_59_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4267_ hold830/X _5546_/A1 _4267_/S VGND VPWR _4267_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6006_ _7003_/Q _5958_/X _5978_/X _6995_/Q VGND VPWR _6006_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3218_ _6829_/Q VGND VPWR _3218_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4198_ _4198_/A0 _5492_/A1 _4201_/S VGND VPWR _4198_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_644 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_154 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6908_ _6908_/CLK _6908_/D fanout475/X VGND VPWR _6908_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6839_ _6865_/CLK _6839_/D fanout464/X VGND VPWR _6839_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_50_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold280 _5188_/X VGND VPWR _6766_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold291/A VGND VPWR hold291/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_677 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_120 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_131 _3925_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_142 _6279_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_647 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_153 _3927_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_164 _4157_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_175 _5975_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_186 _7118_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_524 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_197 hold99/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5170_ hold211/X _5494_/A1 _5170_/S VGND VPWR _5170_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4121_ hold401/X _5526_/A1 _4126_/S VGND VPWR _4121_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4052_ _4110_/A0 _5473_/A1 _4058_/S VGND VPWR _4052_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xinput4 mask_rev_in[0] VGND VPWR input4/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4954_ _4413_/Y _4946_/X _5047_/A _5057_/B _4953_/Y VGND VPWR _4962_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_3905_ _4336_/C _4336_/D _4335_/A _4335_/B VGND VPWR _3906_/C VGND VPWR sky130_fd_sc_hd__nor4_1
X_4885_ _4884_/X _4839_/X _5006_/A _4885_/B2 VGND VPWR _6721_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6624_ _7150_/CLK _6624_/D fanout487/X VGND VPWR _6624_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3836_ _3836_/A _3836_/B VGND VPWR _6416_/D VGND VPWR sky130_fd_sc_hd__nor2_1
X_6555_ _6712_/CLK _6555_/D fanout470/X VGND VPWR _6555_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3767_ _7047_/Q _5505_/A _5166_/A _6751_/Q VGND VPWR _3767_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5506_ _5506_/A0 _5524_/A1 _5513_/S VGND VPWR _5506_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_106_616 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6486_ _3945_/A1 _6486_/D _6375_/X VGND VPWR _6486_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3698_ _3698_/A _3698_/B _3698_/C _3698_/D VGND VPWR _3699_/D VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_160_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput330 hold1373/X VGND VPWR hold1374/A VGND VPWR sky130_fd_sc_hd__buf_12
X_5437_ _5437_/A0 _5524_/A1 _5444_/S VGND VPWR _5437_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput341 hold1331/X VGND VPWR hold1332/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_105_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5368_ hold241/X _5494_/A1 _5372_/S VGND VPWR _5368_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7107_ _7126_/CLK _7107_/D fanout456/X VGND VPWR _7107_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4319_ hold954/X _6355_/A1 _4321_/S VGND VPWR _4319_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5299_ hold669/X _5521_/A1 _5300_/S VGND VPWR _5299_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7038_ _7038_/CLK _7038_/D fanout455/X VGND VPWR _7038_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_74_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_519 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_614 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_190 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4670_ _4928_/A _4676_/B VGND VPWR _4671_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_187_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3621_ _6981_/Q _5427_/A _4020_/A _6463_/Q VGND VPWR _3621_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6340_ _6339_/X _6340_/A1 _6346_/S VGND VPWR _7146_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3552_ _3552_/A _3552_/B _3552_/C _3552_/D VGND VPWR _3581_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_143_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6271_ _6458_/Q _5944_/X _5975_/A _6602_/Q _6270_/X VGND VPWR _6275_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3483_ _6895_/Q _5328_/A _5256_/A _6831_/Q _3482_/X VGND VPWR _3484_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5222_ hold289/X _5465_/A1 _5228_/S VGND VPWR _5222_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5153_ hold564/X _6357_/A1 _5153_/S VGND VPWR _5153_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_57_717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4104_ _4104_/A0 _5492_/A1 _4108_/S VGND VPWR _4104_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_111_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5084_ _5084_/A _5084_/B _5084_/C _5084_/D VGND VPWR _5085_/C VGND VPWR sky130_fd_sc_hd__and4_1
X_4035_ hold948/X _6355_/A1 _4037_/S VGND VPWR _4035_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5986_ _7039_/Q _5971_/C _5982_/X _5985_/X VGND VPWR _5989_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_169_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4937_ _4921_/A _4737_/A _4668_/C _4671_/A _4922_/X VGND VPWR _4996_/C VGND VPWR
+ sky130_fd_sc_hd__a311oi_2
XANTENNA_20 _3494_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_31 _3618_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4868_ _4846_/A _4672_/B _4643_/Y _4694_/Y _4442_/Y VGND VPWR _4869_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XANTENNA_42 _5300_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_53 _5948_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_64 _6051_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6607_ _6707_/CLK _6607_/D fanout447/X VGND VPWR _6607_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA_75 _6276_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3819_ _6555_/Q _4145_/A _3692_/Y _6767_/Q _3818_/X VGND VPWR _3826_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4799_ _4483_/Y _4673_/A _5008_/A _4798_/X VGND VPWR _4799_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XANTENNA_86 _7021_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_97 _6406_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_4_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6538_ _6735_/CLK _6538_/D _6360_/A VGND VPWR _6538_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_146_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6469_ _6654_/CLK hold69/X fanout454/X VGND VPWR _6469_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_121_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput171 _3958_/X VGND VPWR debug_in VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput182 _3207_/Y VGND VPWR mgmt_gpio_oeb[16] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput193 _3197_/Y VGND VPWR mgmt_gpio_oeb[26] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_75_514 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_296 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_761 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5840_ _6450_/Q _5634_/X _5829_/X _5833_/X _5839_/X VGND VPWR _5840_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_34_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5771_ _6871_/Q _5628_/X _5658_/X _6887_/Q VGND VPWR _5771_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_21_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4722_ _4722_/A _4722_/B _4722_/C _4722_/D VGND VPWR _4725_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_174_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4653_ _4716_/A _4653_/B _4653_/C VGND VPWR _4653_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_147_357 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput40 mgmt_gpio_in[13] VGND VPWR input40/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3604_ _3604_/A _3604_/B _3604_/C _3604_/D VGND VPWR _3604_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_162_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput51 mgmt_gpio_in[23] VGND VPWR input51/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput62 mgmt_gpio_in[33] VGND VPWR input62/X VGND VPWR sky130_fd_sc_hd__buf_2
Xhold802 _6966_/Q VGND VPWR hold802/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _4584_/A _5043_/A VGND VPWR _4942_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xinput73 pad_flash_io0_di VGND VPWR _3952_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput84 spimemio_flash_csb VGND VPWR input84/X VGND VPWR sky130_fd_sc_hd__buf_2
Xhold813 _4114_/X VGND VPWR _6528_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput95 usr1_vcc_pwrgood VGND VPWR input95/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xhold824 hold824/A VGND VPWR hold824/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ _6642_/Q _6323_/A2 _6323_/B1 _4230_/B VGND VPWR _6323_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3535_ hold36/X _3571_/B VGND VPWR _4286_/A VGND VPWR sky130_fd_sc_hd__nor2_2
Xhold835 _4312_/X VGND VPWR _6701_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _6456_/Q VGND VPWR hold846/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _5349_/X VGND VPWR _6908_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold868 _6892_/Q VGND VPWR hold868/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold879 _5484_/X VGND VPWR _7028_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _6278_/A0 _6253_/X _6279_/S VGND VPWR _6254_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3466_ _6983_/Q _5427_/A _5247_/A _6823_/Q _3460_/X VGND VPWR _3467_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5205_ _5205_/A0 _5484_/A1 _5210_/S VGND VPWR _5205_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6185_ _6630_/Q _5946_/X _5955_/X _6550_/Q VGND VPWR _6185_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3397_ _3959_/B _4083_/S _5211_/A _6793_/Q _3396_/X VGND VPWR _3409_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1502 _6028_/X VGND VPWR _7120_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1513 _7119_/Q VGND VPWR _6003_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5136_ _6726_/Q _4229_/X _5112_/X _5135_/Y VGND VPWR _5136_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_111_471 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1524 _7109_/Q VGND VPWR _5736_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 _6584_/Q VGND VPWR _4180_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1546 _7115_/Q VGND VPWR _5865_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _7132_/Q VGND VPWR hold1557/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _5134_/B _5066_/X _5006_/Y VGND VPWR _5067_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_57_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1568 _7093_/Q VGND VPWR _5575_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_506 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1579 _6416_/Q VGND VPWR _3835_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4018_ hold756/X _6356_/A1 _4019_/S VGND VPWR _4018_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_274 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5969_ _5969_/A _5979_/A _5969_/C VGND VPWR _5971_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_185_408 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_311 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold109 _3978_/X VGND VPWR _6424_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3320_ hold47/X _3453_/A hold64/X VGND VPWR _3320_/X VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_180_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3251_ _3251_/A _6485_/Q VGND VPWR _3262_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_98_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_555 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3182_ _6489_/Q VGND VPWR _3182_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_94_664 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_314 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6941_ _7054_/CLK _6941_/D fanout461/X VGND VPWR _6941_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_93_185 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6872_ _6920_/CLK _6872_/D fanout473/X VGND VPWR _6872_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_34_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5823_ _6470_/Q _5627_/X _5635_/X _6565_/Q VGND VPWR _5823_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_148_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5754_ _5754_/A _5754_/B _5754_/C VGND VPWR _5754_/Y VGND VPWR sky130_fd_sc_hd__nor3_2
X_4705_ _4689_/A _4644_/Y _4702_/Y _4673_/A _4704_/X VGND VPWR _4706_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5685_ _6979_/Q _5624_/X _5654_/X _6931_/Q _5684_/X VGND VPWR _5690_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4636_ _4636_/A _4646_/A VGND VPWR _4658_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_147_198 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold610 _6511_/Q VGND VPWR hold610/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold621 _3986_/X VGND VPWR _6430_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4567_ _4664_/B _4568_/B VGND VPWR _4737_/A VGND VPWR sky130_fd_sc_hd__and2b_2
Xhold632 _6841_/Q VGND VPWR hold632/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_563 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold643 _4259_/X VGND VPWR _6657_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap362 _3331_/Y VGND VPWR _5202_/B VGND VPWR sky130_fd_sc_hd__buf_6
Xhold654 _6929_/Q VGND VPWR hold654/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6636_/Q _3910_/B _6305_/Y _6306_/B2 VGND VPWR _7132_/D VGND VPWR sky130_fd_sc_hd__a22o_1
Xmax_cap373 _3555_/A VGND VPWR _3554_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold665 hold665/A VGND VPWR hold665/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3518_ _6474_/Q _4032_/A _4038_/A _6479_/Q VGND VPWR _3518_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_1_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xmax_cap384 _5657_/X VGND VPWR _5928_/A2 VGND VPWR sky130_fd_sc_hd__buf_8
Xhold676 _5354_/X VGND VPWR _6913_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4498_/A _4843_/B VGND VPWR _4498_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_143_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold687 _6801_/Q VGND VPWR hold687/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 _6983_/Q VGND VPWR hold698/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6452_/Q _5947_/X _5965_/X _6547_/Q _6236_/X VGND VPWR _6240_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3449_ _3448_/X _3449_/A1 _3829_/B VGND VPWR _6733_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6168_ _6825_/Q _5953_/X _5960_/X _7078_/Q _6167_/X VGND VPWR _6168_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_322 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1310 _4033_/X VGND VPWR _6470_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1321 hold1415/X VGND VPWR hold1321/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 hold1332/A VGND VPWR wb_dat_o[5] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_85_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1343 hold1427/X VGND VPWR hold1343/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5119_ _4465_/B _4644_/B _4975_/B _4450_/Y VGND VPWR _5120_/C VGND VPWR sky130_fd_sc_hd__a31oi_1
XFILLER_84_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1354 hold1354/A VGND VPWR wb_dat_o[12] VGND VPWR sky130_fd_sc_hd__buf_12
X_6099_ _6099_/A _6099_/B _6099_/C _6099_/D VGND VPWR _6100_/C VGND VPWR sky130_fd_sc_hd__nor4_1
Xhold1365 _4189_/A1 VGND VPWR hold1365/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_528 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1376 hold1376/A VGND VPWR wb_dat_o[4] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1387 _7060_/Q VGND VPWR _5520_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 _7145_/Q VGND VPWR _3973_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_46 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VPWR _7113_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_391 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_646 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_599 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_388 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_400 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_102 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5470_ hold750/X _5521_/A1 _5471_/S VGND VPWR _5470_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_124 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4421_ _4753_/A _4607_/A VGND VPWR _4626_/B VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_172_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7140_ _7140_/CLK _7140_/D VGND VPWR _7140_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_4352_ _4633_/B _4352_/B VGND VPWR _4360_/B VGND VPWR sky130_fd_sc_hd__xor2_1
XFILLER_125_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout408 _5509_/A1 VGND VPWR _5545_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_3303_ hold26/X hold46/X VGND VPWR _3303_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
Xfanout419 _5534_/A1 VGND VPWR _5543_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_7071_ _7083_/CLK _7071_/D fanout470/X VGND VPWR _7071_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4283_ _4283_/A0 _5493_/A1 _4285_/S VGND VPWR _4283_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6022_ _6443_/Q _5601_/X _5959_/X _6963_/Q VGND VPWR _6022_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3234_ _6415_/Q _6485_/Q _3234_/C VGND VPWR _3235_/S VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_67_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3165_ _7158_/Q VGND VPWR _3165_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_163 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_528 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6924_ _7006_/CLK _6924_/D fanout458/X VGND VPWR _6924_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_81_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6855_ _6865_/CLK _6855_/D fanout464/X VGND VPWR _6855_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5806_ _7009_/Q _5625_/X _5661_/X _6881_/Q VGND VPWR _5806_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6786_ _7006_/CLK _6786_/D fanout456/X VGND VPWR _6786_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_10_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3998_ hold523/X _5513_/A1 _3998_/S VGND VPWR _3998_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_148_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5737_ _6958_/Q _5638_/X _5661_/X _6878_/Q VGND VPWR _5737_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_13_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5668_ _6890_/Q _5666_/X _5667_/X _6810_/Q _5665_/X VGND VPWR _5669_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_190_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4619_ _4716_/A _4653_/B _4635_/B VGND VPWR _4619_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_151_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5599_ _5597_/B _5598_/Y _5602_/B VGND VPWR _7101_/D VGND VPWR sky130_fd_sc_hd__a21oi_1
Xhold440 _5441_/X VGND VPWR _6990_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold451 _6806_/Q VGND VPWR hold451/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _4235_/X VGND VPWR _6627_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold473 _6918_/Q VGND VPWR hold473/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold484 _5510_/X VGND VPWR _7051_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _6617_/Q VGND VPWR hold495/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1140 _5191_/X VGND VPWR _6768_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1151 _6866_/Q VGND VPWR _5302_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _5473_/X VGND VPWR _7018_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _6555_/Q VGND VPWR _4146_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_111 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1184 _4015_/X VGND VPWR _6455_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 _6850_/Q VGND VPWR _5284_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_168 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_371 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_503 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4970_ _4970_/A _4975_/B VGND VPWR _4970_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_91_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3921_ _3187_/Y input90/X _3921_/S VGND VPWR _3921_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_44_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6640_ _7150_/CLK _6640_/D fanout487/X VGND VPWR _6640_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3852_ _3852_/A _3860_/B VGND VPWR _3853_/B VGND VPWR sky130_fd_sc_hd__nand2_1
X_6571_ _7137_/CLK _6571_/D VGND VPWR _6571_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3783_ _6685_/Q _4292_/A _5490_/A _7034_/Q VGND VPWR _3783_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_118_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5522_ hold313/X _5540_/A1 hold87/X VGND VPWR _5522_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5453_ hold497/X hold22/X _5453_/S VGND VPWR _5453_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4404_ _4408_/B _4448_/B VGND VPWR _4549_/A VGND VPWR sky130_fd_sc_hd__nor2_4
X_5384_ hold301/X _5465_/A1 _5390_/S VGND VPWR _5384_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7123_ _7131_/CLK _7123_/D fanout459/X VGND VPWR _7123_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4335_ _4335_/A _4335_/B _4335_/C _4335_/D VGND VPWR _4338_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_87_715 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_363 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7054_ _7054_/CLK _7054_/D fanout461/X VGND VPWR _7054_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4266_ hold347/X _5518_/A1 _4267_/S VGND VPWR _4266_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_57_csclk _6447_/CLK VGND VPWR _6925_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6005_ _6859_/Q _5943_/X _5981_/X _6915_/Q VGND VPWR _6005_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3217_ _6837_/Q VGND VPWR _3217_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4197_ hold976/X hold666/X _4201_/S VGND VPWR _4197_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_54_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6907_ _7082_/CLK _6907_/D fanout479/X VGND VPWR _6907_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_6838_ _7026_/CLK _6838_/D fanout463/X VGND VPWR _6838_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_7_708 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6769_ _6769_/CLK _6769_/D fanout469/X VGND VPWR _6769_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_7_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold270 _4288_/X VGND VPWR _6681_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6556_/Q VGND VPWR hold281/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _5209_/X VGND VPWR _6784_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_110 _3956_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_121 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_132 _6747_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_143 _5902_/A2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_154 hold6/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_165 _4238_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_176 _5960_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_187 _3957_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_198 _5171_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4120_ hold824/X _6354_/A1 _4126_/S VGND VPWR _4120_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_123_694 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4051_ _6396_/B _3692_/A hold37/X _4050_/X _4322_/B VGND VPWR _4067_/S VGND VPWR
+ sky130_fd_sc_hd__o221a_4
XFILLER_83_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VPWR input5/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_91_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4953_ _4953_/A _5043_/B VGND VPWR _4953_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_51_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3904_ _4335_/C _4335_/D _3904_/C VGND VPWR _3906_/B VGND VPWR sky130_fd_sc_hd__nor3_1
X_4884_ _5006_/A _4884_/B _4884_/C _4884_/D VGND VPWR _4884_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_6623_ _6712_/CLK _6623_/D _6390_/A VGND VPWR _6623_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3835_ _3835_/A _3838_/A VGND VPWR _3836_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_20_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6554_ _6674_/CLK _6554_/D _6383_/A VGND VPWR _6554_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_20_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3766_ input52/X _5193_/A _4220_/A _6619_/Q _3765_/X VGND VPWR _3773_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5505_ _5505_/A _5505_/B VGND VPWR _5513_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_173_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6485_ _3927_/A1 _6485_/D _6374_/X VGND VPWR _6485_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_118_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3697_ _6820_/Q _5247_/A _4298_/A _6692_/Q _3696_/X VGND VPWR _3698_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_628 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5436_ _5436_/A _5505_/B VGND VPWR _5444_/S VGND VPWR sky130_fd_sc_hd__and2_4
Xoutput320 hold1339/X VGND VPWR hold1340/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_105_138 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput331 hold1363/X VGND VPWR hold1364/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_161_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xoutput342 hold1335/X VGND VPWR hold1336/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_121_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5367_ hold325/X _5526_/A1 _5372_/S VGND VPWR _5367_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7106_ _7126_/CLK _7106_/D fanout456/X VGND VPWR _7106_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_114_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4318_ hold814/X _6354_/A1 _4321_/S VGND VPWR _4318_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5298_ hold160/X hold42/X _5300_/S VGND VPWR _5298_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7037_ _7037_/CLK _7037_/D fanout450/X VGND VPWR _7037_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_75_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4249_ hold525/X _5546_/A1 _4249_/S VGND VPWR _4249_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_250 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_325 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3620_ _3620_/A _3620_/B _3620_/C _3620_/D VGND VPWR _3639_/A VGND VPWR sky130_fd_sc_hd__nor4_1
X_3551_ _6830_/Q _5256_/A _4196_/A _6603_/Q _3549_/X VGND VPWR _3552_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6270_ _6468_/Q _5937_/X _5975_/D _6628_/Q VGND VPWR _6270_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_182_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3482_ input57/X _5193_/A _5541_/A _7084_/Q VGND VPWR _3482_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5221_ _5221_/A0 _5524_/A1 _5228_/S VGND VPWR _5221_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5152_ hold728/X _6356_/A1 _5153_/S VGND VPWR _5152_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4103_ _4103_/A0 _5491_/A1 _4108_/S VGND VPWR _4103_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5083_ _5083_/A _5083_/B _5083_/C VGND VPWR _5115_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_111_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4034_ hold876/X _6354_/A1 _4037_/S VGND VPWR _4034_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_65_740 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5985_ _7018_/Q _5937_/X _5944_/X _7026_/Q _5984_/X VGND VPWR _5985_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XPHY_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4936_ _4999_/B _5003_/B _5076_/A VGND VPWR _4944_/B VGND VPWR sky130_fd_sc_hd__and3_1
XANTENNA_10 _3355_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_21 _3504_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4867_ _4902_/B _4639_/Y _4508_/C VGND VPWR _5027_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA_32 _3638_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_43 _5399_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_54 _5976_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6606_ _6746_/CLK _6606_/D fanout447/X VGND VPWR _6606_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3818_ _6898_/Q _5337_/A _4232_/A _6625_/Q VGND VPWR _3818_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XANTENNA_65 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_76 _6276_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4798_ _4627_/B _4638_/Y _4673_/A _4627_/A VGND VPWR _4798_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XANTENNA_87 _7040_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_98 _7157_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6537_ _6537_/CLK _6537_/D fanout464/X VGND VPWR _6537_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_134_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3749_ _6835_/Q _5265_/A _4008_/A _6451_/Q VGND VPWR _3749_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_21_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6468_ _6654_/CLK _6468_/D _6401_/A VGND VPWR _6468_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_161_542 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5419_ _5419_/A0 _5524_/A1 _5426_/S VGND VPWR _5419_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_121_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6399_ _6401_/A _6401_/B VGND VPWR _6399_/X VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput172 _7173_/X VGND VPWR irq[0] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput183 _3206_/Y VGND VPWR mgmt_gpio_oeb[17] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput194 _3196_/Y VGND VPWR mgmt_gpio_oeb[27] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_762 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_507 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_572 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_726 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_480 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5770_ _6983_/Q _5624_/X _5634_/X _6975_/Q _5758_/Y VGND VPWR _5770_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_159_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4721_ _4721_/A _4721_/B _4721_/C VGND VPWR _4722_/D VGND VPWR sky130_fd_sc_hd__and3_1
X_4652_ _4653_/B _4653_/C VGND VPWR _4652_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_147_369 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput30 mask_rev_in[4] VGND VPWR input30/X VGND VPWR sky130_fd_sc_hd__buf_2
X_3603_ _6805_/Q _5229_/A _4145_/A _6558_/Q _3588_/X VGND VPWR _3604_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xinput41 mgmt_gpio_in[14] VGND VPWR input41/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput52 mgmt_gpio_in[24] VGND VPWR input52/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
X_4583_ _4581_/B _4582_/Y _4810_/A VGND VPWR _4583_/X VGND VPWR sky130_fd_sc_hd__a21o_1
Xinput63 mgmt_gpio_in[34] VGND VPWR _3957_/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_162_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold803 _5414_/X VGND VPWR _6966_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VPWR _3953_/B VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold814 _6706_/Q VGND VPWR hold814/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _6643_/Q _6319_/Y _6321_/X _6317_/Y VGND VPWR _6346_/S VGND VPWR sky130_fd_sc_hd__a211o_4
Xinput85 spimemio_flash_io0_do VGND VPWR input85/X VGND VPWR sky130_fd_sc_hd__buf_2
Xhold825 _4120_/X VGND VPWR _6533_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3534_ _6741_/Q _5148_/A hold67/A _6469_/Q _3531_/X VGND VPWR _3538_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_531 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput96 usr1_vdd_pwrgood VGND VPWR input96/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold836 _7152_/Q VGND VPWR hold836/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _4016_/X VGND VPWR _6456_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _7191_/A VGND VPWR hold858/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 _5331_/X VGND VPWR _6892_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ _7128_/Q _6252_/X _6303_/S VGND VPWR _6253_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3465_ _6863_/Q _5292_/A _5154_/A _6747_/Q _3464_/X VGND VPWR _3467_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5204_ hold257/X _5534_/A1 _5210_/S VGND VPWR _5204_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6184_ _6685_/Q _5961_/X _6182_/X _6183_/X VGND VPWR _6189_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3396_ _6441_/Q _3372_/Y _3393_/X _3395_/X VGND VPWR _3396_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_97_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1503 _7130_/Q VGND VPWR _6279_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5135_ _5135_/A _5135_/B _5135_/C VGND VPWR _5135_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
Xhold1514 _7147_/Q VGND VPWR _6343_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1525 hold58/A VGND VPWR _3257_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_483 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1536 hold40/A VGND VPWR _3256_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 _6489_/Q VGND VPWR _3912_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 hold32/A VGND VPWR _3849_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5066_ _5066_/A _5112_/C _5106_/C _5066_/D VGND VPWR _5066_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_38_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1569 _7167_/Q VGND VPWR _3253_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ hold960/X _6355_/A1 _4019_/S VGND VPWR _4017_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5968_ _5968_/A _5969_/C _5979_/C VGND VPWR _5976_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_52_286 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4919_ _5023_/A _5023_/B _5023_/C _4919_/D VGND VPWR _4919_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_21_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5899_ _6658_/Q _5899_/B VGND VPWR _5899_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_166_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_306 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_684 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_323 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_584 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3250_ _3250_/A _3250_/B VGND VPWR _7168_/D VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_112_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_567 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3181_ _4566_/A VGND VPWR _4702_/B VGND VPWR sky130_fd_sc_hd__clkinv_2
XFILLER_79_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_676 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6940_ _7063_/CLK _6940_/D fanout463/X VGND VPWR _6940_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_81_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6871_ _7078_/CLK _6871_/D fanout482/X VGND VPWR _6871_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_179_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_404 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5822_ _3183_/Y _5899_/B _5651_/B VGND VPWR _5822_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_34_275 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5753_ _7006_/Q _5625_/X _5632_/X _6942_/Q _5737_/X VGND VPWR _5754_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4704_ _4460_/A _4626_/B _4616_/Y _4703_/Y VGND VPWR _4704_/X VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_148_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5684_ _6971_/Q _5634_/X _5652_/B _6915_/Q _5651_/Y VGND VPWR _5684_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4635_ _4716_/A _4635_/B _4661_/B VGND VPWR _4689_/B VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_162_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold600 _7056_/Q VGND VPWR hold600/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 _4089_/X VGND VPWR _6511_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4566_ _4566_/A _4566_/B VGND VPWR _4664_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
Xhold622 hold622/A VGND VPWR hold622/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold633 _5273_/X VGND VPWR _6841_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _7080_/Q VGND VPWR hold644/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6636_/Q _6641_/Q _6635_/Q _3910_/B VGND VPWR _6305_/Y VGND VPWR sky130_fd_sc_hd__o31ai_1
XFILLER_89_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xmax_cap363 _4118_/B VGND VPWR _4083_/S VGND VPWR sky130_fd_sc_hd__buf_8
X_3517_ hold74/X _3573_/B VGND VPWR _4038_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_116_575 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold655 _5372_/X VGND VPWR _6929_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 hold666/A VGND VPWR hold666/X VGND VPWR sky130_fd_sc_hd__buf_8
Xmax_cap374 _3571_/A VGND VPWR hold125/A VGND VPWR sky130_fd_sc_hd__buf_12
X_4497_ _4579_/B _5042_/B VGND VPWR _4843_/B VGND VPWR sky130_fd_sc_hd__and2_1
Xmax_cap385 _5655_/X VGND VPWR _5905_/A2 VGND VPWR sky130_fd_sc_hd__buf_6
Xhold677 _6969_/Q VGND VPWR hold677/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold688 _5228_/X VGND VPWR _6801_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 _5433_/X VGND VPWR _6983_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6236_ _6632_/Q _5946_/X _5955_/X _6552_/Q VGND VPWR _6236_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3448_ _3447_/Y _3488_/A1 _3829_/A VGND VPWR _3448_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6167_ _6913_/Q _5973_/A _5948_/X _6953_/Q _6166_/X VGND VPWR _6167_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1300 _5149_/X VGND VPWR _6737_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3379_ _3379_/A hold75/X VGND VPWR _3999_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1311 _6418_/Q VGND VPWR _3966_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 hold1322/A VGND VPWR wb_dat_o[19] VGND VPWR sky130_fd_sc_hd__buf_12
X_5118_ _5118_/A _5118_/B _5118_/C VGND VPWR _5118_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_111_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1333 hold1419/X VGND VPWR hold1333/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 hold1344/A VGND VPWR wb_dat_o[13] VGND VPWR sky130_fd_sc_hd__buf_12
Xclkbuf_0__1177_ _3582_/Y VGND VPWR clkbuf_0__1177_/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6098_ _6814_/Q _5971_/B _5949_/X _6934_/Q _6097_/X VGND VPWR _6099_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1355 _6315_/A1 VGND VPWR hold1355/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1366 hold1366/A VGND VPWR wb_dat_o[1] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1377 _6312_/A1 VGND VPWR hold1377/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _4672_/B _4496_/Y _4542_/A VGND VPWR _5049_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_27_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1388 _7084_/Q VGND VPWR _5547_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 _3973_/X VGND VPWR hold59/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_58 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_770 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_531 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_323 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_315 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_592 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4420_ _4753_/A _4600_/B VGND VPWR _4947_/A VGND VPWR sky130_fd_sc_hd__nand2b_2
XFILLER_144_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4351_ _4352_/B _4351_/B VGND VPWR _4379_/B VGND VPWR sky130_fd_sc_hd__nand2_1
X_3302_ hold72/X _3355_/B _3347_/A VGND VPWR _3555_/A VGND VPWR sky130_fd_sc_hd__nand3b_4
Xfanout409 _5518_/A1 VGND VPWR _5509_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_7070_ _7070_/CLK _7070_/D fanout482/X VGND VPWR _7070_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4282_ _4282_/A0 _5492_/A1 _4285_/S VGND VPWR _4282_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6021_ _7027_/Q _5944_/X _5975_/A _6843_/Q _6020_/X VGND VPWR _6024_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3233_ _3233_/A0 _3251_/A _3233_/S VGND VPWR _7171_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_csclk clkbuf_1_1_1_csclk/A VGND VPWR clkbuf_2_3_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
X_3164_ _7159_/Q VGND VPWR _3164_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_67_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_175 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6923_ _7006_/CLK _6923_/D fanout458/X VGND VPWR _6923_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_35_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6854_ _7081_/CLK _6854_/D fanout478/X VGND VPWR _6854_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5805_ _6953_/Q _5637_/X _5645_/X _7033_/Q VGND VPWR _5805_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6785_ _7076_/CLK _6785_/D fanout481/X VGND VPWR _6785_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3997_ _3997_/A0 hold99/X _3998_/S VGND VPWR _3997_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5736_ _5736_/A1 _6279_/S _5734_/X _5735_/X VGND VPWR _7109_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_148_442 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5667_ _5664_/A _5667_/B _5667_/C VGND VPWR _5667_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_135_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4618_ _4653_/B _4635_/B VGND VPWR _4618_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_163_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5598_ _5598_/A _5602_/A VGND VPWR _5598_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_190_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold430 _5343_/X VGND VPWR _6903_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _6765_/Q VGND VPWR hold441/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4549_/A _4549_/B VGND VPWR _4553_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_89_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold452 _5234_/X VGND VPWR _6806_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _6563_/Q VGND VPWR hold463/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 _5360_/X VGND VPWR _6918_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold485 _6910_/Q VGND VPWR hold485/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold496 _4218_/X VGND VPWR _6617_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6219_ _6646_/Q _5976_/C _5971_/D _6566_/Q VGND VPWR _6219_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_77_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7199_ _7199_/A VGND VPWR _7199_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_621 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1130 _4160_/X VGND VPWR _6567_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _6767_/Q VGND VPWR _5189_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 _5302_/X VGND VPWR _6866_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 _6465_/Q VGND VPWR _4027_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _4146_/X VGND VPWR _6555_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _6882_/Q VGND VPWR _5320_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1196 _5284_/X VGND VPWR _6850_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_166_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_757 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_318 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3920_ _3186_/Y input92/X _3921_/S VGND VPWR _3920_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_32_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3851_ _3850_/Y hold70/A _3851_/C VGND VPWR _3853_/A VGND VPWR sky130_fd_sc_hd__and3b_1
X_6570_ _7137_/CLK _6570_/D VGND VPWR _6570_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3782_ _3782_/A _3782_/B _3782_/C _3782_/D VGND VPWR _3794_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_164_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5521_ hold319/X _5521_/A1 hold87/X VGND VPWR _5521_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5452_ hold112/X hold99/X _5453_/S VGND VPWR _5452_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_765 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4403_ _4633_/B _4389_/Y _4653_/B _4563_/D VGND VPWR _4448_/B VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_145_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5383_ _5383_/A0 hold666/X _5390_/S VGND VPWR _5383_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7122_ _7131_/CLK _7122_/D fanout456/X VGND VPWR _7122_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4334_ _4702_/A _4334_/B _4334_/C VGND VPWR _4434_/B VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_5_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7053_ _7053_/CLK _7053_/D fanout459/X VGND VPWR _7053_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4265_ hold471/X _5544_/A1 _4267_/S VGND VPWR _4265_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6004_ _7040_/Q _5971_/C _5976_/D _6875_/Q VGND VPWR _6004_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3216_ _6845_/Q VGND VPWR _3216_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4196_ _4196_/A _4322_/B VGND VPWR _4201_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_27_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6906_ _6908_/CLK _6906_/D fanout463/X VGND VPWR _6906_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_23_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6837_ _6865_/CLK _6837_/D fanout464/X VGND VPWR _6837_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_145_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_738 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6768_ _6769_/CLK _6768_/D fanout469/X VGND VPWR _6768_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5719_ _7005_/Q _5625_/X _5661_/X _6877_/Q VGND VPWR _5719_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6699_ _6709_/CLK _6699_/D _6360_/A VGND VPWR _6699_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_108_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold260 _5447_/X VGND VPWR _6995_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _6752_/Q VGND VPWR hold271/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _4147_/X VGND VPWR _6556_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_727 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold293 _6851_/Q VGND VPWR hold293/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_100 _7157_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_111 _7199_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_122 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_133 _6739_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_33_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_144 _5902_/A2 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_155 hold60/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_166 _5166_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_177 _5975_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_188 input46/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_199 _5229_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_174_507 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4050_ _6396_/B _5193_/A VGND VPWR _4050_/X VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_49_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput6 mask_rev_in[11] VGND VPWR input6/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4952_ _4542_/B _5043_/B VGND VPWR _5057_/B VGND VPWR sky130_fd_sc_hd__nand2b_1
X_3903_ _4337_/C _4337_/D _4336_/A _4336_/B VGND VPWR _3907_/C VGND VPWR sky130_fd_sc_hd__nor4_1
X_4883_ _5023_/C _4882_/X _5023_/A VGND VPWR _4884_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
X_6622_ _6629_/CLK _6622_/D _6390_/A VGND VPWR _6622_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3834_ _3867_/B _3832_/B _3836_/A _3834_/B2 VGND VPWR _6417_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_118_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6553_ _6659_/CLK _6553_/D fanout469/X VGND VPWR _6553_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_326 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3765_ _7018_/Q hold29/A _5409_/A _6962_/Q VGND VPWR _3765_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5504_ hold311/X _5540_/A1 hold77/X VGND VPWR _5504_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6484_ _6707_/CLK _6484_/D fanout450/X VGND VPWR _6484_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3696_ _6621_/Q _4220_/A _4244_/A _6647_/Q VGND VPWR _3696_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_702 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xpad_flashh_clk_buff_inst _3945_/X VGND VPWR pad_flash_clk VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_5435_ hold143/X hold22/X _5435_/S VGND VPWR _5435_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput310 _3953_/X VGND VPWR spimemio_flash_io1_di VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput321 hold1351/X VGND VPWR hold1352/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput332 hold1357/X VGND VPWR hold1358/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput343 hold1337/X VGND VPWR hold1338/A VGND VPWR sky130_fd_sc_hd__buf_12
X_5366_ hold245/X _5465_/A1 _5372_/S VGND VPWR _5366_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7105_ _7113_/CLK _7105_/D fanout460/X VGND VPWR _7105_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4317_ _4317_/A0 _5491_/A1 _4321_/S VGND VPWR _4317_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5297_ hold180/X _5519_/A1 _5300_/S VGND VPWR _5297_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7036_ _7036_/CLK _7036_/D fanout455/X VGND VPWR _7036_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_59_259 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4248_ hold491/X _5518_/A1 _4249_/S VGND VPWR _4248_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4179_ _3828_/Y _4179_/A1 _4186_/S VGND VPWR _6583_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_23 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_570 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_602 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_csclk clkbuf_opt_3_0_csclk/X VGND VPWR _6967_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_178_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk _6447_/CLK VGND VPWR _6539_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3550_ _3562_/A _3692_/A VGND VPWR _4196_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_143_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3481_ _6855_/Q _5283_/A _5202_/B input40/X _3480_/X VGND VPWR _3484_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5220_ _5220_/A hold17/X VGND VPWR _5227_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_407 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5151_ hold995/X _6355_/A1 _5153_/S VGND VPWR _5151_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4102_ _4102_/A _5541_/B VGND VPWR _4108_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_5082_ _5088_/A _5114_/A _5082_/C VGND VPWR _5087_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_84_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4033_ _4033_/A0 _5491_/A1 _4037_/S VGND VPWR _4033_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5984_ _6794_/Q _5965_/X _5971_/D _6826_/Q VGND VPWR _5984_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_169_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4935_ _4948_/C _4562_/Y _4620_/Y _4638_/Y _4768_/B VGND VPWR _5076_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_3_7_0_csclk clkbuf_3_7_0_csclk/A VGND VPWR clkbuf_3_7_0_csclk/X VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_33_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_11 _5265_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_22 _4220_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4866_ _4948_/C _4496_/Y _4639_/Y _4689_/A VGND VPWR _4870_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_177_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_33 _3688_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_44 _5471_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6605_ _6746_/CLK _6605_/D fanout447/X VGND VPWR _6605_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XANTENNA_55 _5958_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3817_ _3817_/A _3817_/B _3817_/C _3817_/D VGND VPWR _3827_/C VGND VPWR sky130_fd_sc_hd__nor4_1
XANTENNA_66 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_165_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4797_ _4673_/A _4611_/Y _4476_/Y VGND VPWR _5008_/A VGND VPWR sky130_fd_sc_hd__a21o_1
XANTENNA_77 _6276_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_88 _7040_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6536_ _6539_/CLK _6536_/D fanout461/X VGND VPWR _6536_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3748_ _6661_/Q _4262_/A _4127_/A _6541_/Q _3747_/X VGND VPWR _3751_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XANTENNA_99 _7157_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6467_ _6654_/CLK _6467_/D _6401_/A VGND VPWR _6467_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3679_ _3679_/A _3679_/B _3679_/C _3679_/D VGND VPWR _3699_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_134_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5418_/A _5541_/B VGND VPWR _5426_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_6398_ _6401_/A _6401_/B VGND VPWR _6398_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_121_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput173 _3959_/X VGND VPWR irq[1] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput184 _3205_/Y VGND VPWR mgmt_gpio_oeb[18] VGND VPWR sky130_fd_sc_hd__buf_12
X_5349_ hold856/X _5484_/A1 _5354_/S VGND VPWR _5349_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput195 _3195_/Y VGND VPWR mgmt_gpio_oeb[28] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_36 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7019_ _7085_/CLK _7019_/D fanout479/X VGND VPWR _7019_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_28_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_424 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_242 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_223 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_492 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4720_ _4689_/A _4616_/Y _4626_/Y _4483_/Y _4719_/X VGND VPWR _4721_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_159_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4651_ _4441_/A _4484_/Y _4609_/Y _4619_/Y _4650_/Y VGND VPWR _4660_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_147_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput20 mask_rev_in[24] VGND VPWR input20/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_3602_ _6917_/Q _5355_/A _5247_/A _6821_/Q _3601_/X VGND VPWR _3604_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xinput31 mask_rev_in[5] VGND VPWR input31/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4582_ _4992_/A _4582_/B VGND VPWR _4582_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VPWR input42/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VPWR input53/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_128_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput64 mgmt_gpio_in[35] VGND VPWR input64/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput75 porb VGND VPWR input75/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xhold804 _6435_/Q VGND VPWR hold804/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6321_ _6642_/Q _6318_/Y _6320_/Y _6644_/Q _4229_/X VGND VPWR _6321_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3533_ hold74/A hold66/X VGND VPWR hold67/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xinput86 spimemio_flash_io0_oeb VGND VPWR _3947_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xhold815 _4318_/X VGND VPWR _6706_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 _6714_/Q VGND VPWR hold826/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput97 usr2_vcc_pwrgood VGND VPWR input97/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xhold837 _6354_/X VGND VPWR _7152_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold848 _6481_/Q VGND VPWR hold848/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ _6240_/Y _6251_/X _6542_/Q _6226_/B VGND VPWR _6252_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
Xhold859 _5196_/X VGND VPWR _6772_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3464_ _6911_/Q _5346_/A _5391_/A _6951_/Q VGND VPWR _3464_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5203_ _5203_/A0 _5473_/A1 _5210_/S VGND VPWR _5203_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6183_ _6475_/Q _5940_/X _5967_/X _6604_/Q _6181_/X VGND VPWR _6183_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3395_ _6865_/Q _5292_/A _5532_/A _7078_/Q _3394_/X VGND VPWR _3395_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_4
X_5134_ _5134_/A _5134_/B _5134_/C VGND VPWR _5135_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_97_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1504 _7124_/Q VGND VPWR _6129_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1515 _7145_/Q VGND VPWR _6337_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _3257_/X VGND VPWR _7163_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1537 _7112_/Q VGND VPWR _5820_/A2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5065_ _4483_/Y _4625_/B _4650_/Y _4716_/Y _5018_/A VGND VPWR _5066_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
Xhold1548 _3182_/Y VGND VPWR _3869_/A2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 _6635_/Q VGND VPWR _3909_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4016_ hold846/X _6354_/A1 _4019_/S VGND VPWR _4016_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5967_ _5969_/C _5981_/C _5979_/C VGND VPWR _5967_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_52_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4918_ _4918_/A _4918_/B VGND VPWR _4919_/D VGND VPWR sky130_fd_sc_hd__nand2_1
X_5898_ _6563_/Q _5631_/X _5637_/X _6698_/Q _5897_/X VGND VPWR _5906_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4849_ _4483_/Y _4846_/B _4535_/A VGND VPWR _5073_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_193_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6519_ _6668_/CLK _6519_/D _6400_/A VGND VPWR _6519_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_180_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_357 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_596 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3180_ _7101_/Q VGND VPWR _5600_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_140_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_335 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6870_ _7051_/CLK _6870_/D fanout476/X VGND VPWR _6870_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_34_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5821_ _5821_/A1 _6279_/S _5819_/X _5820_/X VGND VPWR _7113_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_50_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_287 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5752_ _7014_/Q _5630_/X _5645_/X _7030_/Q _5751_/X VGND VPWR _5754_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4703_ _4782_/A _4703_/B VGND VPWR _4703_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_30_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5683_ _6923_/Q _5664_/X _5667_/X _6811_/Q _5682_/X VGND VPWR _5690_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4634_ _4716_/A _4635_/B _4661_/B VGND VPWR _4753_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_163_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold601 _5516_/X VGND VPWR _7056_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4563_/D _4653_/B _4595_/A VGND VPWR _4565_/X VGND VPWR sky130_fd_sc_hd__a21o_1
Xhold612 _6672_/Q VGND VPWR hold612/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold623 _4111_/X VGND VPWR _6525_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _6971_/Q VGND VPWR hold634/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6304_/A0 _6303_/X _6304_/S VGND VPWR _7131_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold645 _5543_/X VGND VPWR _7080_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _3573_/A _3814_/B VGND VPWR _4032_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold656 _7015_/Q VGND VPWR hold656/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _4607_/A _4496_/B VGND VPWR _4496_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold667 hold667/A VGND VPWR hold667/X VGND VPWR sky130_fd_sc_hd__buf_8
Xmax_cap386 _5646_/X VGND VPWR _5814_/B1 VGND VPWR sky130_fd_sc_hd__buf_8
Xhold678 _5417_/X VGND VPWR _6969_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold689 _6423_/Q VGND VPWR hold689/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6687_/Q _5961_/X _6232_/X _6234_/X VGND VPWR _6240_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3447_ _3447_/A _3447_/B _3447_/C VGND VPWR _3447_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_6166_ _6905_/Q _5976_/C _5971_/D _6833_/Q VGND VPWR _6166_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3378_ _3586_/A hold75/X VGND VPWR hold76/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_69_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1301 _6434_/Q VGND VPWR _3991_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1312 _3966_/X VGND VPWR _6418_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1323 hold1416/X VGND VPWR hold1323/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _4482_/B _4695_/Y _4858_/X _4823_/A VGND VPWR _5118_/C VGND VPWR sky130_fd_sc_hd__o211a_1
Xhold1334 hold1334/A VGND VPWR wb_dat_o[11] VGND VPWR sky130_fd_sc_hd__buf_12
X_6097_ hold79/A _5601_/X _5959_/X _6966_/Q VGND VPWR _6097_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold1345 hold1428/X VGND VPWR hold1345/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 hold1356/A VGND VPWR wb_dat_o[31] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1367 _4190_/A1 VGND VPWR hold1367/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _4672_/B _4496_/Y _4413_/Y VGND VPWR _5057_/C VGND VPWR sky130_fd_sc_hd__a21o_1
Xhold1378 hold1378/A VGND VPWR wb_dat_o[28] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1389 _6788_/Q VGND VPWR _5214_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6999_ _6999_/CLK _6999_/D fanout465/X VGND VPWR _6999_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_43_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_471 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_671 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_419 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4350_ _4661_/A _4357_/B _4631_/D VGND VPWR _4351_/B VGND VPWR sky130_fd_sc_hd__a21o_1
X_3301_ _3586_/A _3562_/A VGND VPWR _5283_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_4281_ _4281_/A0 _6353_/A1 _4285_/S VGND VPWR _4281_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6020_ _7019_/Q _5937_/X _5975_/D _6883_/Q VGND VPWR _6020_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3232_ _3867_/A _3829_/A VGND VPWR _3233_/S VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_140_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_658 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6922_ _6926_/CLK _6922_/D fanout458/X VGND VPWR _6922_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_120_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6853_ _6951_/CLK _6853_/D fanout474/X VGND VPWR _6853_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_35_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5804_ _6849_/Q _5616_/X _5655_/X _6801_/Q _5803_/X VGND VPWR _5804_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6784_ _7076_/CLK _6784_/D fanout481/X VGND VPWR _6784_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3996_ hold574/X _5469_/A1 _3998_/S VGND VPWR _3996_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5735_ _6507_/Q _5735_/A2 _6103_/B1 VGND VPWR _5735_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_30_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_616 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5666_ _5664_/A _5666_/B _5666_/C VGND VPWR _5666_/X VGND VPWR sky130_fd_sc_hd__and3b_4
X_4617_ _4627_/A _4846_/B VGND VPWR _4646_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_135_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5597_ _5600_/A _5597_/B VGND VPWR _5602_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold420 _5535_/X VGND VPWR _7073_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6712_/Q VGND VPWR hold431/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _4500_/A _4947_/C _4464_/Y _4902_/A _5114_/A VGND VPWR _4548_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold442 _5187_/X VGND VPWR _6765_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _6557_/Q VGND VPWR hold453/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _4155_/X VGND VPWR _6563_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _6870_/Q VGND VPWR hold475/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _5351_/X VGND VPWR _6910_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _4653_/C VGND VPWR _4479_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_104_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold497 _7001_/Q VGND VPWR hold497/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6218_/A _6218_/B _6218_/C VGND VPWR _6226_/C VGND VPWR sky130_fd_sc_hd__nor3_1
X_7198_ _7198_/A VGND VPWR _7198_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_58_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1120 _5493_/X VGND VPWR _7036_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _6816_/Q _5971_/B _5949_/X _6936_/Q _6148_/X VGND VPWR _6150_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_666 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1131 _6580_/Q VGND VPWR _4175_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1142 _5189_/X VGND VPWR _6767_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 _6826_/Q VGND VPWR _5257_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1164 _4027_/X VGND VPWR _6465_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 hold1590/X VGND VPWR _4053_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 _5320_/X VGND VPWR _6882_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1197 _6888_/Q VGND VPWR _5326_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_332 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_633 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3850_ _6488_/Q _3854_/S VGND VPWR _3850_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_3781_ _6946_/Q _3781_/A2 _5523_/A _7063_/Q _3780_/X VGND VPWR _3782_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5520_ _5520_/A0 hold42/X hold87/A VGND VPWR hold88/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_762 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5451_ hold726/X _5469_/A1 _5453_/S VGND VPWR _5451_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4402_ _4661_/A _4653_/B VGND VPWR _4627_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_5382_ _5382_/A hold17/X VGND VPWR _5390_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_7121_ _7126_/CLK _7121_/D fanout456/X VGND VPWR _7121_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4333_ hold902/X _6357_/A1 _4333_/S VGND VPWR _4333_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7052_ _7086_/CLK _7052_/D fanout482/X VGND VPWR _7052_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4264_ hold267/X _5534_/A1 _4267_/S VGND VPWR _4264_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3215_ _6853_/Q VGND VPWR _3215_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6003_ _6001_/X _6002_/Y _6003_/B1 _6103_/B1 VGND VPWR _7119_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_4195_ _3410_/Y _4195_/A1 _4195_/S VGND VPWR _6598_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_474 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6905_ _7076_/CLK _6905_/D fanout481/X VGND VPWR _6905_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_35_360 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_499 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6836_ _7065_/CLK _6836_/D fanout463/X VGND VPWR _6836_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_10_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6767_ _6890_/CLK _6767_/D fanout470/X VGND VPWR _6767_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3979_ hold20/X hold172/X _6624_/Q VGND VPWR _3979_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5718_ _6821_/Q _5818_/A2 _5642_/X _6965_/Q VGND VPWR _5718_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_164_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_722 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6698_ _6735_/CLK _6698_/D fanout445/X VGND VPWR _6698_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_163_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5649_ _5658_/B _5667_/C VGND VPWR _5652_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_151_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold250 _5402_/X VGND VPWR _6955_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold261 _7072_/Q VGND VPWR hold261/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _5168_/X VGND VPWR _6752_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _6859_/Q VGND VPWR hold283/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _5285_/X VGND VPWR _6851_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_101 _7157_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_112 _7199_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_123 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_134 _6428_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_145 _5513_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_156 hold99/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_167 _3700_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_178 _6301_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_159_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_189 _6423_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_0_csclk clkbuf_0_csclk/X VGND VPWR clkbuf_1_1_1_csclk/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_167_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_732 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput7 mask_rev_in[12] VGND VPWR input7/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_64_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_499 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4951_ _5114_/A _4951_/B VGND VPWR _5047_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_17_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3902_ _4337_/A _4337_/B VGND VPWR _3907_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_4882_ _5023_/D _4882_/B _4882_/C VGND VPWR _4882_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_6621_ _6629_/CLK _6621_/D _6390_/A VGND VPWR _6621_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3833_ _6416_/Q _3838_/A VGND VPWR _3836_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_6552_ _6632_/CLK _6552_/D fanout454/X VGND VPWR _6552_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_146_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3764_ _3763_/X _3764_/A1 _3829_/B VGND VPWR _3764_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_118_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5503_ hold910/X _5548_/A1 hold77/X VGND VPWR _5503_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6483_ _6704_/CLK _6483_/D fanout450/X VGND VPWR _6483_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3695_ _3251_/A _4083_/S _3358_/Y input13/X _3694_/X VGND VPWR _3698_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_161_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput300 _6754_/Q VGND VPWR pwr_ctrl_out[3] VGND VPWR sky130_fd_sc_hd__buf_12
X_5434_ hold521/X hold99/X _5435_/S VGND VPWR _5434_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput311 _7199_/X VGND VPWR spimemio_flash_io2_di VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput322 hold1347/X VGND VPWR hold1348/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput333 hold1349/X VGND VPWR hold1350/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_99_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput344 hold1329/X VGND VPWR hold1330/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_126_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5365_ _5365_/A0 _5524_/A1 _5372_/S VGND VPWR _5365_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_csclk clkbuf_3_3_0_csclk/A VGND VPWR _7001_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_7104_ _7131_/CLK _7104_/D fanout460/X VGND VPWR _7104_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4316_ _4316_/A _6352_/B VGND VPWR _4321_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_5296_ hold916/X _5509_/A1 _5300_/S VGND VPWR _5296_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7035_ _7037_/CLK _7035_/D fanout455/X VGND VPWR _7035_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4247_ hold638/X _5544_/A1 _4249_/S VGND VPWR _4247_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4178_ _6637_/Q _6307_/B VGND VPWR _4186_/S VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_28_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A VGND VPWR clkbuf_3_1_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
X_6819_ _6884_/CLK _6819_/D fanout475/X VGND VPWR _6819_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_50_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_582 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_479 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_702 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_633 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3480_ _7060_/Q hold86/A _5505_/A _7052_/Q VGND VPWR _3480_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5150_ hold890/X _6354_/A1 _5153_/S VGND VPWR _5150_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4101_ hold720/X _4100_/X _4101_/S VGND VPWR _4101_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5081_ _4902_/A _4902_/B _4689_/A _4464_/Y VGND VPWR _5082_/C VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_2_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4032_ _4032_/A _5490_/B VGND VPWR _4037_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_56_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5983_ _6842_/Q _5975_/A _5959_/X _6962_/Q VGND VPWR _5983_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_17_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4934_ _4542_/D _4562_/Y _4620_/Y _4652_/Y _4770_/B VGND VPWR _5003_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_178_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_694 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4865_ _4652_/Y _4700_/Y _4518_/C VGND VPWR _5034_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA_12 _5265_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_32_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_23 _4220_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_34 _3742_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_177_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6604_ _6746_/CLK _6604_/D fanout447/X VGND VPWR _6604_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3816_ _6826_/Q _5256_/A _4244_/A _6645_/Q _3815_/X VGND VPWR _3817_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XANTENNA_45 _5627_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_177_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_56 _5965_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4796_ _4796_/A _5064_/A _4796_/C _4796_/D VGND VPWR _4804_/A VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_67 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_78 _6542_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6535_ _6925_/CLK _6535_/D fanout460/X VGND VPWR _6535_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_89 _6664_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3747_ _7072_/Q _5532_/A _5490_/A _7035_/Q VGND VPWR _3747_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6466_ _6653_/CLK _6466_/D _6401_/A VGND VPWR _6466_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_133_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3678_ _6980_/Q _5427_/A _4238_/A _6632_/Q _3677_/X VGND VPWR _3679_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5417_ hold677/X _5540_/A1 _5417_/S VGND VPWR _5417_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6397_ _6400_/A _6400_/B VGND VPWR _6397_/X VGND VPWR sky130_fd_sc_hd__and2_1
Xoutput174 _3960_/X VGND VPWR irq[2] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5348_ hold572/X _5543_/A1 _5354_/S VGND VPWR _5348_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput185 _3204_/Y VGND VPWR mgmt_gpio_oeb[19] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput196 _3194_/Y VGND VPWR mgmt_gpio_oeb[29] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_87_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5279_ hold467/X _5528_/A1 _5282_/S VGND VPWR _5279_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7018_ _7051_/CLK _7018_/D fanout476/X VGND VPWR _7018_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_56_731 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_614 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_599 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xfanout390 _4372_/X VGND VPWR _4716_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_143_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4650_ _4650_/A _5043_/A VGND VPWR _4650_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xinput10 mask_rev_in[15] VGND VPWR input10/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_3601_ _7050_/Q _5505_/A _5541_/A _7082_/Q VGND VPWR _3601_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xinput21 mask_rev_in[25] VGND VPWR input21/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_190_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput32 mask_rev_in[6] VGND VPWR input32/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _4810_/A _4581_/B VGND VPWR _4581_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xinput43 mgmt_gpio_in[16] VGND VPWR input43/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VPWR input54/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6320_ _6320_/A _6320_/B VGND VPWR _6320_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_155_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput65 mgmt_gpio_in[36] VGND VPWR _7199_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xhold805 _3992_/X VGND VPWR _6435_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ hold85/X _3714_/B VGND VPWR _5148_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xinput76 qspi_enabled VGND VPWR _3921_/S VGND VPWR sky130_fd_sc_hd__clkbuf_8
Xhold816 _7083_/Q VGND VPWR hold816/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VPWR _7198_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VPWR input98/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold827 _4327_/X VGND VPWR _6714_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _6694_/Q VGND VPWR hold838/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold849 _4046_/X VGND VPWR _6481_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ _6243_/X _6251_/B _6301_/C VGND VPWR _6251_/X VGND VPWR sky130_fd_sc_hd__and3b_1
X_3463_ _6431_/Q _3981_/A _3381_/Y input31/X _3462_/X VGND VPWR _3467_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_5202_ _6396_/B _5202_/B _5505_/B VGND VPWR _5210_/S VGND VPWR sky130_fd_sc_hd__and3b_4
X_6182_ _7151_/Q _5958_/X _5978_/X _6480_/Q VGND VPWR _6182_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3394_ input42/X _5202_/B _3999_/A _6449_/Q VGND VPWR _3394_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_111_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5133_ _4628_/Y _4970_/Y _5010_/Y _4631_/Y _4796_/D VGND VPWR _5134_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_96_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1505 _6588_/Q VGND VPWR _4184_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1516 _7105_/Q VGND VPWR _5609_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _7141_/Q VGND VPWR _6325_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1538 hold97/A VGND VPWR _3255_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5064_ _5064_/A _5064_/B _5064_/C VGND VPWR _5106_/C VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1549 _7099_/Q VGND VPWR _5592_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4015_ _4015_/A0 _6353_/A1 _4019_/S VGND VPWR _4015_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_65_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5966_ _5966_/A _5981_/B _5981_/C VGND VPWR _5971_/C VGND VPWR sky130_fd_sc_hd__and3_4
X_4917_ _4359_/Y _4887_/A _4384_/A _4887_/B _4872_/B VGND VPWR _5033_/A VGND VPWR
+ sky130_fd_sc_hd__o41a_1
X_5897_ _6648_/Q _5621_/X _5913_/B1 _6553_/Q VGND VPWR _5897_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_32_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4848_ _4469_/A _4689_/A _4490_/B VGND VPWR _5029_/A VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_165_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4779_ _4902_/B _4611_/Y _4500_/A VGND VPWR _5068_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_107_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6518_ _6755_/CLK _6518_/D _6360_/A VGND VPWR _6518_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_134_555 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6449_ _7070_/CLK _6449_/D fanout473/X VGND VPWR _6449_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_csclk _6888_/CLK VGND VPWR _6951_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xclkbuf_2_0_0_csclk clkbuf_2_1_0_csclk/A VGND VPWR clkbuf_3_1_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_189_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_369 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_255 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_602 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_146 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_588 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5820_ _6507_/Q _5820_/A2 _5611_/Y VGND VPWR _5820_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_34_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5751_ _6950_/Q _5637_/X _5660_/X _6806_/Q VGND VPWR _5751_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_187_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4702_ _4702_/A _4702_/B _4702_/C _4965_/B VGND VPWR _4702_/Y VGND VPWR sky130_fd_sc_hd__nand4_2
XFILLER_148_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5682_ _6867_/Q _5628_/X _5666_/X _6891_/Q VGND VPWR _5682_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4633_ _4631_/D _4633_/B VGND VPWR _4661_/B VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_163_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4564_ _4564_/A _4773_/A VGND VPWR _4566_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_118_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold602 _7040_/Q VGND VPWR hold602/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold613 _4277_/X VGND VPWR _6672_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _7130_/Q _6302_/X _6303_/S VGND VPWR _6303_/X VGND VPWR sky130_fd_sc_hd__mux2_2
Xhold624 _6849_/Q VGND VPWR hold624/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 _5420_/X VGND VPWR _6971_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3515_ _3555_/A _3562_/B VGND VPWR _4214_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold646 _6445_/Q VGND VPWR hold646/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _4495_/A _4632_/B VGND VPWR _5042_/B VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold657 _5469_/X VGND VPWR _7015_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmax_cap376 _5611_/Y VGND VPWR _6103_/B1 VGND VPWR sky130_fd_sc_hd__buf_4
Xhold668 _5174_/X VGND VPWR _6756_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap387 _5631_/X VGND VPWR _5818_/A2 VGND VPWR sky130_fd_sc_hd__buf_8
Xhold679 _6833_/Q VGND VPWR hold679/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6477_/Q _5940_/X _5967_/X _6606_/Q _6231_/X VGND VPWR _6234_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3446_ _3446_/A _3446_/B _3446_/C _3446_/D VGND VPWR _3446_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_170_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6165_ _6165_/A _6165_/B _6165_/C VGND VPWR _6176_/C VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_134_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3377_ _3455_/A hold28/X VGND VPWR _5541_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1302 _3991_/X VGND VPWR _6434_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ _5116_/A VGND VPWR _5116_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_97_483 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1313 _7034_/Q VGND VPWR _5491_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1324 hold1324/A VGND VPWR wb_dat_o[21] VGND VPWR sky130_fd_sc_hd__buf_12
X_6096_ _7030_/Q _5944_/X _5975_/A _6846_/Q _6095_/X VGND VPWR _6099_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_196 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1335 hold1418/X VGND VPWR hold1335/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 hold1346/A VGND VPWR wb_dat_o[14] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_27_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1357 _6310_/A1 VGND VPWR hold1357/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 hold1368/A VGND VPWR wb_dat_o[2] VGND VPWR sky130_fd_sc_hd__buf_12
X_5047_ _5047_/A _5096_/B VGND VPWR _5122_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_84_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1379 hold1557/X VGND VPWR hold1379/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_712 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_406 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6998_ _7065_/CLK _6998_/D fanout465/X VGND VPWR _6998_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5949_ _5978_/A _5981_/A _5981_/B VGND VPWR _5949_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_43_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_483 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_572 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_734 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_726 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_190 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_671 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3300_ _3355_/B _3311_/C VGND VPWR _3300_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
X_4280_ _4280_/A _5490_/B VGND VPWR _4285_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_140_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3231_ _3837_/A _3234_/C VGND VPWR _3829_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_82_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6921_ _7001_/CLK _6921_/D fanout464/X VGND VPWR _6921_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_704 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6852_ _7049_/CLK _6852_/D fanout456/X VGND VPWR _6852_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_50_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5803_ _6993_/Q _5627_/X _5635_/X _6833_/Q VGND VPWR _5803_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6783_ _6890_/CLK _6783_/D fanout476/X VGND VPWR _6783_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3995_ hold586/X _6357_/A1 _3998_/S VGND VPWR _3995_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5734_ _6789_/Q _5652_/Y _5728_/X _5733_/X _3178_/Y VGND VPWR _5734_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5665_ _6858_/Q _5663_/X _5664_/X _6922_/Q VGND VPWR _5665_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_175_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_628 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4616_ _4716_/A _4698_/C VGND VPWR _4616_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
X_5596_ _5596_/A1 _5574_/Y _5597_/B _5595_/X VGND VPWR _7100_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_135_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold410 _5517_/X VGND VPWR _7057_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _6671_/Q VGND VPWR hold421/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _4881_/B _4576_/B VGND VPWR _5114_/A VGND VPWR sky130_fd_sc_hd__nand2_4
Xhold432 _4325_/X VGND VPWR _6712_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 _7193_/A VGND VPWR hold443/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _4148_/X VGND VPWR _6557_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 _6878_/Q VGND VPWR hold465/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _5306_/X VGND VPWR _6870_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4642_/A _4739_/A VGND VPWR _4653_/C VGND VPWR sky130_fd_sc_hd__and2b_4
Xhold487 _6621_/Q VGND VPWR hold487/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _5453_/X VGND VPWR _7001_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6217_ _6461_/Q _5945_/X _5975_/C _6579_/Q _6216_/X VGND VPWR _6218_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3429_ input59/X _5193_/A _3358_/Y input18/X _3418_/X VGND VPWR _3429_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7197_ _7197_/A VGND VPWR _7197_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6148_ _6448_/Q _5601_/X _5959_/X _6968_/Q VGND VPWR _6148_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_58_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1110 _5413_/X VGND VPWR _6965_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 _6717_/Q VGND VPWR _4331_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 _4175_/X VGND VPWR _6580_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1143 _6565_/Q VGND VPWR _4158_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 _5257_/X VGND VPWR _6826_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6079_ _7014_/Q _5940_/X _5967_/X _6854_/Q VGND VPWR _6079_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_45_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1165 hold1576/X VGND VPWR _4110_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1176 _4053_/X VGND VPWR _6490_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _6442_/Q VGND VPWR _4000_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1198 _5326_/X VGND VPWR _6888_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_344 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_464 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_136 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3780_ input93/X _5190_/A _3355_/X _5283_/A _6850_/Q VGND VPWR _3780_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_158_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5450_ hold152/X hold60/X _5453_/S VGND VPWR _5450_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4401_ _4633_/B _4631_/D VGND VPWR _4653_/B VGND VPWR sky130_fd_sc_hd__and2b_4
X_5381_ hold307/X _5540_/A1 _5381_/S VGND VPWR _5381_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A VGND VPWR _7131_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_7120_ _7126_/CLK _7120_/D fanout466/X VGND VPWR _7120_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4332_ hold373/X _5494_/A1 _4333_/S VGND VPWR _4332_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7051_ _7051_/CLK _7051_/D fanout485/X VGND VPWR _7051_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_87_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4263_ _4263_/A0 hold667/X _4267_/S VGND VPWR _4263_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6002_ _6786_/Q _6226_/B _5610_/Y VGND VPWR _6002_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
X_3214_ _6861_/Q VGND VPWR _3214_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4194_ _3447_/Y _4194_/A1 _4195_/S VGND VPWR _6597_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_762 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_486 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6904_ _7069_/CLK _6904_/D fanout482/X VGND VPWR _6904_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6835_ _7063_/CLK _6835_/D fanout463/X VGND VPWR _6835_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_23_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6766_ _6890_/CLK _6766_/D fanout470/X VGND VPWR _6766_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3978_ _3978_/A0 hold99/X _3980_/S VGND VPWR _3978_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5717_ _3207_/Y _5899_/B _5651_/B VGND VPWR _5717_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_109_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6697_ _6755_/CLK _6697_/D fanout445/X VGND VPWR _6697_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_40_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR _3945_/A1 VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_164_734 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5648_ _5664_/A _5658_/B _5663_/C VGND VPWR _5648_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_108_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5579_ _6508_/Q _5658_/B _5667_/C VGND VPWR _5583_/S VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_151_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold240 _4082_/X VGND VPWR _6504_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 _6787_/Q VGND VPWR hold251/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _5534_/X VGND VPWR _7072_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold273 _6620_/Q VGND VPWR hold273/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _5294_/X VGND VPWR _6859_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _6931_/Q VGND VPWR hold295/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_102 _7157_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_113 input64/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_124 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_135 _6431_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_146 _5513_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_157 hold99/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_168 _3700_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_179 _5978_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_556 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput8 mask_rev_in[13] VGND VPWR input8/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_49_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4950_ _4574_/A _4723_/B _4581_/Y _4810_/Y VGND VPWR _4950_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_3901_ _4374_/A _4702_/C _3901_/C _3901_/D VGND VPWR _3907_/A VGND VPWR sky130_fd_sc_hd__and4b_1
X_4881_ _4881_/A _4881_/B VGND VPWR _4882_/C VGND VPWR sky130_fd_sc_hd__nand2_1
X_6620_ _6712_/CLK _6620_/D fanout470/X VGND VPWR _6620_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3832_ _3837_/A _3832_/B VGND VPWR _3838_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_6551_ _6632_/CLK _6551_/D fanout454/X VGND VPWR _6551_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3763_ _3762_/Y _6727_/Q _3829_/A VGND VPWR _3763_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5502_ _5502_/A0 hold42/X hold77/X VGND VPWR hold78/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_6482_ _6707_/CLK _6482_/D fanout450/X VGND VPWR _6482_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3694_ _7057_/Q hold86/A _4232_/A _6627_/Q VGND VPWR _3694_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5433_ hold698/X _5469_/A1 _5435_/S VGND VPWR _5433_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput301 _3788_/Y VGND VPWR reset VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput312 _7200_/X VGND VPWR spimemio_flash_io3_di VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput323 hold1319/X VGND VPWR hold1320/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput334 hold1377/X VGND VPWR hold1378/A VGND VPWR sky130_fd_sc_hd__buf_12
X_5364_ _5364_/A hold17/X VGND VPWR _5372_/S VGND VPWR sky130_fd_sc_hd__and2_4
Xoutput345 hold1341/X VGND VPWR hold1342/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_113_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7103_ _7131_/CLK _7103_/D fanout460/X VGND VPWR _7103_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4315_ hold614/X _6357_/A1 _4315_/S VGND VPWR _4315_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5295_ hold407/X _5544_/A1 _5300_/S VGND VPWR _5295_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7034_ _7037_/CLK _7034_/D fanout450/X VGND VPWR _7034_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4246_ hold415/X _5534_/A1 _4249_/S VGND VPWR _4246_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_710 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4177_ hold562/X _6357_/A1 _4177_/S VGND VPWR _4177_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_364 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6818_ _7067_/CLK _6818_/D fanout476/X VGND VPWR _6818_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_51_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6749_ _6749_/CLK _6749_/D fanout449/X VGND VPWR _6749_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_183_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_714 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_386 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_299 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4100_ hold341/X _5540_/A1 _5202_/B VGND VPWR _4100_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5080_ _5080_/A _5080_/B _5080_/C VGND VPWR _5087_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_150_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4031_ _4031_/A0 hold60/X hold68/X VGND VPWR hold69/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5982_ _6810_/Q _5971_/B _5946_/X _6890_/Q VGND VPWR _5982_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4933_ _5068_/C _5002_/C _4933_/C _5138_/A VGND VPWR _4944_/A VGND VPWR sky130_fd_sc_hd__and4_1
X_4864_ _4618_/Y _4694_/Y _5084_/A VGND VPWR _4864_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA_13 _5265_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_24 _3508_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6603_ _6674_/CLK _6603_/D _6383_/A VGND VPWR _6603_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3815_ _7002_/Q _3370_/Y _5184_/A _6764_/Q VGND VPWR _3815_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XANTENNA_35 _3828_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_46 _5627_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4795_ _4546_/Y _4631_/Y _4697_/Y VGND VPWR _4796_/D VGND VPWR sky130_fd_sc_hd__o21a_1
XANTENNA_57 _5971_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_192_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_68 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6534_ _6539_/CLK _6534_/D fanout461/X VGND VPWR _6534_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_79 _6787_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_118_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3746_ _6762_/Q _5182_/S _4304_/A _6696_/Q _3745_/X VGND VPWR _3751_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6465_ _6654_/CLK _6465_/D _6401_/A VGND VPWR _6465_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3677_ _7028_/Q hold49/A _5505_/A _7049_/Q VGND VPWR _3677_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_173_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5416_ hold924/X _5548_/A1 _5417_/S VGND VPWR _5416_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6396_ _6396_/A _6396_/B VGND VPWR _6396_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5347_ _5347_/A0 _5473_/A1 _5354_/S VGND VPWR _5347_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_770 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput175 _3935_/X VGND VPWR mgmt_gpio_oeb[0] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput186 _3934_/X VGND VPWR mgmt_gpio_oeb[1] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_623 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput197 _3220_/Y VGND VPWR mgmt_gpio_oeb[2] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5278_ hold914/X _5509_/A1 _5282_/S VGND VPWR _5278_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7017_ _7017_/CLK _7017_/D fanout461/X VGND VPWR _7017_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4229_ _6640_/Q _4230_/B VGND VPWR _4229_/X VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_56_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_475 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3600_ _6893_/Q _5328_/A _5166_/A _6754_/Q _3591_/X VGND VPWR _3604_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xinput11 mask_rev_in[16] VGND VPWR input11/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 mask_rev_in[26] VGND VPWR input22/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4580_ _4561_/B _4611_/B _4948_/D _4578_/X _4575_/Y VGND VPWR _4580_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
Xinput33 mask_rev_in[7] VGND VPWR input33/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput44 mgmt_gpio_in[17] VGND VPWR input44/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput55 mgmt_gpio_in[27] VGND VPWR input55/X VGND VPWR sky130_fd_sc_hd__buf_2
X_3531_ _6564_/Q _4151_/A _4262_/A _6664_/Q VGND VPWR _3531_/X VGND VPWR sky130_fd_sc_hd__a22o_2
Xinput66 mgmt_gpio_in[37] VGND VPWR _7200_/A VGND VPWR sky130_fd_sc_hd__buf_4
Xinput77 ser_tx VGND VPWR input77/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xhold806 _7075_/Q VGND VPWR hold806/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _5546_/X VGND VPWR _7083_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VPWR _3949_/B VGND VPWR sky130_fd_sc_hd__buf_4
Xhold828 _6427_/Q VGND VPWR hold828/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wb_adr_i[0] VGND VPWR _4563_/A VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold839 _4303_/X VGND VPWR _6694_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6250_ _6250_/A _6250_/B _6250_/C _6250_/D VGND VPWR _6251_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_115_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3462_ _6975_/Q _5418_/A _5373_/A _6935_/Q VGND VPWR _3462_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_5201_ hold395/X _5540_/A1 _5201_/S VGND VPWR _5201_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_131_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6181_ _6609_/Q _5943_/X _5981_/X _6655_/Q VGND VPWR _6181_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3393_ _6953_/Q _3781_/A2 _3358_/Y input19/X _3383_/X VGND VPWR _3393_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5132_ _5087_/A _5120_/X _5131_/X _5116_/Y VGND VPWR _5143_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_123_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_367 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1506 _7131_/Q VGND VPWR _6304_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1517 _7128_/Q VGND VPWR _6229_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5063_ _4619_/Y _5010_/Y _4974_/B VGND VPWR _5064_/C VGND VPWR sky130_fd_sc_hd__o21a_1
Xhold1528 _7161_/Q VGND VPWR _3259_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _7150_/Q VGND VPWR _6351_/A2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4014_ _4014_/A _6352_/B VGND VPWR _4019_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_65_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5965_ _5979_/A _5981_/B _5969_/C VGND VPWR _5965_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_12_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4916_ _5118_/A _4916_/B _4916_/C VGND VPWR _4918_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_5896_ _5896_/A _5896_/B _5896_/C VGND VPWR _5896_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_4847_ _4847_/A VGND VPWR _4847_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4778_ _5023_/B _5039_/B _4777_/X _4593_/Y VGND VPWR _4884_/B VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_165_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6517_ _7076_/CLK _6517_/D fanout481/X VGND VPWR _6517_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3729_ _3729_/A _3729_/B _3729_/C _3729_/D VGND VPWR _3730_/C VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_146_372 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6448_ _7086_/CLK _6448_/D fanout483/X VGND VPWR _6448_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_134_567 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6379_ _6401_/A _6401_/B VGND VPWR _6379_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5750_ _6838_/Q _5928_/A2 _5740_/X _5749_/X VGND VPWR _5754_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_4701_ _4702_/A _4702_/B _4702_/C VGND VPWR _4701_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
X_5681_ _5681_/A _5681_/B _5681_/C VGND VPWR _5681_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_4632_ _4753_/B _4632_/B VGND VPWR _4632_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_163_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4563_ _4563_/A _4631_/D _4633_/B _4563_/D VGND VPWR _4773_/A VGND VPWR sky130_fd_sc_hd__and4_1
Xhold603 _5498_/X VGND VPWR _7040_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold614 _6704_/Q VGND VPWR hold614/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ _6289_/Y _6301_/X _6544_/Q _6226_/B VGND VPWR _6302_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3514_ _6649_/Q _4244_/A _3511_/Y _3513_/X _3414_/Y VGND VPWR _3523_/B VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_116_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold625 _5282_/X VGND VPWR _6849_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _6952_/Q VGND VPWR hold636/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _5010_/A _4881_/B VGND VPWR _4494_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold647 _4003_/X VGND VPWR _6445_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _6945_/Q VGND VPWR hold658/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ _6692_/Q _5954_/X _5976_/D _6621_/Q _6230_/X VGND VPWR _6250_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xmax_cap377 hold74/X VGND VPWR hold75/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold669 _6864_/Q VGND VPWR hold669/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3445_ _6968_/Q _5409_/A _3365_/Y input9/X _3444_/X VGND VPWR _3446_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xmax_cap388 _5616_/X VGND VPWR _5902_/A2 VGND VPWR sky130_fd_sc_hd__buf_8
X_6164_ _6985_/Q _5945_/X _5975_/C _6841_/Q _6157_/X VGND VPWR _6165_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3376_ _3717_/B _3376_/B VGND VPWR _3964_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_85_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5115_ _5115_/A _5115_/B _5115_/C _5115_/D VGND VPWR _5116_/A VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1303 _6540_/Q VGND VPWR _4128_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1314 _5491_/X VGND VPWR _7034_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6095_ _7022_/Q _5937_/X _5975_/D _6886_/Q VGND VPWR _6095_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_97_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1325 hold1422/X VGND VPWR hold1325/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1336 hold1336/A VGND VPWR wb_dat_o[6] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1347 hold1429/X VGND VPWR hold1347/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _5046_/A _5046_/B _5046_/C VGND VPWR _5096_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_27_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1358 hold1358/A VGND VPWR wb_dat_o[26] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1369 _4191_/A1 VGND VPWR hold1369/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6997_ _6997_/CLK _6997_/D fanout465/X VGND VPWR _6997_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_13_418 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5948_ _5969_/A _5981_/A _5981_/C VGND VPWR _5948_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_138_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5879_ _6452_/Q _5634_/X _5876_/X _5878_/X VGND VPWR _5879_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_126_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_746 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_444 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_215 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_738 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3230_ _6417_/Q _6416_/Q VGND VPWR _3234_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_140_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_318 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6920_ _6920_/CLK _6920_/D fanout473/X VGND VPWR _6920_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_6851_ _6963_/CLK _6851_/D fanout456/X VGND VPWR _6851_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5802_ _3228_/Y _5899_/B _5651_/B VGND VPWR _5802_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
X_6782_ _6969_/CLK _6782_/D fanout481/X VGND VPWR _6782_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3994_ hold772/X _6356_/A1 _3998_/S VGND VPWR _3994_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5733_ _6805_/Q _5660_/X _5729_/X _5731_/X _5732_/X VGND VPWR _5733_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
XFILLER_50_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5664_ _5664_/A _5667_/C _5666_/C VGND VPWR _5664_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4615_ _4661_/A _4615_/B VGND VPWR _4615_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_5595_ _6508_/Q _5969_/A _5968_/A VGND VPWR _5595_/X VGND VPWR sky130_fd_sc_hd__and3_1
Xhold400 _5385_/X VGND VPWR _6940_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 _7076_/Q VGND VPWR hold411/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4562_/A _4753_/B VGND VPWR _4546_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold422 _4276_/X VGND VPWR _6671_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold433 _6522_/Q VGND VPWR hold433/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _5198_/X VGND VPWR _6774_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _7022_/Q VGND VPWR hold455/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _5315_/X VGND VPWR _6878_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _5010_/A _4650_/A VGND VPWR _5088_/A VGND VPWR sky130_fd_sc_hd__nand2_4
Xhold477 _6934_/Q VGND VPWR hold477/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold488 _4223_/X VGND VPWR _6621_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _6658_/Q VGND VPWR hold499/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk _7001_/CLK VGND VPWR _7026_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6216_ _6666_/Q _5938_/X _5952_/X _6706_/Q VGND VPWR _6216_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3428_ _6928_/Q _5364_/A _3981_/A _6432_/Q _3427_/X VGND VPWR _3428_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7196_ _7196_/A VGND VPWR _7196_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6147_ _7032_/Q _5944_/X _5975_/A _6848_/Q _6146_/X VGND VPWR _6150_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1100 _5230_/X VGND VPWR _6802_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3359_ _3562_/A hold28/X VGND VPWR _5256_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1111 _6677_/Q VGND VPWR _4283_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 _4331_/X VGND VPWR _6717_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _6818_/Q VGND VPWR _5248_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 _4158_/X VGND VPWR _6565_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ _6078_/A0 _6077_/X _6279_/S VGND VPWR _6078_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1155 _6670_/Q VGND VPWR _4275_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _4110_/X VGND VPWR _6524_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1177 _6665_/Q VGND VPWR _4269_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _5029_/A _5029_/B VGND VPWR _5083_/C VGND VPWR sky130_fd_sc_hd__and2_1
Xhold1188 _4000_/X VGND VPWR _6442_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 _6962_/Q VGND VPWR _5410_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_532 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4400_ _4631_/D _4400_/B VGND VPWR _4408_/B VGND VPWR sky130_fd_sc_hd__xnor2_2
XFILLER_145_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5380_ hold930/X _5548_/A1 _5381_/S VGND VPWR _5380_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4331_ _4331_/A0 _5493_/A1 _4333_/S VGND VPWR _4331_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7050_ _7086_/CLK _7050_/D fanout483/X VGND VPWR _7050_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A _4322_/B VGND VPWR _4267_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_140_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6001_ _5992_/X _6226_/B _6001_/C _6001_/D VGND VPWR _6001_/X VGND VPWR sky130_fd_sc_hd__and4b_1
X_3213_ _6869_/Q VGND VPWR _3213_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4193_ _3486_/Y _4193_/A1 _4195_/S VGND VPWR _6596_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6903_ _7076_/CLK _6903_/D fanout481/X VGND VPWR _6903_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6834_ _7026_/CLK _6834_/D fanout463/X VGND VPWR _6834_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_62_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6765_ _6890_/CLK _6765_/D fanout470/X VGND VPWR _6765_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3977_ hold97/X hold106/X _6624_/Q VGND VPWR _3977_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_149_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5716_ _6445_/Q _5614_/X _5666_/X _6893_/Q VGND VPWR _5716_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_148_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6696_ _6755_/CLK _6696_/D _6360_/A VGND VPWR _6696_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_109_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5647_ _7026_/Q _5645_/X _5646_/X _6906_/Q _5644_/X VGND VPWR _5669_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_16 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_757 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5578_ _7095_/Q _7094_/Q VGND VPWR _5667_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_151_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold230 _4285_/X VGND VPWR _6679_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _6925_/Q VGND VPWR hold241/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _5213_/X VGND VPWR _6787_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4413_/Y _4724_/A VGND VPWR _4529_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_6_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold263 _6443_/Q VGND VPWR hold263/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _4222_/X VGND VPWR _6620_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold285 _6827_/Q VGND VPWR hold285/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _5375_/X VGND VPWR _6931_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7179_ _7179_/A VGND VPWR _7179_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_105_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_103 _7173_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_114 _3957_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_125 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 _6432_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_147 _6357_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_158 hold99/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_169 _3803_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_41_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput9 mask_rev_in[14] VGND VPWR input9/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_52_619 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3900_ input118/X input119/X _3900_/C _3900_/D VGND VPWR _3901_/D VGND VPWR sky130_fd_sc_hd__and4bb_1
XFILLER_32_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4880_ _4951_/B _5086_/B _5073_/A _4880_/D VGND VPWR _4882_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_177_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3831_ _3837_/B _3837_/C VGND VPWR _3832_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_177_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6550_ _6654_/CLK _6550_/D fanout454/X VGND VPWR _6550_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3762_ _3762_/A _3762_/B VGND VPWR _3762_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_5501_ hold182/X _5519_/A1 hold77/A VGND VPWR _5501_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6481_ _6704_/CLK _6481_/D fanout450/X VGND VPWR _6481_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3693_ _6542_/Q _4127_/A _3692_/Y _6765_/Q _3691_/X VGND VPWR _3698_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5432_ hold147/X hold60/X _5435_/S VGND VPWR _5432_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_133_418 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput302 _3956_/X VGND VPWR ser_rx VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput313 hold1379/X VGND VPWR wb_ack_o VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_610 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput324 hold1321/X VGND VPWR hold1322/A VGND VPWR sky130_fd_sc_hd__buf_12
X_5363_ hold489/X hold22/X _5363_/S VGND VPWR _5363_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput335 hold1361/X VGND VPWR hold1362/A VGND VPWR sky130_fd_sc_hd__buf_12
X_7102_ _7113_/CLK _7102_/D fanout464/X VGND VPWR _7102_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4314_ hold782/X _6356_/A1 _4315_/S VGND VPWR _4314_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5294_ hold283/X _5465_/A1 _5300_/S VGND VPWR _5294_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_376 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7033_ _7033_/CLK _7033_/D fanout464/X VGND VPWR _7033_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4245_ _4245_/A0 hold667/X _4249_/S VGND VPWR _4245_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4176_ hold734/X _6356_/A1 _4177_/S VGND VPWR _4176_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_287 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6817_ _7070_/CLK _6817_/D fanout473/X VGND VPWR _6817_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_50_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_540 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6748_ _6926_/CLK _6748_/D fanout449/X VGND VPWR _6748_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_137_702 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6679_ _7036_/CLK _6679_/D fanout455/X VGND VPWR _6679_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_151_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xmgmt_gpio_14_buff_inst _3937_/X VGND VPWR mgmt_gpio_out[14] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_73_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_746 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4030_ _4030_/A0 _5494_/A1 hold68/X VGND VPWR _4030_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5981_ _5981_/A _5981_/B _5981_/C VGND VPWR _5981_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_64_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4932_ _4542_/A _4562_/Y _4673_/A _4628_/Y _4755_/X VGND VPWR _5138_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4542_/B _4496_/Y _4618_/Y _4700_/Y VGND VPWR _4877_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_14 _5505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6602_ _6769_/CLK _6602_/D fanout469/X VGND VPWR _6602_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_25 _4202_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_178_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3814_ _3814_/A _3814_/B VGND VPWR _5184_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XANTENNA_36 _4084_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4794_ _4846_/B _4616_/Y _4619_/Y _4689_/A VGND VPWR _4796_/C VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_47 _5631_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_58 _6301_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_177_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_69 _6075_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6533_ _6755_/CLK _6533_/D _6360_/A VGND VPWR _6533_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3745_ _6859_/Q _5292_/A _3370_/Y _7003_/Q VGND VPWR _3745_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_146_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6464_ _6668_/CLK _6464_/D _6360_/A VGND VPWR _6464_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3676_ _6900_/Q _5337_/A _5301_/A _6868_/Q _3675_/X VGND VPWR _3679_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5415_ hold469/X _5469_/A1 _5417_/S VGND VPWR _5415_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6395_ _6396_/A _6396_/B VGND VPWR _6395_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_114_451 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5346_ _5346_/A _5541_/B VGND VPWR _5354_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput176 _3213_/Y VGND VPWR mgmt_gpio_oeb[10] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput187 _3203_/Y VGND VPWR mgmt_gpio_oeb[20] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput198 _3193_/Y VGND VPWR mgmt_gpio_oeb[30] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_102_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5277_ _5277_/A0 _5484_/A1 _5282_/S VGND VPWR _5277_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7016_ _7016_/CLK _7016_/D fanout474/X VGND VPWR _7016_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4228_ _6638_/Q _4228_/B VGND VPWR _4228_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
XFILLER_46_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4159_ hold810/X _6354_/A1 _4162_/S VGND VPWR _4159_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_73 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout392 hold22/X VGND VPWR _5513_/A1 VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_46_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput12 mask_rev_in[17] VGND VPWR input12/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput23 mask_rev_in[27] VGND VPWR input23/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput34 mask_rev_in[8] VGND VPWR input34/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VPWR input45/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_3530_ hold36/X hold66/X VGND VPWR _4262_/A VGND VPWR sky130_fd_sc_hd__nor2_8
Xinput56 mgmt_gpio_in[28] VGND VPWR input56/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput67 mgmt_gpio_in[3] VGND VPWR _3268_/C VGND VPWR sky130_fd_sc_hd__buf_6
Xhold807 _5537_/X VGND VPWR _7075_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput78 spi_csb VGND VPWR input78/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
Xinput89 spimemio_flash_io2_do VGND VPWR input89/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xhold818 _6696_/Q VGND VPWR hold818/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold829 _3983_/X VGND VPWR _6427_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ _6967_/Q _5409_/A _3964_/A _6423_/Q _3456_/X VGND VPWR _3467_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5200_ hold365/X _5521_/A1 _5201_/S VGND VPWR _5200_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6180_ _6660_/Q _5976_/B _5971_/C _6710_/Q VGND VPWR _6180_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3392_ _3392_/A _3392_/B _3392_/C _3392_/D VGND VPWR _3392_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_69_302 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5131_ _5131_/A _5131_/B _5131_/C VGND VPWR _5131_/X VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1507 _7108_/Q VGND VPWR _5735_/A2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _5062_/A _5062_/B _5062_/C _5062_/D VGND VPWR _5134_/B VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1518 _7111_/Q VGND VPWR _5778_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _3258_/X VGND VPWR _7162_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ hold978/X _5546_/A1 _4013_/S VGND VPWR _4013_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_338 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5964_ _5964_/A _5969_/C _5981_/C VGND VPWR _5975_/D VGND VPWR sky130_fd_sc_hd__and3_4
X_4915_ _4906_/Y _4915_/B _4915_/C _4915_/D VGND VPWR _4916_/C VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_178_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5895_ _6688_/Q _5632_/X _5892_/X _5894_/X VGND VPWR _5896_/C VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_20_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4846_ _4846_/A _4846_/B VGND VPWR _4847_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_166_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4777_ _4753_/A _4602_/Y _5114_/B _4776_/X VGND VPWR _4777_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_6516_ _7076_/CLK _6516_/D fanout481/X VGND VPWR _6516_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_107_716 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3728_ _6939_/Q _5382_/A _4196_/A _6600_/Q _3727_/X VGND VPWR _3729_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_180_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_395 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6447_ _6447_/CLK _6447_/D fanout461/X VGND VPWR _6447_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_106_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3659_ _6908_/Q _5346_/A _5355_/A _6916_/Q VGND VPWR _3659_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_134_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6378_ _6400_/A _6400_/B VGND VPWR _6378_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_0_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5329_ _5329_/A0 _5473_/A1 _5336_/S VGND VPWR _5329_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_307 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_703 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4700_ _4716_/A _4911_/B VGND VPWR _4700_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_5680_ _7019_/Q _5619_/X _5677_/X _5679_/X VGND VPWR _5681_/C VGND VPWR sky130_fd_sc_hd__a211o_2
XFILLER_148_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4633_/B _4716_/A _4653_/C _4631_/D VGND VPWR _4631_/Y VGND VPWR sky130_fd_sc_hd__nand4b_4
XFILLER_8_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4562_ _4562_/A _4600_/B VGND VPWR _4562_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold604 _6811_/Q VGND VPWR hold604/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6301_ _6292_/X _6301_/B _6301_/C VGND VPWR _6301_/X VGND VPWR sky130_fd_sc_hd__and3b_1
Xhold615 _4315_/X VGND VPWR _6704_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ _7067_/Q _5523_/A _4020_/A _6464_/Q VGND VPWR _3513_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_143_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold626 _7017_/Q VGND VPWR hold626/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4493_ _5010_/A _4493_/B VGND VPWR _5083_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold637 _5398_/X VGND VPWR _6952_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _7007_/Q VGND VPWR hold648/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold659 _5390_/X VGND VPWR _6945_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _7153_/Q _5958_/X _5978_/X _6482_/Q VGND VPWR _6232_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xmax_cap378 _3543_/A VGND VPWR _3573_/A VGND VPWR sky130_fd_sc_hd__buf_12
X_3444_ _6952_/Q _5391_/A hold29/A _7024_/Q VGND VPWR _3444_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_103_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_696 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6163_ _6977_/Q _5947_/X _5965_/X _6801_/Q _6162_/X VGND VPWR _6165_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3375_ _3375_/A _3415_/B VGND VPWR _3814_/B VGND VPWR sky130_fd_sc_hd__nand2_8
X_5114_ _5114_/A _5114_/B _5114_/C _5114_/D VGND VPWR _5115_/D VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1304 _4128_/X VGND VPWR _6540_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6094_ _7067_/Q _5934_/X _5975_/B _6870_/Q _6093_/X VGND VPWR _6094_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_84_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1315 hold1412/X VGND VPWR hold1315/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1326 hold1326/A VGND VPWR wb_dat_o[10] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1337 hold1421/X VGND VPWR hold1337/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1348 hold1348/A VGND VPWR wb_dat_o[17] VGND VPWR sky130_fd_sc_hd__buf_12
X_5045_ _4947_/B _4453_/B _4570_/Y VGND VPWR _5046_/C VGND VPWR sky130_fd_sc_hd__a21o_1
Xhold1359 _4168_/A1 VGND VPWR hold1359/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6996_ _7063_/CLK _6996_/D fanout463/X VGND VPWR _6996_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_43_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5947_ _5969_/A _5968_/A _5981_/A VGND VPWR _5947_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_178_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5878_ _6647_/Q _5621_/X _5648_/X _6606_/Q _5877_/X VGND VPWR _5878_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4829_ _4456_/Y _4810_/B _4818_/X _4820_/X VGND VPWR _4829_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_138_148 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_758 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_402 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_227 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VPWR hold1/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_444 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6850_ _6926_/CLK _6850_/D fanout457/X VGND VPWR _6850_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5801_ _6905_/Q _5621_/X _5648_/X _6857_/Q VGND VPWR _5801_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6781_ _6969_/CLK _6781_/D fanout473/X VGND VPWR _6781_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3993_ hold984/X _6355_/A1 _3998_/S VGND VPWR _3993_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5732_ _6925_/Q _5664_/X _5716_/X _5718_/X VGND VPWR _5732_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_5663_ _5664_/A _5666_/C _5663_/C VGND VPWR _5663_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_163_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4614_ _4661_/A _4615_/B VGND VPWR _4698_/C VGND VPWR sky130_fd_sc_hd__and2_2
X_5594_ _5594_/A _5964_/A VGND VPWR _5597_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_191_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold401 _6534_/Q VGND VPWR hold401/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4545_ _4562_/A _4753_/B VGND VPWR _4576_/B VGND VPWR sky130_fd_sc_hd__and2_2
Xhold412 _5538_/X VGND VPWR _7076_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _6769_/Q VGND VPWR hold423/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _4107_/X VGND VPWR _6522_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold445 _6950_/Q VGND VPWR hold445/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold456 _5477_/X VGND VPWR _7022_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _4984_/A _4710_/A VGND VPWR _4476_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold467 _6846_/Q VGND VPWR hold467/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 _5378_/X VGND VPWR _6934_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _6921_/Q VGND VPWR hold489/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6451_/Q _5947_/X _5965_/X _6546_/Q _6214_/X VGND VPWR _6218_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3427_ input69/X _4083_/S _5532_/A _7077_/Q VGND VPWR _3427_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7195_ _7195_/A VGND VPWR _7195_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6146_ _7024_/Q _5937_/X _5975_/D _6888_/Q VGND VPWR _6146_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3358_ _3511_/A _3573_/B VGND VPWR _3358_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
Xhold1101 _6869_/Q VGND VPWR _5305_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1112 _4283_/X VGND VPWR _6677_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1123 _6632_/Q VGND VPWR _4241_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1134 _5248_/X VGND VPWR _6818_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ _7121_/Q _6076_/X _6303_/S VGND VPWR _6077_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1145 _6512_/Q VGND VPWR _4091_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3289_ hold32/X _6488_/Q _3288_/Y VGND VPWR hold33/A VGND VPWR sky130_fd_sc_hd__a21bo_1
Xhold1156 _4275_/X VGND VPWR _6670_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _6550_/Q VGND VPWR _4140_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1178 _4269_/X VGND VPWR _6665_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ _4623_/Y _4695_/Y _4875_/A _4522_/D VGND VPWR _5085_/B VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_38_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1189 _7151_/Q VGND VPWR _6353_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_110_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6979_ _7063_/CLK _6979_/D fanout463/X VGND VPWR _6979_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_80_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_435 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold990 _6763_/Q VGND VPWR hold990/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_544 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_600 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4330_ _4330_/A0 _5492_/A1 _4333_/S VGND VPWR _4330_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_153_482 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_633 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4261_ hold970/X _5546_/A1 _4261_/S VGND VPWR _4261_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6000_ _6000_/A _6000_/B _6000_/C _6000_/D VGND VPWR _6001_/D VGND VPWR sky130_fd_sc_hd__nor4_1
X_3212_ _6877_/Q VGND VPWR _3212_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_140_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4192_ _4192_/A0 _4192_/A1 _4195_/S VGND VPWR _6595_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6902_ _7079_/CLK _6902_/D fanout478/X VGND VPWR _6902_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6833_ _6969_/CLK _6833_/D fanout473/X VGND VPWR _6833_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_24_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6764_ _6926_/CLK _6764_/D fanout457/X VGND VPWR _6764_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3976_ hold689/X _5469_/A1 _3980_/S VGND VPWR _3976_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5715_ _6845_/Q _5902_/A2 _5928_/A2 _6837_/Q VGND VPWR _5715_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6695_ _6735_/CLK _6695_/D fanout445/X VGND VPWR _6695_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_191_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5646_ _5664_/A _5667_/B _5666_/B VGND VPWR _5646_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_164_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5577_ _7094_/Q _5576_/B _5574_/Y _5576_/Y VGND VPWR _7094_/D VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold220 _5449_/X VGND VPWR _6997_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold231 _6981_/Q VGND VPWR hold231/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _4542_/B _4947_/B _4902_/A _4413_/Y _4527_/X VGND VPWR _4528_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold242 _5368_/X VGND VPWR _6925_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _7003_/Q VGND VPWR hold253/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _4001_/X VGND VPWR _6443_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold275 _7011_/Q VGND VPWR hold275/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _5258_/X VGND VPWR _6827_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4459_/A _4459_/B VGND VPWR _4542_/D VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_104_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold297 _6835_/Q VGND VPWR hold297/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7178_ _7178_/A VGND VPWR _7178_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_131_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_390 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6129_ _6129_/A0 _6128_/X _6304_/S VGND VPWR _7124_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_104 user_clock VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_61_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_115 _3251_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_126 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_137 _6433_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_148 _5528_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_159 hold666/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_81_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_674 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_327 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_712 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3830_ _3830_/A1 _3829_/B _3828_/Y _3829_/Y VGND VPWR _6727_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_189_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_68_csclk _7001_/CLK VGND VPWR _7063_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_32_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3761_ _3733_/X _3761_/B _3761_/C _3761_/D VGND VPWR _3762_/B VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_13_591 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5500_ hold590/X _5509_/A1 hold77/X VGND VPWR _5500_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6480_ _6707_/CLK _6480_/D fanout450/X VGND VPWR _6480_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3692_ _3692_/A _3714_/B VGND VPWR _3692_/Y VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_145_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5431_ hold231/X _5494_/A1 _5435_/S VGND VPWR _5431_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_173_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput303 _5606_/A VGND VPWR serial_clock VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput314 hold1371/X VGND VPWR hold1372/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_161_739 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5362_ hold718/X _5521_/A1 _5363_/S VGND VPWR _5362_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput325 hold1365/X VGND VPWR hold1366/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput336 hold1367/X VGND VPWR hold1368/A VGND VPWR sky130_fd_sc_hd__buf_12
X_7101_ _7113_/CLK _7101_/D fanout464/X VGND VPWR _7101_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4313_ hold972/X _6355_/A1 _4315_/S VGND VPWR _4313_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_666 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5293_ _5293_/A0 _6353_/A1 _5300_/S VGND VPWR _5293_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7032_ _7086_/CLK _7032_/D fanout483/X VGND VPWR _7032_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4244_ _4244_/A _4322_/B VGND VPWR _4249_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_141_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4175_ _4175_/A0 _6355_/A1 _4177_/S VGND VPWR _4175_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_406 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_480 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6816_ _7069_/CLK _6816_/D fanout482/X VGND VPWR _6816_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_11_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6747_ _6747_/CLK _6747_/D fanout447/X VGND VPWR _6747_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3959_ _6768_/Q _3959_/B VGND VPWR _3959_/X VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_149_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6678_ _7037_/CLK _6678_/D fanout455/X VGND VPWR _6678_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_164_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5629_ _6986_/Q _5627_/X _5628_/X _6866_/Q _5626_/X VGND VPWR _5641_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_151_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_496 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_620 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_322 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_576 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_539 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5980_ _6850_/Q _5967_/X _5979_/X _6986_/Q VGND VPWR _5980_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_52_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_428 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4931_ _4741_/A _4741_/B _4921_/Y _4612_/Y _4663_/Y VGND VPWR _4933_/C VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_33_642 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4862_ _4456_/Y _4496_/Y _4689_/Y VGND VPWR _4872_/B VGND VPWR sky130_fd_sc_hd__o21ba_1
XFILLER_177_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6601_ _6601_/CLK _6601_/D fanout469/X VGND VPWR _6601_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_177_135 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3813_ _6858_/Q _5292_/A _5328_/A _6890_/Q _3812_/X VGND VPWR _3817_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XANTENNA_15 _5505_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_26 _4127_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4793_ _4846_/B _4619_/Y _4645_/Y _4689_/A VGND VPWR _5064_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XANTENNA_37 _4108_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_20_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_48 _5637_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_119_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6532_ _6735_/CLK _6532_/D _3946_/B VGND VPWR _6532_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XANTENNA_59 _6301_/C VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3744_ _6743_/Q _5154_/A _4214_/A _6615_/Q _3743_/X VGND VPWR _3751_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6463_ _6668_/CLK _6463_/D _6400_/A VGND VPWR _6463_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3675_ _6924_/Q _5364_/A _4316_/A _6707_/Q VGND VPWR _3675_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_173_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5414_ hold802/X _5546_/A1 _5417_/S VGND VPWR _5414_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6394_ _6396_/A _6396_/B VGND VPWR _6394_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_161_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5345_ hold331/X _5540_/A1 _5345_/S VGND VPWR _5345_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_463 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput177 _3212_/Y VGND VPWR mgmt_gpio_oeb[11] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput188 _3202_/Y VGND VPWR mgmt_gpio_oeb[21] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput199 _3192_/Y VGND VPWR mgmt_gpio_oeb[31] VGND VPWR sky130_fd_sc_hd__buf_12
X_5276_ hold560/X _5543_/A1 _5282_/S VGND VPWR _5276_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7015_ _7017_/CLK _7015_/D fanout461/X VGND VPWR _7015_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_102_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4227_ _6636_/Q _6637_/Q _6639_/Q VGND VPWR _4228_/B VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_56_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4158_ _4158_/A0 _5491_/A1 _4162_/S VGND VPWR _4158_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_43_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4089_ hold610/X _4088_/X _4101_/S VGND VPWR _4089_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_192_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout393 hold22/X VGND VPWR _5540_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_46_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput13 mask_rev_in[18] VGND VPWR input13/X VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_128_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput24 mask_rev_in[28] VGND VPWR input24/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput35 mask_rev_in[9] VGND VPWR input35/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput46 mgmt_gpio_in[19] VGND VPWR input46/X VGND VPWR sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VPWR input57/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VPWR _3956_/A VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xhold808 _6541_/Q VGND VPWR hold808/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 spi_enabled VGND VPWR _3957_/B VGND VPWR sky130_fd_sc_hd__clkbuf_4
Xhold819 _4306_/X VGND VPWR _6696_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3460_ input49/X _4058_/S _5523_/A _7068_/Q VGND VPWR _3460_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3391_ _6921_/Q _5355_/A _5274_/A _6849_/Q _3390_/X VGND VPWR _3392_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_314 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5130_ _4691_/A _4631_/Y _4855_/Y _4895_/B _4518_/B VGND VPWR _5131_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_123_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1508 _6586_/Q VGND VPWR _4182_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _5061_/A1 _4229_/X _5022_/Y _5060_/X VGND VPWR _6723_/D VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_96_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1519 _5778_/X VGND VPWR _7111_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ hold507/X _5518_/A1 _4013_/S VGND VPWR _4012_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5963_ _5978_/A _5969_/A _5969_/C VGND VPWR _5975_/C VGND VPWR sky130_fd_sc_hd__and3_4
Xclkbuf_opt_4_0_csclk _6888_/CLK VGND VPWR clkbuf_opt_4_0_csclk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_52_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4914_ _5114_/B _5083_/B _5114_/C VGND VPWR _4915_/D VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_80_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5894_ _6568_/Q _5635_/X _5654_/X _6678_/Q _5893_/X VGND VPWR _5894_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4845_ _4907_/B _5042_/B _4644_/B _4911_/B VGND VPWR _4845_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_32_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4776_ _5088_/A _5114_/A _4776_/C VGND VPWR _4776_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_165_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6515_ _6890_/CLK _6515_/D fanout476/X VGND VPWR _6515_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3727_ _7040_/Q hold76/A _6352_/A _7152_/Q VGND VPWR _3727_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_174_672 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6446_ _7081_/CLK hold80/X fanout478/X VGND VPWR hold79/A VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3658_ _6796_/Q _3326_/Y _5154_/A _6744_/Q _3657_/X VGND VPWR _3661_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_161_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6377_ _6400_/A _6400_/B VGND VPWR _6377_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3589_ _7058_/Q hold86/A _4274_/A _6673_/Q VGND VPWR _3589_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_88_623 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5328_ _5328_/A _5541_/B VGND VPWR _5336_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5259_ hold844/X _5484_/A1 _5264_/S VGND VPWR _5259_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_564 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_575 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4630_ _4633_/B _4716_/A _4653_/C _4631_/D VGND VPWR _4630_/X VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_8_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4561_ _4690_/A _4561_/B VGND VPWR _5043_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_190_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6300_ _6300_/A _6300_/B _6300_/C _6300_/D VGND VPWR _6301_/B VGND VPWR sky130_fd_sc_hd__nor4_1
X_3512_ _3546_/A _3573_/A VGND VPWR _4020_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold605 _5240_/X VGND VPWR _6811_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 _6459_/Q VGND VPWR hold616/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _4739_/A _4911_/A _4896_/A _4492_/D VGND VPWR _4881_/B VGND VPWR sky130_fd_sc_hd__and4b_4
Xhold627 _5471_/X VGND VPWR _7017_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _6647_/Q VGND VPWR hold638/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 _5460_/X VGND VPWR _7007_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _6611_/Q _5943_/X _5981_/X _6657_/Q VGND VPWR _6231_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_143_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3443_ input41/X _5202_/B _5274_/A _6848_/Q _3442_/X VGND VPWR _3446_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_366 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xmax_cap368 _5391_/A VGND VPWR _3781_/A2 VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_131_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6162_ _6897_/Q _5946_/X _5955_/X _6809_/Q VGND VPWR _6162_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_97_420 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3374_ _3374_/A hold85/X VGND VPWR _5301_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5113_ _5113_/A1 _4229_/X _5109_/Y _5112_/X VGND VPWR _5113_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6093_ _7051_/Q _5971_/A _5979_/X _6990_/Q VGND VPWR _6093_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold1305 _6518_/Q VGND VPWR _4103_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1316 hold1316/A VGND VPWR wb_dat_o[22] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_111_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1327 hold1424/X VGND VPWR hold1327/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5044_ _4948_/C _5042_/Y _5043_/Y _4948_/B VGND VPWR _5058_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_84_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_520 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1338 hold1338/A VGND VPWR wb_dat_o[7] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1349 _6311_/A1 VGND VPWR hold1349/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6995_ _7017_/CLK _6995_/D fanout458/X VGND VPWR _6995_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_41_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5946_ _5979_/A _5964_/A _5969_/C VGND VPWR _5946_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_43_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5877_ _6616_/Q _5628_/X _5910_/B1 _6627_/Q VGND VPWR _5877_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_166_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4828_ _4948_/B _4562_/Y _4827_/X _5027_/A VGND VPWR _4828_/X VGND VPWR sky130_fd_sc_hd__o211a_1
X_4759_ _4542_/A _4672_/B _4626_/Y _4689_/B VGND VPWR _4999_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_153_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6429_ _7155_/CLK _6429_/D fanout449/X VGND VPWR _6429_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_134_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_128 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_756 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_297 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_672 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_174 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_550 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold5/X VGND VPWR hold6/A VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_181_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5800_ _5799_/Y _5798_/X _6279_/S _5820_/A2 VGND VPWR _7112_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_6780_ _6969_/CLK _6780_/D fanout473/X VGND VPWR _6780_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3992_ hold804/X _6354_/A1 _3998_/S VGND VPWR _3992_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5731_ _6797_/Q _5905_/A2 _5715_/X _5730_/X VGND VPWR _5731_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_31_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_403 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5662_ _6802_/Q _5913_/B1 _5661_/X _6874_/Q _5659_/X VGND VPWR _5669_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4613_ _4716_/A _4636_/A VGND VPWR _4613_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_175_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5593_ _7100_/Q _7099_/Q VGND VPWR _5964_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_4544_ _4948_/A _4413_/Y _4561_/B _4562_/A VGND VPWR _4589_/B VGND VPWR sky130_fd_sc_hd__a211o_1
Xhold402 _4121_/X VGND VPWR _6534_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold413 _6626_/Q VGND VPWR hold413/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _5192_/X VGND VPWR _6769_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _7067_/Q VGND VPWR hold435/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 _5396_/X VGND VPWR _6950_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _4984_/A _4710_/A VGND VPWR _4650_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_144_686 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold457 _6692_/Q VGND VPWR hold457/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold468 _5279_/X VGND VPWR _6846_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6214_ _6631_/Q _5946_/X _5955_/X _6551_/Q VGND VPWR _6214_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold479 _6894_/Q VGND VPWR hold479/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _6832_/Q _5256_/A _3423_/X _3425_/X VGND VPWR _3426_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_7194_ hold91/A VGND VPWR _7194_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6145_ _7069_/Q _5934_/X _5975_/B _6872_/Q _6144_/X VGND VPWR _6145_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3357_ hold65/X _3454_/A VGND VPWR _3573_/B VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_112_572 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1102 _5305_/X VGND VPWR _6869_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_434 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1113 _7187_/A VGND VPWR _4065_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 _4241_/X VGND VPWR _6632_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6076_ _6789_/Q _6226_/B _6075_/X VGND VPWR _6076_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
Xhold1135 _6799_/Q VGND VPWR _5226_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ _6488_/Q _6414_/Q VGND VPWR _3288_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold1146 _4091_/X VGND VPWR _6512_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1157 _6874_/Q VGND VPWR _5311_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5027_ _5027_/A _5027_/B _5027_/C VGND VPWR _5080_/B VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1168 _4140_/X VGND VPWR _6550_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1179 _6858_/Q VGND VPWR _5293_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6978_ _7012_/CLK _6978_/D fanout458/X VGND VPWR _6978_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_179_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5929_ _6544_/Q _5652_/Y _5920_/X _5928_/X _6303_/S VGND VPWR _5929_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_179_594 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_756 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold980 _7153_/Q VGND VPWR hold980/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold991 _5182_/X VGND VPWR _5183_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_314 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_762 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4260_ hold499/X _5518_/A1 _4261_/S VGND VPWR _4260_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3211_ _6885_/Q VGND VPWR _3211_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4191_ _3640_/Y _4191_/A1 _4195_/S VGND VPWR _6594_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_79_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6901_ _7076_/CLK _6901_/D fanout481/X VGND VPWR _6901_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_47_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6832_ _6951_/CLK _6832_/D fanout474/X VGND VPWR _6832_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_6763_ _6953_/CLK _6763_/D fanout460/X VGND VPWR _6763_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3975_ hold40/X hold52/X _3975_/S VGND VPWR hold53/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_5714_ _5735_/A2 _5713_/X _6279_/S VGND VPWR _7108_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_6694_ _6714_/CLK _6694_/D fanout470/X VGND VPWR _6694_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_149_756 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5645_ _5664_/A _5666_/B _5660_/C VGND VPWR _5645_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_40_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_439 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5576_ _7094_/Q _5576_/B VGND VPWR _5576_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_117_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold210 _5177_/X VGND VPWR _6758_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 _6957_/Q VGND VPWR hold221/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _4542_/B _4453_/B _4525_/X _5084_/B VGND VPWR _4527_/X VGND VPWR sky130_fd_sc_hd__o211a_1
Xhold232 _5431_/X VGND VPWR _6981_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold243 hold243/A VGND VPWR hold243/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _5456_/X VGND VPWR _7003_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _6711_/Q VGND VPWR hold265/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold276 _5465_/X VGND VPWR _7011_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _4551_/A _4813_/A _4459_/B VGND VPWR _4953_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_49_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold287 _6819_/Q VGND VPWR hold287/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold298 _5267_/X VGND VPWR _6835_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_678 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3409_ _3409_/A _3409_/B wire357/X VGND VPWR _3410_/B VGND VPWR sky130_fd_sc_hd__nor3b_1
X_7177_ _7177_/A VGND VPWR _7177_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4389_ _4631_/D _4661_/A _4441_/B VGND VPWR _4389_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
X_6128_ _6128_/A0 _6127_/X _6303_/S VGND VPWR _6128_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_58_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6059_ _7058_/Q _5954_/X _5976_/D _6877_/Q _6058_/X VGND VPWR _6074_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_105 user_clock VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_116 _3251_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_127 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_138 _6440_/Q VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_54_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_149 _5494_/A1 VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_53_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_356 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_339 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_732 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_686 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_710 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_339 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_754 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_724 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_334 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_676 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3760_ _3760_/A _3760_/B _3760_/C _3760_/D VGND VPWR _3761_/D VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_9_530 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3691_ _7004_/Q _3370_/Y _4038_/A _6477_/Q VGND VPWR _3691_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_187_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5430_ hold357/X _5526_/A1 _5435_/S VGND VPWR _5430_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput304 _3450_/X VGND VPWR serial_data_1 VGND VPWR sky130_fd_sc_hd__buf_12
X_5361_ hold708/X _5469_/A1 _5363_/S VGND VPWR _5361_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput315 hold1325/X VGND VPWR hold1326/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput326 hold1359/X VGND VPWR hold1360/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput337 hold1327/X VGND VPWR hold1328/A VGND VPWR sky130_fd_sc_hd__buf_12
X_7100_ _7113_/CLK _7100_/D fanout464/X VGND VPWR _7100_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4312_ hold834/X _6354_/A1 _4315_/S VGND VPWR _4312_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5292_ _5292_/A _5505_/B VGND VPWR _5300_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_678 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7031_ _7086_/CLK hold51/X fanout484/X VGND VPWR _7031_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_113_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4243_ hold974/X _5546_/A1 _4243_/S VGND VPWR _4243_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4174_ _4174_/A0 _5492_/A1 _4177_/S VGND VPWR _4174_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_82_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6815_ _6969_/CLK _6815_/D fanout473/X VGND VPWR _6815_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_51_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6746_ _6746_/CLK _6746_/D fanout447/X VGND VPWR _6746_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3958_ _3958_/A input1/X VGND VPWR _3958_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_50_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6677_ _6677_/CLK _6677_/D fanout450/X VGND VPWR _6677_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3889_ _7097_/Q _7098_/Q VGND VPWR _5978_/A VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_136_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5628_ _5638_/A _5660_/C _5663_/C VGND VPWR _5628_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_164_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5559_ _7088_/Q _7089_/Q VGND VPWR _5604_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_183_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VPWR _7130_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
XPHY_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4930_ _4482_/B _4562_/Y _4741_/A _5099_/B _4758_/X VGND VPWR _4930_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_18_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4465_/B _4845_/X _4847_/A VGND VPWR _4869_/C VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_32_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6600_ _7036_/CLK _6600_/D fanout455/X VGND VPWR _6600_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3812_ _7173_/A _3320_/X _3355_/X _4268_/A _6665_/Q VGND VPWR _3812_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XANTENNA_16 _3571_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_177_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4792_ _4576_/B _4703_/B _4689_/Y VGND VPWR _4796_/A VGND VPWR sky130_fd_sc_hd__a21oi_2
XFILLER_193_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _4304_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_38 _4108_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_49 _5643_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6531_ _6990_/CLK hold39/X fanout479/X VGND VPWR _6531_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3743_ _6819_/Q _5247_/A _4032_/A _6471_/Q VGND VPWR _3743_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6462_ _6668_/CLK _6462_/D _6400_/A VGND VPWR _6462_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3674_ input22/X _3367_/Y _4310_/A _6702_/Q _3673_/X VGND VPWR _3679_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_134_718 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5413_ _5413_/A0 _5545_/A1 _5417_/S VGND VPWR _5413_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6393_ _6396_/A _6396_/B VGND VPWR _6393_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5344_ hold932/X _5548_/A1 _5345_/S VGND VPWR _5344_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput178 _3211_/Y VGND VPWR mgmt_gpio_oeb[12] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput189 _3201_/Y VGND VPWR mgmt_gpio_oeb[22] VGND VPWR sky130_fd_sc_hd__buf_12
X_5275_ _5275_/A0 hold666/X _5282_/S VGND VPWR _5275_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7014_ _7049_/CLK _7014_/D fanout457/X VGND VPWR _7014_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4226_ _6643_/Q _6642_/Q _6644_/Q VGND VPWR _4230_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_101_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4157_ _4157_/A _6352_/B VGND VPWR _4162_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_95_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_705 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4088_ hold257/X _5534_/A1 _5202_/B VGND VPWR _4088_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_587 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_350 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6729_ _3945_/A1 _6729_/D _6381_/X VGND VPWR _6729_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_109_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_52_csclk _7001_/CLK VGND VPWR _6537_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_164_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_540 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout394 hold174/X VGND VPWR hold22/A VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_27_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_440 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_698 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput14 mask_rev_in[19] VGND VPWR input14/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_167_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput25 mask_rev_in[29] VGND VPWR input25/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput36 mgmt_gpio_in[0] VGND VPWR _3958_/A VGND VPWR sky130_fd_sc_hd__buf_6
Xinput47 mgmt_gpio_in[1] VGND VPWR input47/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput58 mgmt_gpio_in[2] VGND VPWR _3251_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_183_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput69 mgmt_gpio_in[6] VGND VPWR input69/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold809 _4129_/X VGND VPWR _6541_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3390_ _6873_/Q _5301_/A _5541_/A _7086_/Q VGND VPWR _3390_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_170_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5060_ _5069_/A _5004_/Y _5038_/X _5059_/X VGND VPWR _5060_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_28_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1509 _7106_/Q VGND VPWR _5672_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4011_ _4011_/A0 _6355_/A1 _4013_/S VGND VPWR _4011_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_532 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5962_ _5978_/A _5969_/C _5979_/C VGND VPWR _5975_/B VGND VPWR sky130_fd_sc_hd__and3_4
X_4913_ _5051_/A _4782_/A _4881_/B VGND VPWR _5114_/C VGND VPWR sky130_fd_sc_hd__o21ai_1
X_5893_ _7037_/Q _5614_/X _5630_/X _6478_/Q VGND VPWR _5893_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_21_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_484 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4844_ _4686_/Y _5041_/C _4887_/A VGND VPWR _4869_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_138_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4775_ _4912_/A _4775_/B _5074_/A _4775_/D VGND VPWR _4776_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_20_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6514_ _6969_/CLK _6514_/D fanout473/X VGND VPWR _7180_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3726_ _6971_/Q _5418_/A _3585_/Y input96/X _3725_/X VGND VPWR _3729_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_684 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6445_ _7082_/CLK _6445_/D fanout483/X VGND VPWR _6445_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3657_ _7153_/Q _6352_/A _4014_/A _6457_/Q VGND VPWR _3657_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_164_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6376_ _6401_/A _6401_/B VGND VPWR _6376_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3588_ _6813_/Q _5238_/A _4157_/A _6568_/Q VGND VPWR _3588_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_102_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5327_ hold681/X _5540_/A1 _5327_/S VGND VPWR _5327_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5258_ hold285/X _5534_/A1 _5264_/S VGND VPWR _5258_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4209_ _4209_/A0 _6353_/A1 _4213_/S VGND VPWR _4209_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5189_ _5189_/A0 hold667/X _5189_/S VGND VPWR _5189_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_537 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_311 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_275 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4560_ _4563_/A _4631_/D _4563_/D VGND VPWR _4595_/A VGND VPWR sky130_fd_sc_hd__nand3_1
X_3511_ _3511_/A _3571_/B VGND VPWR _3511_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold606 _6865_/Q VGND VPWR hold606/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4491_ _4739_/A _4492_/D VGND VPWR _4491_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold617 _4019_/X VGND VPWR _6459_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _6877_/Q VGND VPWR hold628/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 _4247_/X VGND VPWR _6647_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6662_/Q _5976_/B _5971_/C _6712_/Q VGND VPWR _6230_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3442_ _6888_/Q _5319_/A _5301_/A _6872_/Q VGND VPWR _3442_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xmax_cap369 _3814_/A VGND VPWR _3455_/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_170_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_378 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6161_ _6945_/Q _5961_/X _6159_/X _6160_/X VGND VPWR _6165_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3373_ _3374_/A _3373_/B VGND VPWR _5319_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5112_ _5112_/A _5112_/B _5112_/C _5112_/D VGND VPWR _5112_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_6092_ _6822_/Q _5953_/X _5960_/X _7075_/Q _6091_/X VGND VPWR _6092_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1306 _4103_/X VGND VPWR _6518_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 hold1413/X VGND VPWR hold1317/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5043_ _5043_/A _5043_/B VGND VPWR _5043_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold1328 hold1328/A VGND VPWR wb_dat_o[30] VGND VPWR sky130_fd_sc_hd__buf_12
Xhold1339 hold1423/X VGND VPWR hold1339/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck _7149_/Q VGND VPWR clkbuf_0_wbbd_sck/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_53_524 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6994_ _7012_/CLK _6994_/D fanout458/X VGND VPWR _6994_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_179_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5945_ _5981_/A _5981_/C _5979_/C VGND VPWR _5945_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5876_ _6462_/Q _5624_/X _5654_/X _6677_/Q _5866_/Y VGND VPWR _5876_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_178_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_117 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4827_ _4948_/C _4810_/B _4825_/Y _4826_/X _4574_/Y VGND VPWR _4827_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_4758_ _4607_/A _4413_/Y _4947_/A _4611_/Y _4616_/Y VGND VPWR _4758_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_147_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3709_ _3709_/A _3709_/B _3709_/C VGND VPWR _3730_/A VGND VPWR sky130_fd_sc_hd__nor3_1
X_4689_ _4689_/A _4689_/B VGND VPWR _4689_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_161_120 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6428_ _7155_/CLK _6428_/D fanout449/X VGND VPWR _6428_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_161_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6359_ _6400_/A _6400_/B VGND VPWR _6359_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_88_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VPWR hold3/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3991_ _3991_/A0 _5491_/A1 _3998_/S VGND VPWR _3991_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_50_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5730_ _6989_/Q _5627_/X _5635_/X _6829_/Q VGND VPWR _5730_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_95_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5661_ _5638_/A _5667_/B _5663_/C VGND VPWR _5661_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_129_640 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4612_ _4975_/A _5010_/B VGND VPWR _4612_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_191_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5592_ _5592_/A1 _5594_/A _5591_/Y VGND VPWR _7099_/D VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_129_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4543_ _4948_/C _4456_/Y _4542_/X _4561_/B VGND VPWR _4589_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_128_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold403 _7052_/Q VGND VPWR hold403/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _4234_/X VGND VPWR _6626_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold425 _6631_/Q VGND VPWR hold425/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _5528_/X VGND VPWR _7067_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_507 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4474_ _4615_/B _4638_/A VGND VPWR _4710_/A VGND VPWR sky130_fd_sc_hd__and2_1
Xhold447 _6613_/Q VGND VPWR hold447/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _4301_/X VGND VPWR _6692_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 _6967_/Q VGND VPWR hold469/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6686_/Q _5961_/X _6207_/X _6212_/X VGND VPWR _6218_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_131_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3425_ input50/X _4058_/S _5211_/A _6792_/Q _3424_/X VGND VPWR _3425_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7193_ _7193_/A VGND VPWR _7193_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_131_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6144_ _7053_/Q _5971_/A _5979_/X _6992_/Q VGND VPWR _6144_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3356_ _3356_/A _3356_/B VGND VPWR _3511_/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_97_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1103 _7066_/Q VGND VPWR _5527_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _4065_/X VGND VPWR _6496_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6075_ _6069_/X _6301_/C _6075_/C _6075_/D VGND VPWR _6075_/X VGND VPWR sky130_fd_sc_hd__and4b_2
X_3287_ _3975_/S hold101/X _3285_/X VGND VPWR _3287_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
Xhold1125 _6452_/Q VGND VPWR _4011_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 _5226_/X VGND VPWR _6799_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 _6914_/Q VGND VPWR _5356_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 _5311_/X VGND VPWR _6874_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _4638_/Y _4695_/Y _4915_/B VGND VPWR _5027_/C VGND VPWR sky130_fd_sc_hd__o21a_1
Xhold1169 hold1593/X VGND VPWR _4070_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6977_ _7033_/CLK _6977_/D fanout464/X VGND VPWR _6977_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_81_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5928_ _6582_/Q _5928_/A2 _5923_/X _5927_/X VGND VPWR _5928_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_5859_ _6686_/Q _5632_/X _5642_/X _6716_/Q _5858_/X VGND VPWR _5862_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold970 _6659_/Q VGND VPWR hold970/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold981 _6355_/X VGND VPWR _7153_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_741 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold992 _5183_/X VGND VPWR _6763_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_326 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_376 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3210_ _6893_/Q VGND VPWR _3210_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4190_ _3700_/Y _4190_/A1 _4195_/S VGND VPWR _6593_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_178 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_424 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6900_ _6990_/CLK _6900_/D fanout479/X VGND VPWR _6900_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_35_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6831_ _6951_/CLK _6831_/D fanout474/X VGND VPWR _6831_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6762_ _6953_/CLK _6762_/D fanout460/X VGND VPWR _6762_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3974_ hold640/X _6357_/A1 _3980_/S VGND VPWR _3974_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5713_ _5713_/A0 _5712_/X _6303_/S VGND VPWR _5713_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6693_ _6714_/CLK _6693_/D fanout470/X VGND VPWR _6693_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_31_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5644_ _6962_/Q _5642_/X _5643_/X _6994_/Q VGND VPWR _5644_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_136_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5575_ _5610_/B _5658_/B _5667_/B _5575_/B1 _5568_/Y VGND VPWR _7093_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_191_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold200 _6797_/Q VGND VPWR hold200/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 _6754_/Q VGND VPWR hold211/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4526_ _4542_/B _4531_/B VGND VPWR _5084_/B VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold222 _5404_/X VGND VPWR _6957_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6569_/Q VGND VPWR hold233/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold244 _4122_/X VGND VPWR _6535_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _6762_/Q VGND VPWR hold255/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _4324_/X VGND VPWR _6711_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4459_/A _4724_/A _4579_/B VGND VPWR _4508_/C VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_131_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold277 _6691_/Q VGND VPWR hold277/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold288 _5249_/X VGND VPWR _6819_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold299 _6979_/Q VGND VPWR hold299/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _3408_/A _3408_/B _3408_/C _3408_/D VGND VPWR _3408_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_172_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7176_ _7176_/A VGND VPWR _7176_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4388_ _4642_/A _4441_/B VGND VPWR _4396_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_98_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6127_ _6791_/Q _6226_/B _6126_/X VGND VPWR _6127_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
X_3339_ hold36/X _3692_/A VGND VPWR hold37/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_39_660 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6058_ _7082_/Q _5976_/B _5971_/C _7042_/Q VGND VPWR _6058_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_39_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5009_ _4625_/B _4702_/Y _4981_/A VGND VPWR _5112_/C VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_73_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA_106 user_clock VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_117 input45/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_128 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_139 _3581_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_471 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_96 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_167 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_736 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_490 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_688 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3690_ _7065_/Q _5523_/A _3365_/Y input5/X _3689_/X VGND VPWR _3698_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput305 _3417_/X VGND VPWR serial_data_2 VGND VPWR sky130_fd_sc_hd__buf_12
X_5360_ hold473/X _5528_/A1 _5363_/S VGND VPWR _5360_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput316 hold1333/X VGND VPWR hold1334/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput327 hold1323/X VGND VPWR hold1324/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput338 hold1355/X VGND VPWR hold1356/A VGND VPWR sky130_fd_sc_hd__buf_12
X_4311_ _4311_/A0 _6353_/A1 _4315_/S VGND VPWR _4311_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5291_ hold327/X _5540_/A1 _5291_/S VGND VPWR _5291_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7030_ _7080_/CLK _7030_/D fanout478/X VGND VPWR _7030_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0__f__1177_ clkbuf_0__1177_/X VGND VPWR _4192_/A0 VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4242_ hold509/X _5518_/A1 _4243_/S VGND VPWR _4242_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4173_ hold999/X hold666/X _4177_/S VGND VPWR _4173_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6814_ _7058_/CLK _6814_/D fanout480/X VGND VPWR _6814_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_51_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6745_ _6746_/CLK _6745_/D fanout447/X VGND VPWR _6745_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3957_ _3957_/A _3957_/B VGND VPWR _3957_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_6676_ _7036_/CLK _6676_/D fanout455/X VGND VPWR _6676_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3888_ _6303_/S _3887_/Y _5610_/B VGND VPWR _6507_/D VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_109_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5627_ _5638_/A _5666_/C _5663_/C VGND VPWR _5627_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5558_ _5555_/Y _5564_/A _5558_/C VGND VPWR _7088_/D VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_3_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4509_ _4947_/B _4948_/C _4456_/Y _4496_/Y VGND VPWR _4509_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_132_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5489_ hold690/X _5513_/A1 hold50/X VGND VPWR _5489_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_120_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_178 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7159_ _3927_/A1 _7159_/D _6389_/X VGND VPWR _7159_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_100_340 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_563 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4860_ _4685_/A _5042_/B _4504_/X VGND VPWR _5023_/D VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3811_ _3958_/A _4118_/B _4250_/A _6650_/Q _3810_/X VGND VPWR _3817_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4791_ _4791_/A _4791_/B _5106_/A _4791_/D VGND VPWR _4791_/X VGND VPWR sky130_fd_sc_hd__and4_1
XANTENNA_17 _5154_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_28 _3585_/Y VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_39 _5291_/S VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_6530_ _6990_/CLK _6530_/D fanout479/X VGND VPWR _6530_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3742_ _3742_/A _3742_/B _3742_/C _3742_/D VGND VPWR _3761_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_146_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_671 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6461_ _6668_/CLK _6461_/D _6400_/A VGND VPWR _6461_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_173_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3673_ _6452_/Q _4008_/A _4304_/A _6697_/Q VGND VPWR _3673_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5412_ hold321/X _5526_/A1 _5417_/S VGND VPWR _5412_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_161_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6392_ _6396_/A _6396_/B VGND VPWR _6392_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5343_ hold429/X _5538_/A1 _5345_/S VGND VPWR _5343_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_143 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xoutput179 _3210_/Y VGND VPWR mgmt_gpio_oeb[13] VGND VPWR sky130_fd_sc_hd__buf_12
X_5274_ _5274_/A _5541_/B VGND VPWR _5282_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_7013_ _7082_/CLK _7013_/D fanout480/X VGND VPWR _7013_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4225_ hold820/X _5546_/A1 _4225_/S VGND VPWR _4225_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_563 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4156_ hold946/X _5546_/A1 _4156_/S VGND VPWR _4156_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4087_ _4087_/A0 _4086_/X _4101_/S VGND VPWR _4087_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_599 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4989_ _4542_/A _4428_/Y _4846_/B _4628_/Y VGND VPWR _4999_/C VGND VPWR sky130_fd_sc_hd__o22a_1
X_6728_ _3945_/A1 _6728_/D _6380_/X VGND VPWR _6728_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_183_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_362 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6659_ _6659_/CLK _6659_/D fanout468/X VGND VPWR _6659_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_125_708 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xfanout395 _5521_/A1 VGND VPWR _5548_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_74_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_599 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_452 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput15 mask_rev_in[1] VGND VPWR input15/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VPWR input26/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_167_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput37 mgmt_gpio_in[10] VGND VPWR input37/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput48 mgmt_gpio_in[20] VGND VPWR input48/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VPWR input59/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_183_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_270 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4010_ _4010_/A0 _5492_/A1 _4013_/S VGND VPWR _4010_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_77_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_544 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_257 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_503 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5961_ _5968_/A _5981_/A _5981_/B VGND VPWR _5961_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_547 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4912_ _4912_/A _5073_/A _4912_/C VGND VPWR _5083_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_33_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5892_ _6483_/Q _5643_/X _5910_/B1 _6628_/Q VGND VPWR _5892_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_772 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4843_ _4959_/A _4843_/B VGND VPWR _5041_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_33_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_660 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4774_ _5002_/A _4774_/B _4774_/C _5002_/B VGND VPWR _4775_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6513_ _6969_/CLK _6513_/D fanout473/X VGND VPWR _7179_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_20_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_535 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3725_ _6716_/Q _4328_/A _4322_/A _6711_/Q VGND VPWR _3725_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_174_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6444_ _7081_/CLK _6444_/D fanout479/X VGND VPWR _6444_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3656_ _6828_/Q _5256_/A _3654_/Y _3655_/X VGND VPWR _3661_/B VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_174_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6375_ _6400_/A _6400_/B VGND VPWR _6375_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3587_ _6997_/Q _5445_/A hold67/A _6468_/Q VGND VPWR _3587_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_774 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5326_ _5326_/A0 _5548_/A1 _5327_/S VGND VPWR _5326_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5257_ _5257_/A0 _5473_/A1 _5264_/S VGND VPWR _5257_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4208_ _4208_/A _4322_/B VGND VPWR _4213_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_180_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5188_ hold279/X _5534_/A1 _5189_/S VGND VPWR _5188_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4139_ _4139_/A _4322_/B VGND VPWR _4144_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_11_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_622 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_346 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_379 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_400 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_332 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3510_ _3555_/A _3577_/B VGND VPWR _4244_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_7_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4490_ _4689_/A _4490_/B VGND VPWR _4490_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold607 _5300_/X VGND VPWR _6865_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _6899_/Q VGND VPWR hold618/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _5314_/X VGND VPWR _6877_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ _6976_/Q _5418_/A _3326_/Y _6800_/Q _3440_/X VGND VPWR _3446_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6160_ _7017_/Q _5940_/X _5967_/X _6857_/Q _6158_/X VGND VPWR _6160_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3372_ _3546_/A _3717_/B VGND VPWR _3372_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_111_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5111_ _4482_/A _4625_/B _4615_/Y _4650_/Y _5110_/X VGND VPWR _5112_/D VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6091_ _6910_/Q _5973_/A _5948_/X _6950_/Q _6090_/X VGND VPWR _6091_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_85_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1307 _6545_/Q VGND VPWR _4134_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 hold1318/A VGND VPWR wb_dat_o[23] VGND VPWR sky130_fd_sc_hd__buf_12
X_5042_ _5051_/A _5042_/B VGND VPWR _5042_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_78_680 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1329 hold1425/X VGND VPWR hold1329/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_363 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6993_ _7053_/CLK _6993_/D fanout459/X VGND VPWR _6993_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_53_536 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_csclk _7001_/CLK VGND VPWR _6865_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_80_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5944_ _5978_/A _5964_/A _5981_/A VGND VPWR _5944_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5875_ _6557_/Q _5667_/X _5870_/X _5872_/X _5874_/X VGND VPWR _5875_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_33_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4826_ _4902_/A _4810_/B _4948_/B VGND VPWR _4826_/X VGND VPWR sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_66_csclk _6447_/CLK VGND VPWR _7012_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4757_ _4581_/B _4542_/D _4611_/Y _4653_/Y VGND VPWR _4770_/B VGND VPWR sky130_fd_sc_hd__o22a_1
X_3708_ _6947_/Q _3781_/A2 _3964_/A _6419_/Q _3707_/X VGND VPWR _3709_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4688_ _4689_/A _4619_/Y _4631_/Y _4902_/B _5108_/A VGND VPWR _4722_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_107_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6427_ _6747_/CLK _6427_/D fanout449/X VGND VPWR _6427_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_162_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3639_ _3639_/A _3639_/B _3639_/C VGND VPWR _3640_/D VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_161_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6358_ _6400_/A _6400_/B VGND VPWR _6358_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_88_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5309_ hold738/X _5540_/A1 _5309_/S VGND VPWR _5309_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6289_ _6289_/A _6289_/B _6289_/C VGND VPWR _6289_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_88_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6890_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_95 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_116 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VPWR hold4/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xnet399_2 net399_2/A VGND VPWR _3941_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_3990_ _3990_/A _6352_/B VGND VPWR _3998_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_62_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5660_ _5664_/A _5667_/C _5660_/C VGND VPWR _5660_/X VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_31_764 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4611_ _4753_/B _4611_/B VGND VPWR _4611_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
X_5591_ _7099_/Q _5574_/Y _5594_/A VGND VPWR _5591_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_129_652 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4542_ _4542_/A _4542_/B _4948_/B _4542_/D VGND VPWR _4542_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_129_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold404 _5511_/X VGND VPWR _7052_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold415 _6646_/Q VGND VPWR hold415/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _4240_/X VGND VPWR _6631_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4739_/A _4642_/A VGND VPWR _4638_/A VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_116_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold437 _6974_/Q VGND VPWR hold437/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _4213_/X VGND VPWR _6613_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold459 _6854_/Q VGND VPWR hold459/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6476_/Q _5940_/X _5967_/X _6605_/Q _6206_/X VGND VPWR _6212_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3424_ _6856_/Q _5283_/A _3370_/Y _7008_/Q VGND VPWR _3424_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7192_ _7192_/A VGND VPWR _7192_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6143_ _6824_/Q _5953_/X _5960_/X _7077_/Q _6142_/X VGND VPWR _6143_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3355_ _3356_/A _3355_/B hold72/X VGND VPWR _3355_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_97_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1104 _5527_/X VGND VPWR _7066_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6074_ _6074_/A _6074_/B _6074_/C _6074_/D VGND VPWR _6075_/D VGND VPWR sky130_fd_sc_hd__nor4_1
Xhold1115 _7179_/A VGND VPWR _4093_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3286_ _3975_/S hold101/X hold204/X VGND VPWR _3286_/X VGND VPWR sky130_fd_sc_hd__a21o_4
Xhold1126 _4011_/X VGND VPWR _6452_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 _7192_/A VGND VPWR _5197_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5025_ _4413_/Y _4902_/A _4616_/Y _4691_/A _4877_/B VGND VPWR _5118_/B VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold1148 _5356_/X VGND VPWR _6914_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _7189_/A VGND VPWR _5194_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6976_ _7082_/CLK _6976_/D fanout483/X VGND VPWR _6976_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_41_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_9 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5927_ _6689_/Q _5632_/X _5924_/X _5926_/X VGND VPWR _5927_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_22_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5858_ _6561_/Q _5631_/X _5667_/X _6556_/Q VGND VPWR _5858_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_70_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4809_ _4992_/A _4886_/B VGND VPWR _4810_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_5789_ _7016_/Q _5630_/X _5658_/X _6888_/Q _5788_/X VGND VPWR _5797_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_107_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold960 _6457_/Q VGND VPWR hold960/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold971 _4261_/X VGND VPWR _6659_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _6618_/Q VGND VPWR hold982/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _6428_/Q VGND VPWR hold993/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_666 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_539 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_672 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6830_ _6884_/CLK _6830_/D fanout475/X VGND VPWR _6830_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_62_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6761_ _6953_/CLK _6761_/D fanout459/X VGND VPWR _6761_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_16_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3973_ hold58/X _3973_/A1 _3975_/S VGND VPWR _3973_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_50_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5712_ _5706_/Y _5711_/Y _6788_/Q _5652_/Y VGND VPWR _5712_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_6692_ _6714_/CLK _6692_/D fanout470/X VGND VPWR _6692_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_31_583 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5643_ _5664_/A _5660_/C _5663_/C VGND VPWR _5643_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_176_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_460 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5574_ _6506_/Q _5610_/B VGND VPWR _5574_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold201 _5224_/X VGND VPWR _6797_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _4948_/A _4453_/B _4522_/X _5084_/A VGND VPWR _4525_/X VGND VPWR sky130_fd_sc_hd__o211a_1
Xhold212 _5170_/X VGND VPWR _6754_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _6837_/Q VGND VPWR hold223/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_463 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold234 _4162_/X VGND VPWR _6569_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _6923_/Q VGND VPWR hold245/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold256 _5181_/X VGND VPWR _6762_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4456_/A _4579_/B VGND VPWR _4456_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_131_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold267 _6661_/Q VGND VPWR hold267/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _4300_/X VGND VPWR _6691_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 _6795_/Q VGND VPWR hold289/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ _6913_/Q _5346_/A _5238_/A _6817_/Q _3406_/X VGND VPWR _3408_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7175_ _7175_/A VGND VPWR _7175_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4387_ _4661_/A _4441_/B VGND VPWR _4400_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_131_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6126_ _6118_/X _6226_/B _6126_/C _6126_/D VGND VPWR _6126_/X VGND VPWR sky130_fd_sc_hd__and4b_2
XFILLER_100_511 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3338_ _3454_/B _3415_/B VGND VPWR _3692_/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_100_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6057_ _6813_/Q _5971_/B _5949_/X _6933_/Q _6056_/X VGND VPWR _6074_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3269_ _6390_/A _6396_/B VGND VPWR _3269_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_73_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5008_ _5008_/A _5008_/B _5008_/C _5008_/D VGND VPWR _5112_/B VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_39_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_107 wb_clk_i VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_118 input38/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_129 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_121_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_303 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_483 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6959_ _6999_/CLK _6959_/D fanout465/X VGND VPWR _6959_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_14_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold790 _6831_/Q VGND VPWR hold790/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1490 _6078_/X VGND VPWR _7122_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_494 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_509 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VPWR _3927_/A1 VGND
+ VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput306 _3940_/X VGND VPWR serial_load VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput317 hold1353/X VGND VPWR hold1354/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput328 hold1315/X VGND VPWR hold1316/A VGND VPWR sky130_fd_sc_hd__buf_12
X_4310_ _4310_/A _6352_/B VGND VPWR _4315_/S VGND VPWR sky130_fd_sc_hd__and2_2
Xoutput339 hold1369/X VGND VPWR hold1370/A VGND VPWR sky130_fd_sc_hd__buf_12
X_5290_ hold141/X hold99/X _5291_/S VGND VPWR _5290_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4241_ _4241_/A0 _5493_/A1 _4243_/S VGND VPWR _4241_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4172_ _4172_/A _5490_/B VGND VPWR _4177_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_95_575 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6813_ _7076_/CLK _6813_/D fanout481/X VGND VPWR _6813_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_90_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6744_ _6746_/CLK _6744_/D _3946_/B VGND VPWR _6744_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3956_ _3956_/A _3956_/B VGND VPWR _3956_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_188_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_380 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_19 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6675_ _7036_/CLK _6675_/D fanout455/X VGND VPWR _6675_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3887_ _5606_/A _3887_/B VGND VPWR _3887_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_5626_ _6978_/Q _5624_/X _5625_/X _7002_/Q VGND VPWR _5626_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_136_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5557_ _7088_/Q _5562_/D VGND VPWR _5558_/C VGND VPWR sky130_fd_sc_hd__nand2_1
X_4508_ _4507_/X _5027_/A _4508_/C _4508_/D VGND VPWR _4508_/X VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_117_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5488_ hold894/X _5548_/A1 hold50/X VGND VPWR _5488_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4439_ _4615_/B _4635_/B VGND VPWR _4672_/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_132_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_712 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7158_ _3927_/A1 _7158_/D _6388_/X VGND VPWR _7158_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_59_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6109_ _7015_/Q _5940_/X _5967_/X _6855_/Q _6107_/X VGND VPWR _6109_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7089_ _7113_/CLK _7089_/D fanout460/X VGND VPWR _7089_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_73_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_344 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_680 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_586 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_686 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3810_ input71/X _3331_/Y _4196_/A _6599_/Q VGND VPWR _3810_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4790_ _4556_/A _4632_/B _4482_/A _4672_/A _4789_/X VGND VPWR _4791_/D VGND VPWR
+ sky130_fd_sc_hd__o41a_1
XANTENNA_18 _5164_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_29 _5166_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3741_ input47/X _4118_/B _4310_/A _6701_/Q _3740_/X VGND VPWR _3742_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_650 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6460_ _6668_/CLK _6460_/D _6400_/A VGND VPWR _6460_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3672_ _6547_/Q _4133_/A _5490_/A _7036_/Q _3671_/X VGND VPWR _3679_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5411_ _5411_/A0 hold13/X _5417_/S VGND VPWR _5411_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6391_ _6396_/A _6396_/B VGND VPWR _6391_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5342_ hold184/X _5519_/A1 _5345_/S VGND VPWR _5342_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_126_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5273_ hold632/X _5513_/A1 _5273_/S VGND VPWR _5273_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7012_ _7012_/CLK _7012_/D fanout466/X VGND VPWR _7012_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_99_188 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4224_ hold309/X _5518_/A1 _4225_/S VGND VPWR _4224_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_101_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4155_ hold463/X _5518_/A1 _4156_/S VGND VPWR _4155_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4086_ _5203_/A0 _5473_/A1 _5202_/B VGND VPWR _4086_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_450 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4988_ _4919_/X _4945_/Y _4987_/X _5006_/A _4988_/B2 VGND VPWR _6722_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_6727_ _3568_/A1 _6727_/D _6379_/X VGND VPWR _6727_/Q VGND VPWR sky130_fd_sc_hd__dfrtn_1
X_3939_ _7103_/Q _6759_/Q _6762_/Q VGND VPWR _3939_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_149_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_160 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6658_ _6659_/CLK _6658_/D fanout469/X VGND VPWR _6658_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5609_ _5609_/A1 _5606_/B _5608_/X _3886_/B VGND VPWR _7105_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_124_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6589_ _7137_/CLK _6589_/D VGND VPWR _6589_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_152_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout396 hold99/X VGND VPWR _5521_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_143_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_133 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_464 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput16 mask_rev_in[20] VGND VPWR input16/X VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput27 mask_rev_in[30] VGND VPWR input27/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput38 mgmt_gpio_in[11] VGND VPWR input38/X VGND VPWR sky130_fd_sc_hd__clkbuf_4
XFILLER_116_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput49 mgmt_gpio_in[21] VGND VPWR input49/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_182_152 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_398 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5960_ _5969_/A _5966_/A _5981_/C VGND VPWR _5960_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_18_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4911_ _4911_/A _4911_/B _4911_/C VGND VPWR _4912_/C VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_80_559 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5891_ _6473_/Q _5627_/X _5667_/X _6558_/Q _5890_/X VGND VPWR _5896_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4842_ _4947_/B _4542_/D _4623_/Y _4694_/Y VGND VPWR _4875_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_193_406 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4773_ _4773_/A _4928_/A VGND VPWR _5002_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_119_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6512_ _6969_/CLK _6512_/D fanout473/X VGND VPWR _6512_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3724_ input53/X _5193_/A _4145_/A _6556_/Q _3723_/X VGND VPWR _3729_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_547 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6443_ _7017_/CLK _6443_/D fanout458/X VGND VPWR _6443_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3655_ _6844_/Q _5274_/A _5166_/A _6753_/Q VGND VPWR _3655_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_161_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6374_ _6401_/A _6401_/B VGND VPWR _6374_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3586_ _3586_/A _3814_/A VGND VPWR _5166_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5325_ hold788/X _5538_/A1 _5327_/S VGND VPWR _5325_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5256_ _5256_/A _5505_/B VGND VPWR _5264_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_102_458 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4207_ hold529/X _6357_/A1 _4207_/S VGND VPWR _4207_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5187_ hold441/X _5544_/A1 _5189_/S VGND VPWR _5187_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4138_ hold962/X _5546_/A1 _4138_/S VGND VPWR _4138_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4069_ _4119_/A0 _5491_/A1 _4118_/B VGND VPWR _4069_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_366 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_667 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_648 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_762 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_652 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold608 _6544_/Q VGND VPWR hold608/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold619 _5339_/X VGND VPWR _6899_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _6992_/Q _5436_/A _5373_/A _6936_/Q VGND VPWR _3440_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3371_ _3586_/A _3717_/B VGND VPWR _3981_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5110_ _4483_/Y _4625_/B _4716_/Y _4484_/Y _5006_/A VGND VPWR _5110_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_88_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6090_ _6902_/Q _5976_/C _5971_/D _6830_/Q VGND VPWR _6090_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5041_ _5041_/A _5041_/B _5041_/C VGND VPWR _5041_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_69_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1308 _4134_/X VGND VPWR _6545_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1319 hold1414/X VGND VPWR hold1319/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VPWR clkbuf_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_375 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6992_ _7069_/CLK _6992_/D fanout482/X VGND VPWR _6992_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_53_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5943_ _5979_/A _5969_/C _5979_/C VGND VPWR _5943_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_34_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5874_ _6482_/Q _5643_/X _5664_/X _6667_/Q _5873_/X VGND VPWR _5874_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4825_ _4551_/A _4815_/Y _4812_/Y VGND VPWR _4825_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_193_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4756_ _4542_/B _4672_/B _4626_/Y _4645_/Y VGND VPWR _4771_/C VGND VPWR sky130_fd_sc_hd__o22a_1
X_3707_ _6851_/Q _5283_/A _5409_/A _6963_/Q VGND VPWR _3707_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4687_ _4469_/A _4644_/Y _4663_/Y _4689_/A VGND VPWR _5108_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_162_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6426_ _6747_/CLK _6426_/D fanout449/X VGND VPWR _6426_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3638_ _3638_/A _3638_/B _3638_/C _3638_/D VGND VPWR _3639_/C VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_162_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6357_ hold566/X _6357_/A1 _6357_/S VGND VPWR _6357_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3569_ _3573_/A _3692_/A VGND VPWR _4008_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5308_ hold716/X _5521_/A1 _5309_/S VGND VPWR _5308_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_391 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6288_ _6464_/Q _5945_/X _5975_/C _6582_/Q _6287_/X VGND VPWR _6289_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_102_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5239_ _5239_/A0 hold667/X _5246_/S VGND VPWR _5239_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_102_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_331 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_303 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_358 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VPWR hold5/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4610_ _4753_/B _4611_/B VGND VPWR _5010_/B VGND VPWR sky130_fd_sc_hd__and2_2
X_5590_ _5610_/B _5978_/A _5979_/A _5568_/Y _5590_/B2 VGND VPWR _7098_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_4541_ _4661_/A _4724_/A _4959_/B _3962_/A VGND VPWR _4541_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_190_217 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire380 _4674_/Y VGND VPWR wire380/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xhold405 hold405/A VGND VPWR hold405/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 _4246_/X VGND VPWR _6646_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ _4472_/A _4489_/B VGND VPWR _4472_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_143_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold427 _6656_/Q VGND VPWR hold427/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _5423_/X VGND VPWR _6974_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _6911_/Q VGND VPWR hold449/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6691_/Q _5954_/X _5976_/D _6620_/Q _6210_/X VGND VPWR _6225_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_3423_ _6864_/Q _5292_/A _5337_/A _6904_/Q VGND VPWR _3423_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7191_ _7191_/A VGND VPWR _7191_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6142_ _6912_/Q _5973_/A _5948_/X _6952_/Q _6141_/X VGND VPWR _6142_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3354_ _3571_/A _3373_/B VGND VPWR _5247_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_6073_ _7029_/Q _5944_/X _5975_/A _6845_/Q _6072_/X VGND VPWR _6074_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_57_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1105 _6917_/Q VGND VPWR _5359_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3285_ _3975_/S _3285_/B VGND VPWR _3285_/X VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_100_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1116 _4093_/X VGND VPWR _6513_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 _6552_/Q VGND VPWR _4142_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5024_ _5051_/B _5024_/B VGND VPWR _5086_/C VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold1138 _5197_/X VGND VPWR _6773_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 _6906_/Q VGND VPWR _5347_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6975_ _7016_/CLK _6975_/D fanout474/X VGND VPWR _6975_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_13_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5926_ _6479_/Q _5630_/X _5638_/X _6709_/Q _5925_/X VGND VPWR _5926_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5857_ _6651_/Q _5646_/X _5928_/A2 _6579_/Q _5856_/X VGND VPWR _5862_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4808_ _5068_/B _4805_/X _4964_/A VGND VPWR _4884_/C VGND VPWR sky130_fd_sc_hd__a21bo_1
XFILLER_186_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5788_ _6448_/Q _5614_/X _5814_/B1 _6912_/Q VGND VPWR _5788_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4739_ _4739_/A _4739_/B VGND VPWR _4740_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_5_419 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6409_ _3568_/A1 _6409_/D _6365_/X VGND VPWR hold81/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xhold950 _6744_/Q VGND VPWR hold950/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _4017_/X VGND VPWR _6457_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _6702_/Q VGND VPWR hold972/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _4219_/X VGND VPWR _6618_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_531 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold994 _3984_/X VGND VPWR _6428_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_404 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_383 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_676 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_707 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_678 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk _7001_/CLK VGND VPWR _6999_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_140_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_65_csclk _6447_/CLK VGND VPWR _7006_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_94_289 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6760_ _6953_/CLK _6760_/D fanout459/X VGND VPWR _6760_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_90_495 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3972_ hold784/X _6356_/A1 _3980_/S VGND VPWR _3972_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5711_ _5711_/A _5711_/B _5711_/C VGND VPWR _5711_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_50_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6691_ _6712_/CLK _6691_/D fanout470/X VGND VPWR _6691_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_148_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5642_ _5664_/A _5657_/B _5660_/C VGND VPWR _5642_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5573_ _6506_/Q _5610_/B VGND VPWR _5602_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_129_483 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold202 _6488_/Q VGND VPWR hold202/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _4584_/A _4724_/A VGND VPWR _5084_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold213 _6464_/Q VGND VPWR hold213/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _5269_/X VGND VPWR _6837_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VPWR _7083_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold235 _7038_/Q VGND VPWR hold235/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _5366_/X VGND VPWR _6923_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ _4498_/A _4579_/B VGND VPWR _4948_/C VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold257 _6779_/Q VGND VPWR hold257/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_188 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold268 _4264_/X VGND VPWR _6661_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 _6766_/Q VGND VPWR hold279/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _6881_/Q _5310_/A _5229_/A _6809_/Q VGND VPWR _3406_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7174_ _7174_/A VGND VPWR _7174_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4386_ _4661_/A _4441_/B VGND VPWR _4563_/D VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_131_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6125_ _6125_/A _6125_/B _6125_/C _6125_/D VGND VPWR _6126_/D VGND VPWR sky130_fd_sc_hd__nor4_1
X_3337_ _3453_/A hold64/X _3415_/B VGND VPWR _5186_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_100_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6056_ _6445_/Q _5601_/X _5959_/X _6965_/Q VGND VPWR _6056_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3268_ _6764_/Q _6813_/Q _3268_/C VGND VPWR _3268_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_100_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5007_ _4576_/Y _4710_/Y _4482_/A VGND VPWR _5008_/D VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_73_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3199_ _6981_/Q VGND VPWR _3199_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_38_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_108 input92/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XANTENNA_119 _3899_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_14_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6958_ _7065_/CLK _6958_/D fanout465/X VGND VPWR _6958_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_81_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5909_ _5908_/Y _5907_/X _6279_/S _5909_/B2 VGND VPWR _7117_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_6889_ _6969_/CLK _6889_/D fanout475/X VGND VPWR _6889_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_139_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_559 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold780 _6847_/Q VGND VPWR hold780/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold791 _5262_/X VGND VPWR _6831_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_404 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1480 _6638_/Q VGND VPWR _3880_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _7121_/Q VGND VPWR _6053_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_698 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_375 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _3939_/X VGND VPWR serial_resetn VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_153_250 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput318 hold1343/X VGND VPWR hold1344/A VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput329 hold1317/X VGND VPWR hold1318/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_114_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_434 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4240_ hold425/X _5534_/A1 _4243_/S VGND VPWR _4240_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4171_ _3410_/Y _4171_/A1 _4171_/S VGND VPWR _6577_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6812_ _6990_/CLK _6812_/D fanout478/X VGND VPWR _6812_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_23_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6743_ _6746_/CLK _6743_/D _3946_/B VGND VPWR _6743_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3955_ _6643_/Q _3961_/B VGND VPWR _6637_/D VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_176_342 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6674_ _6674_/CLK _6674_/D fanout468/X VGND VPWR _6674_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3886_ _7088_/Q _3886_/B _7090_/Q _7091_/Q VGND VPWR _3887_/B VGND VPWR sky130_fd_sc_hd__nand4b_1
XFILLER_137_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5625_ _5638_/A _5667_/B _5663_/C VGND VPWR _5625_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5556_ _5552_/B _3887_/B _5554_/Y _6509_/Q VGND VPWR _5564_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_4507_ _4782_/A _4493_/B _4472_/X _4502_/X _4450_/Y VGND VPWR _4507_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
X_5487_ _5487_/A0 hold42/X hold50/X VGND VPWR hold51/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4438_ _4615_/B _4635_/B VGND VPWR _4965_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7157_ _7157_/CLK _7157_/D _3269_/X VGND VPWR _7157_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4369_ _4556_/A _4441_/A VGND VPWR _4454_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_59_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6108_ _7007_/Q _5958_/X _5978_/X _6999_/Q VGND VPWR _6108_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_58_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7088_ _7113_/CLK _7088_/D fanout460/X VGND VPWR _7088_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_58_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6039_ _6980_/Q _5945_/X _5975_/C _6836_/Q _6038_/X VGND VPWR _6040_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_73_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_495 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_392 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_112 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _5164_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_3740_ _6795_/Q _3326_/Y _4292_/A _6686_/Q VGND VPWR _3740_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_186_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3671_ _6932_/Q _5373_/A _4274_/A _6672_/Q VGND VPWR _3671_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5410_ _5410_/A0 _5524_/A1 _5417_/S VGND VPWR _5410_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6390_ _6390_/A _6396_/B VGND VPWR _6390_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_5341_ _5341_/A0 _5545_/A1 _5345_/S VGND VPWR _5341_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5272_ hold135/X hold99/X _5273_/S VGND VPWR _5272_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7011_ _7011_/CLK _7011_/D fanout456/X VGND VPWR _7011_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4223_ hold487/X _5544_/A1 _4225_/S VGND VPWR _4223_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4154_ hold596/X _5544_/A1 _4156_/S VGND VPWR _4154_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4085_ _6367_/B _3379_/A _5202_/B _4050_/X _4322_/B VGND VPWR _4101_/S VGND VPWR
+ sky130_fd_sc_hd__o221a_4
XFILLER_55_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_462 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4987_ _5039_/A _5039_/C _4963_/Y _4986_/X VGND VPWR _4987_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_11_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6726_ _7140_/CLK _6726_/D _6307_/B VGND VPWR _6726_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3938_ _6515_/Q input93/X _6767_/Q VGND VPWR _3938_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_109_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6657_ _6659_/CLK _6657_/D fanout468/X VGND VPWR _6657_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3869_ _3911_/B1 _3869_/A2 _3832_/B _6405_/Q VGND VPWR _6405_/D VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_164_334 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5608_ _7088_/Q _6509_/Q _5608_/C VGND VPWR _5608_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_6588_ _7137_/CLK _6588_/D VGND VPWR _6588_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_127_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5539_ hold898/X _5548_/A1 _5540_/S VGND VPWR _5539_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_133_765 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xfanout375 _6304_/S VGND VPWR _6279_/S VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_101_662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout397 hold108/X VGND VPWR hold99/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_59_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xinput17 mask_rev_in[21] VGND VPWR input17/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_168_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput28 mask_rev_in[31] VGND VPWR input28/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput39 mgmt_gpio_in[12] VGND VPWR _3960_/B VGND VPWR sky130_fd_sc_hd__buf_2
XFILLER_183_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_727 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4910_ _4691_/A _4482_/A _4672_/A _4964_/B _4909_/Y VGND VPWR _4915_/C VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_45_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5890_ _6708_/Q _5638_/X _5928_/A2 _6581_/Q VGND VPWR _5890_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4841_ _4493_/B _4911_/B _4472_/X VGND VPWR _4841_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_21_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_284 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4772_ _4772_/A _5099_/C _4772_/C _4772_/D VGND VPWR _4774_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_159_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6511_ _6969_/CLK _6511_/D fanout473/X VGND VPWR _6511_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3723_ _6769_/Q _5190_/A _5190_/B _4274_/A _6671_/Q VGND VPWR _3723_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6442_ _6926_/CLK _6442_/D fanout458/X VGND VPWR _6442_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3654_ hold85/A _3562_/B _3511_/A VGND VPWR _3654_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_173_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6373_ _6400_/A _6400_/B VGND VPWR _6373_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_161_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_0_0_wb_clk_i clkbuf_3_1_0_wb_clk_i/A VGND VPWR _7126_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_3585_ hold48/A _3714_/B VGND VPWR _3585_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5324_ hold798/X _5528_/A1 _5327_/S VGND VPWR _5324_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5255_ hold746/X _5540_/A1 _5255_/S VGND VPWR _5255_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4206_ hold730/X _6356_/A1 _4207_/S VGND VPWR _4206_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5186_ _5186_/A _5190_/B hold16/X VGND VPWR _5189_/S VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_56_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4137_ hold760/X _6356_/A1 _4138_/S VGND VPWR _4137_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4068_ _6396_/B _3546_/A _4118_/B _4050_/X _4322_/B VGND VPWR _4084_/S VGND VPWR
+ sky130_fd_sc_hd__o221a_4
XFILLER_83_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6709_ _6709_/CLK _6709_/D fanout445/X VGND VPWR _6709_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_137_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_378 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_679 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_30 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold609 _4132_/X VGND VPWR _6544_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3370_ _3370_/A hold74/X VGND VPWR _3370_/Y VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_170_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5040_ _4574_/A _4816_/Y _4950_/X VGND VPWR _5089_/B VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_26_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1309 _6470_/Q VGND VPWR _4033_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6991_ _7086_/CLK _6991_/D fanout484/X VGND VPWR _6991_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_93_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5942_ _7099_/Q _7100_/Q VGND VPWR _5979_/C VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_80_379 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5873_ _6562_/Q _5631_/X _5646_/X _6652_/Q VGND VPWR _5873_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4824_ _4542_/D _4562_/Y _4522_/D VGND VPWR _4824_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_193_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4755_ _4542_/A _4581_/B _4611_/Y _4628_/Y VGND VPWR _4755_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_3706_ input35/X _3365_/Y _5301_/A _6867_/Q _3705_/X VGND VPWR _3709_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4686_ _4911_/B _4686_/B VGND VPWR _4686_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_134_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_624 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6425_ _6926_/CLK _6425_/D fanout457/X VGND VPWR _6425_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_174_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3637_ _7029_/Q hold49/A _4328_/A _6718_/Q _3636_/X VGND VPWR _3638_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_146_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6356_ hold768/X _6356_/A1 _6357_/S VGND VPWR _6356_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3568_ _3568_/A1 _4118_/B hold37/A input48/X _3567_/X VGND VPWR _3580_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_88_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5307_ hold513/X _5538_/A1 _5309_/S VGND VPWR _5307_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6287_ _6669_/Q _5938_/X _5952_/X _6709_/Q VGND VPWR _6287_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3499_ _3573_/A _3562_/B VGND VPWR _4280_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_88_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5238_ _5238_/A _5541_/B VGND VPWR _5246_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_29_535 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5169_ hold367/X _5526_/A1 _5170_/S VGND VPWR _5169_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_343 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_202 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_654 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_87 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold6 hold6/A VGND VPWR hold6/X VGND VPWR sky130_fd_sc_hd__buf_8
XFILLER_59_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_516 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_265 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4540_ _4661_/A _4724_/A _4959_/B _3962_/A VGND VPWR _5039_/A VGND VPWR sky130_fd_sc_hd__a31oi_4
XFILLER_156_451 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_698 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_229 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire381 _5975_/Y VGND VPWR _5977_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold406 _4080_/X VGND VPWR _6503_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ _4702_/C _4471_/B _4471_/C VGND VPWR _4489_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_128_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold417 _6895_/Q VGND VPWR hold417/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _4258_/X VGND VPWR _6656_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold439 _6990_/Q VGND VPWR hold439/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6661_/Q _5976_/B _5971_/C _6711_/Q VGND VPWR _6210_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3422_ _6840_/Q _5265_/A _3414_/Y _3419_/X _3421_/X VGND VPWR _3431_/A VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
X_7190_ _7190_/A VGND VPWR _7190_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6141_ _6904_/Q _5976_/C _5971_/D _6832_/Q VGND VPWR _6141_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3353_ _3814_/A _3373_/B VGND VPWR _5532_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6072_ _7021_/Q _5937_/X _5975_/D _6885_/Q VGND VPWR _6072_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3284_ hold62/X hold202/X _3283_/Y VGND VPWR _3284_/X VGND VPWR sky130_fd_sc_hd__a21bo_1
Xhold1106 _5359_/X VGND VPWR _6917_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 _6667_/Q VGND VPWR _4271_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 _4142_/X VGND VPWR _6552_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _5023_/A _5023_/B _5023_/C _5023_/D VGND VPWR _5115_/A VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1139 _6768_/Q VGND VPWR _5191_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6974_ _6990_/CLK _6974_/D fanout480/X VGND VPWR _6974_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5925_ _7155_/Q _5625_/X _5661_/X _6623_/Q VGND VPWR _5925_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5856_ _6551_/Q _5913_/B1 _5855_/Y _5652_/B VGND VPWR _5856_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4807_ _4846_/B _4645_/Y _4653_/Y _4689_/A VGND VPWR _4807_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_5787_ _5787_/A _5787_/B _5787_/C VGND VPWR _5787_/Y VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_119_131 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4738_ _4738_/A VGND VPWR _4738_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_119_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4669_ _4739_/A _5043_/A _4747_/B _4739_/B VGND VPWR _4676_/B VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_174_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6408_ _3568_/A1 _6408_/D _6364_/X VGND VPWR hold24/A VGND VPWR sky130_fd_sc_hd__dfrtp_2
Xhold940 _6896_/Q VGND VPWR hold940/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _5157_/X VGND VPWR _6744_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _6549_/Q VGND VPWR hold962/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_370 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold973 _4313_/X VGND VPWR _6702_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 _6436_/Q VGND VPWR hold984/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6642_/Q _6339_/A2 _6339_/B1 _6350_/A2 _6338_/X VGND VPWR _6339_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold995 _6739_/Q VGND VPWR hold995/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_395 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_151 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_154 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_101 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_630 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3971_ hold93/X hold154/X _3975_/S VGND VPWR _3971_/X VGND VPWR sky130_fd_sc_hd__mux2_8
X_5710_ _7012_/Q _5630_/X _5645_/X _7028_/Q _5709_/X VGND VPWR _5711_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6690_ _6714_/CLK _6690_/D fanout470/X VGND VPWR _6690_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5641_ _5641_/A _5641_/B _5641_/C VGND VPWR _5670_/A VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_148_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5572_ _7093_/Q _7092_/Q VGND VPWR _5667_/B VGND VPWR sky130_fd_sc_hd__and2_2
Xclkbuf_1_0_1_csclk clkbuf_1_0_1_csclk/A VGND VPWR clkbuf_2_1_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_191_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4523_ _4584_/A _5042_/B VGND VPWR _4523_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_144_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold203 _3284_/X VGND VPWR _3285_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _4025_/X VGND VPWR _6464_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _6789_/Q VGND VPWR hold225/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _5495_/X VGND VPWR _7038_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _4454_/A _4626_/B VGND VPWR _4947_/C VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_132_616 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold247 _6419_/Q VGND VPWR hold247/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold258 _5204_/X VGND VPWR _6779_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _6681_/Q VGND VPWR hold269/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ input51/X _4058_/S _5337_/A _6905_/Q _3404_/X VGND VPWR _3408_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_7173_ _7173_/A VGND VPWR _7173_/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4385_ _4556_/A _4753_/A _4607_/A VGND VPWR _4441_/B VGND VPWR sky130_fd_sc_hd__and3_4
X_6124_ _7060_/Q _5954_/X _5976_/D _6879_/Q _6106_/X VGND VPWR _6125_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3336_ hold26/X hold46/X VGND VPWR _3415_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_682 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6055_ _7005_/Q _5958_/X _5978_/X _6997_/Q VGND VPWR _6055_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3267_ _3868_/A1 _3265_/X _3870_/S _3251_/A VGND VPWR _7158_/D VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_100_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5006_ _5006_/A _5112_/A VGND VPWR _5006_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_54_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3198_ _6989_/Q VGND VPWR _3198_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA_109 _3959_/B VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_26_335 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6957_ _6997_/CLK _6957_/D fanout463/X VGND VPWR _6957_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_157_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5908_ _5552_/B _7116_/Q _6103_/B1 VGND VPWR _5908_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_179_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6888_ _6888_/CLK _6888_/D fanout473/X VGND VPWR _6888_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5839_ _6685_/Q _5632_/X _5835_/X _5838_/X VGND VPWR _5839_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_10_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_741 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold770 _6429_/Q VGND VPWR hold770/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 _5280_/X VGND VPWR _6847_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _7186_/A VGND VPWR hold792/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_20 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_416 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_600 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1470 _7107_/Q VGND VPWR _5713_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _6575_/Q VGND VPWR _4169_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 _6053_/X VGND VPWR _7121_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_95 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput308 _3957_/X VGND VPWR spi_sdi VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_5_751 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput319 hold1345/X VGND VPWR hold1346/A VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_126_487 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_638 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4170_ _3447_/Y _4170_/A1 _4171_/S VGND VPWR _6576_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_750 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6811_ _7080_/CLK _6811_/D fanout479/X VGND VPWR _6811_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6742_ _6746_/CLK _6742_/D _3946_/B VGND VPWR _6742_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3954_ _3954_/A _3961_/B VGND VPWR _6638_/D VGND VPWR sky130_fd_sc_hd__and2_1
X_6673_ _6674_/CLK _6673_/D fanout468/X VGND VPWR _6673_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3885_ _5552_/B _5606_/A VGND VPWR _3885_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_31_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5624_ _5638_/A _5658_/B _5663_/C VGND VPWR _5624_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_176_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5555_ _7088_/Q _5562_/D VGND VPWR _5555_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4506_ _4469_/A _4887_/A _4672_/A _4846_/A _4672_/B VGND VPWR _4508_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
X_5486_ hold503/X _5528_/A1 hold50/X VGND VPWR _5486_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4437_ _4739_/A _4642_/A VGND VPWR _4635_/B VGND VPWR sky130_fd_sc_hd__nor2_8
X_7156_ _3945_/A1 _7156_/D _6387_/X VGND VPWR hold15/A VGND VPWR sky130_fd_sc_hd__dfrtn_1
XFILLER_86_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4368_ _4500_/A _4469_/A _6644_/Q VGND VPWR _5023_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_59_736 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6107_ _6863_/Q _5943_/X _5981_/X _6919_/Q VGND VPWR _6107_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3319_ _3453_/A hold64/X VGND VPWR _3454_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_59_769 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7087_ _7131_/CLK _7087_/D fanout460/X VGND VPWR _7087_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4299_ _4299_/A0 hold667/X _4303_/S VGND VPWR _4299_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6038_ _6924_/Q _5938_/X _5952_/X _6956_/Q VGND VPWR _6038_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XPHY_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_500 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_64_csclk _6447_/CLK VGND VPWR _7049_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_10_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_32 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_251 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_79_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6735_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_89_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VPWR _7079_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_122_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3670_ _3670_/A _3670_/B _3670_/C _3670_/D VGND VPWR _3670_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_185_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5340_ hold862/X _5484_/A1 _5345_/S VGND VPWR _5340_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5271_ hold704/X _5469_/A1 _5273_/S VGND VPWR _5271_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_141_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7010_ _7049_/CLK _7010_/D fanout457/X VGND VPWR _7010_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_4222_ hold273/X _5534_/A1 _4225_/S VGND VPWR _4222_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4153_ _4153_/A0 _5492_/A1 _4156_/S VGND VPWR _4153_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4084_ hold986/X _4083_/X _4084_/S VGND VPWR _4084_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4986_ _5005_/B _4985_/Y _4229_/X VGND VPWR _4986_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_6725_ _7140_/CLK _6725_/D _6307_/B VGND VPWR _6725_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3937_ _6516_/Q _3937_/A1 _6765_/Q VGND VPWR _3937_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_177_652 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6656_ _6659_/CLK _6656_/D fanout469/X VGND VPWR _6656_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3868_ _6406_/Q _3868_/A1 _3868_/S VGND VPWR _6406_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_149_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5607_ _5607_/A1 _5606_/B _5606_/Y _5552_/B VGND VPWR _7104_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6587_ _7137_/CLK _6587_/D VGND VPWR _6587_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_164_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3799_ _6737_/Q _5148_/A hold67/A _6465_/Q VGND VPWR _3799_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5538_ hold411/X _5538_/A1 _5540_/S VGND VPWR _5538_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_435 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5469_ hold656/X _5469_/A1 _5471_/S VGND VPWR _5469_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_457 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7139_ _7140_/CLK _7139_/D VGND VPWR _7139_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
Xfanout398 hold42/X VGND VPWR _5469_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_86_374 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xinput18 mask_rev_in[22] VGND VPWR input18/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_128_549 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput29 mask_rev_in[3] VGND VPWR input29/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_316 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_374 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4840_ _5051_/B _4911_/B VGND VPWR _5086_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_60_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_639 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4771_ _4771_/A _4995_/A _4771_/C _4771_/D VGND VPWR _4772_/D VGND VPWR sky130_fd_sc_hd__and4_1
X_6510_ _6951_/CLK _6510_/D fanout473/X VGND VPWR _6510_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_174_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3722_ _6907_/Q _5346_/A _4058_/S input44/X _3721_/X VGND VPWR _3729_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6441_ _6747_/CLK _6441_/D fanout449/X VGND VPWR _6441_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3653_ _6860_/Q _5292_/A _4151_/A _6562_/Q _3652_/X VGND VPWR _3661_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6372_ _6400_/A _6400_/B VGND VPWR _6372_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3584_ _3583_/X _6731_/Q _3829_/B VGND VPWR _6731_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_5323_ hold896/X _5509_/A1 _5327_/S VGND VPWR _5323_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5254_ hold714/X _5521_/A1 _5255_/S VGND VPWR _5254_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4205_ hold936/X _6355_/A1 _4207_/S VGND VPWR _4205_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5185_ _6353_/A1 _5185_/A1 _5185_/S VGND VPWR _5185_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clkbuf_3_7_0_csclk/A VGND VPWR _6888_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_4136_ hold866/X _5493_/A1 _4138_/S VGND VPWR _4136_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4067_ hold732/X _4066_/X _4067_/S VGND VPWR _4067_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_274 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4969_ _4969_/A _4969_/B VGND VPWR _4969_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_11_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6708_ _6709_/CLK _6708_/D fanout445/X VGND VPWR _6708_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_20_672 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6639_ _3937_/A1 _6639_/D fanout487/X VGND VPWR _6639_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_192_452 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_42 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_558 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6990_ _6990_/CLK _6990_/D fanout480/X VGND VPWR _6990_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_93_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5941_ _5968_/A _5964_/A _5969_/C VGND VPWR _5973_/A VGND VPWR sky130_fd_sc_hd__and3_4
X_5872_ _7036_/Q _5614_/X _5871_/X VGND VPWR _5872_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_61_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_758 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4823_ _4823_/A _5099_/A VGND VPWR _4823_/X VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_147_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4754_ _4581_/B _4456_/Y _4611_/Y _4689_/B VGND VPWR _4768_/C VGND VPWR sky130_fd_sc_hd__o22a_1
X_3705_ _7056_/Q hold86/A _5436_/A _6987_/Q VGND VPWR _3705_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4685_ _4685_/A _5042_/B VGND VPWR _4964_/B VGND VPWR sky130_fd_sc_hd__nand2_2
XFILLER_146_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6424_ _6926_/CLK _6424_/D fanout457/X VGND VPWR _6424_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3636_ _3268_/C _4118_/B _4262_/A _6663_/Q _3635_/X VGND VPWR _3636_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6355_ hold980/X _6355_/A1 _6357_/S VGND VPWR _6355_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3567_ _3960_/B _3331_/Y _4316_/A _6709_/Q VGND VPWR _3567_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_108_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5306_ hold475/X _5528_/A1 _5309_/S VGND VPWR _5306_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_115_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6286_ _6454_/Q _5947_/X _5965_/X _6549_/Q _6285_/X VGND VPWR _6289_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_3498_ _6894_/Q _5328_/A _4220_/A _6623_/Q VGND VPWR _3498_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_130_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5237_ hold391/X _5540_/A1 _5237_/S VGND VPWR _5237_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5168_ hold271/X _5465_/A1 _5170_/S VGND VPWR _5168_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_631 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4119_ _4119_/A0 _5491_/A1 _4126_/S VGND VPWR _4119_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5099_ _5099_/A _5099_/B _5099_/C _5099_/D VGND VPWR _5099_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_56_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_425 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold7 hold7/A VGND VPWR hold7/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_491 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_152 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_463 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire360 _5906_/Y VGND VPWR wire360/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
X_4470_ _4702_/C _4471_/C VGND VPWR _4664_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold407 _6860_/Q VGND VPWR hold407/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold418 _5334_/X VGND VPWR _6895_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_135 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold429 _6903_/Q VGND VPWR hold429/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3421_ _6944_/Q _5382_/A _3372_/Y _6440_/Q _3420_/X VGND VPWR _3421_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6140_ _6140_/A _6140_/B _6140_/C VGND VPWR _6140_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_3352_ _3374_/A hold28/X VGND VPWR _5328_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6071_ _7066_/Q _5934_/X _5975_/B _6869_/Q _6070_/X VGND VPWR _6074_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3283_ hold202/X hold70/X VGND VPWR _3283_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
Xhold1107 _6462_/Q VGND VPWR _4023_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _5112_/B _5021_/X _5006_/Y VGND VPWR _5022_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
Xhold1118 _4271_/X VGND VPWR _6667_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 _6567_/Q VGND VPWR _4160_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_322 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6973_ _6990_/CLK _6973_/D fanout480/X VGND VPWR _6973_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_53_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5924_ _6699_/Q _5637_/X _5645_/X _6459_/Q VGND VPWR _5924_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5855_ _6656_/Q _5899_/B VGND VPWR _5855_/Y VGND VPWR sky130_fd_sc_hd__nand2b_1
X_4806_ _4504_/X _5039_/B VGND VPWR _4964_/C VGND VPWR sky130_fd_sc_hd__and2b_1
X_5786_ _7008_/Q _5625_/X _5783_/X _5785_/X VGND VPWR _5787_/C VGND VPWR sky130_fd_sc_hd__a211o_1
X_4737_ _4737_/A _4737_/B VGND VPWR _4738_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_119_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_316 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4668_ _4921_/A _4928_/A _4668_/C VGND VPWR _5002_/A VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_134_124 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_455 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6407_ _3568_/A1 _6407_/D _6363_/X VGND VPWR hold44/A VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3619_ _6740_/Q _5148_/A _4014_/A _6458_/Q _3618_/X VGND VPWR _3620_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold930 _6936_/Q VGND VPWR hold930/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _5335_/X VGND VPWR _6896_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _4563_/A _4396_/A _4598_/Y VGND VPWR _4739_/B VGND VPWR sky130_fd_sc_hd__a21oi_2
Xhold952 _6542_/Q VGND VPWR hold952/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold963 _4138_/X VGND VPWR _6549_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold974 _6634_/Q VGND VPWR hold974/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6338_ _6644_/Q _6338_/A2 _6338_/B1 _6643_/Q VGND VPWR _6338_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold985 _3993_/X VGND VPWR _6436_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold996 _5151_/X VGND VPWR _6739_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6269_ _6683_/Q _5934_/X _5975_/B _6617_/Q _6268_/X VGND VPWR _6275_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_588 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_csclk clkbuf_2_3_0_csclk/A VGND VPWR clkbuf_3_7_0_csclk/A VGND VPWR
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_716 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_214 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_453 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3970_ hold988/X _6355_/A1 _3980_/S VGND VPWR _3970_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_514 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5640_ _7010_/Q _5630_/X _5633_/X _5639_/X VGND VPWR _5641_/C VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_176_558 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5571_ _6508_/Q _5658_/B VGND VPWR _5576_/B VGND VPWR sky130_fd_sc_hd__nand2_1
X_4522_ _4522_/A _4522_/B _4522_/C _4522_/D VGND VPWR _4522_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_116_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold204 _3285_/X VGND VPWR hold204/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _7081_/Q VGND VPWR hold215/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 _5215_/X VGND VPWR _6789_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _4607_/A _4453_/B VGND VPWR _4886_/B VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold237 hold237/A VGND VPWR hold237/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold248 _3968_/X VGND VPWR _6419_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 _6995_/Q VGND VPWR hold259/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _6897_/Q _5328_/A _5247_/A _6825_/Q VGND VPWR _3404_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_132_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4384_ _4384_/A _4892_/A VGND VPWR _4907_/B VGND VPWR sky130_fd_sc_hd__nor2_1
X_6123_ _6815_/Q _5971_/B _5949_/X _6935_/Q _6122_/X VGND VPWR _6125_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3335_ _3370_/A _3573_/A VGND VPWR _5382_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_58_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6054_ _6861_/Q _5943_/X _5981_/X _6917_/Q VGND VPWR _6054_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_85_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3266_ _6415_/Q _3266_/B VGND VPWR _3870_/S VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_105_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5005_ _5068_/B _5005_/B _5069_/B VGND VPWR _5112_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_100_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3197_ _6997_/Q VGND VPWR _3197_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_81_420 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6956_ _6981_/CLK _6956_/D fanout463/X VGND VPWR _6956_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5907_ _3223_/Y _5651_/Y _5896_/Y wire360/X _5552_/B VGND VPWR _5907_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6887_ _6951_/CLK _6887_/D fanout474/X VGND VPWR _6887_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_139_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5838_ _7034_/Q _5614_/X _5836_/X _5837_/X VGND VPWR _5838_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_5769_ _6815_/Q _5667_/X _5764_/X _5765_/X _5768_/X VGND VPWR _5769_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
XFILLER_108_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold760 _6548_/Q VGND VPWR hold760/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold771 _3985_/X VGND VPWR _6429_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 _6703_/Q VGND VPWR hold782/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold793 _4063_/X VGND VPWR _6495_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_32 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_428 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1460 _3488_/X VGND VPWR _6732_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1471 _5693_/X VGND VPWR _7107_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1482 _7127_/Q VGND VPWR _6204_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 _7171_/Q VGND VPWR _3233_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_431 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xoutput309 _3952_/X VGND VPWR spimemio_flash_io0_di VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_763 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_306 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_499 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_691 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6810_ _7058_/CLK _6810_/D _6396_/A VGND VPWR _6810_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_50_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6741_ _6746_/CLK _6741_/D _3946_/B VGND VPWR _6741_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3953_ _6403_/Q _3953_/B VGND VPWR _3953_/X VGND VPWR sky130_fd_sc_hd__and2b_4
X_6672_ _6674_/CLK _6672_/D fanout468/X VGND VPWR _6672_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3884_ _3894_/B2 _3174_/Y _3883_/X VGND VPWR _6506_/D VGND VPWR sky130_fd_sc_hd__a21o_1
X_5623_ _7094_/Q _7095_/Q VGND VPWR _5663_/C VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_164_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5554_ _5562_/D VGND VPWR _5554_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4505_ _5010_/A _4972_/A VGND VPWR _4912_/A VGND VPWR sky130_fd_sc_hd__nand2_1
X_5485_ _5485_/A0 _5545_/A1 hold50/X VGND VPWR _5485_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4436_ _4631_/D _4633_/B VGND VPWR _4615_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_160_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7155_ _7155_/CLK _7155_/D fanout450/X VGND VPWR _7155_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4367_ _4562_/A _4690_/B VGND VPWR _4469_/A VGND VPWR sky130_fd_sc_hd__nand2_4
X_6106_ _7084_/Q _5976_/B _5971_/C _7044_/Q VGND VPWR _6106_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3318_ _3555_/A _3714_/A VGND VPWR _5292_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_7086_ _7086_/CLK hold23/X fanout483/X VGND VPWR _7086_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_86_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4298_ _4298_/A _4322_/B VGND VPWR _4303_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_112_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6037_ _6972_/Q _5947_/X _5965_/X _6796_/Q _6036_/X VGND VPWR _6040_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3249_ _3249_/A _3249_/B VGND VPWR _3250_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_86_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_472 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6939_ _6981_/CLK _6939_/D fanout463/X VGND VPWR _6939_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_csclk _3942_/X VGND VPWR clkbuf_0_csclk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_135_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold590 _7042_/Q VGND VPWR hold590/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_534 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_480 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_0_0_csclk clkbuf_0_csclk/X VGND VPWR clkbuf_1_0_1_csclk/A VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_18_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1290 _4281_/X VGND VPWR _6675_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_152 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5270_ hold166/X hold60/X _5273_/S VGND VPWR _5270_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4221_ _4221_/A0 hold667/X _4225_/S VGND VPWR _4221_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_87_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4152_ _4152_/A0 _6353_/A1 _4156_/S VGND VPWR _4152_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4083_ hold555/X _5513_/A1 _4083_/S VGND VPWR _4083_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4985_ _5068_/B _5069_/B _5008_/B _4985_/D VGND VPWR _4985_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_168_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6724_ _7150_/CLK _6724_/D _6307_/B VGND VPWR _6724_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3936_ _6517_/Q user_clock _6766_/Q VGND VPWR _3936_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_149_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_2_0_csclk clkbuf_3_3_0_csclk/A VGND VPWR _6447_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_8
X_6655_ _6655_/CLK _6655_/D fanout468/X VGND VPWR _6655_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_137_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3867_ _3867_/A _3867_/B VGND VPWR _3868_/S VGND VPWR sky130_fd_sc_hd__nor2_1
X_5606_ _5606_/A _5606_/B VGND VPWR _5606_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_6586_ _7137_/CLK _6586_/D VGND VPWR _6586_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3798_ _6434_/Q _3372_/Y _3511_/Y _3796_/X _3797_/X VGND VPWR _3798_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_118_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5537_ hold806/X _5546_/A1 _5540_/S VGND VPWR _5537_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5468_ hold131/X hold60/X _5471_/S VGND VPWR _5468_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_9 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4419_ _4556_/A _4563_/A VGND VPWR _4561_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_5399_ hold592/X _5513_/A1 _5399_/S VGND VPWR _5399_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7138_ _7140_/CLK _7138_/D VGND VPWR _7138_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_143_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_504 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout399 hold42/X VGND VPWR _5538_/A1 VGND VPWR sky130_fd_sc_hd__buf_6
X_7069_ _7069_/CLK _7069_/D fanout482/X VGND VPWR _7069_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_100_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_386 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_428 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xinput19 mask_rev_in[23] VGND VPWR input19/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_10_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_586 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_710 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_272 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4770_ _4942_/C _4770_/B _5003_/A _4770_/D VGND VPWR _4771_/D VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_158_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3721_ _6899_/Q _5337_/A _5166_/A _6752_/Q VGND VPWR _3721_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6440_ _6747_/CLK _6440_/D fanout447/X VGND VPWR _6440_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_174_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3652_ _6657_/Q _4256_/A _4214_/A _6616_/Q VGND VPWR _3652_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_127_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6371_ _6400_/A _6400_/B VGND VPWR _6371_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3583_ _4192_/A0 _3642_/A1 _3829_/A VGND VPWR _3583_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5322_ _5322_/A0 _5484_/A1 _5327_/S VGND VPWR _5322_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5253_ hold800/X _5538_/A1 _5255_/S VGND VPWR _5253_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4204_ hold822/X _6354_/A1 _4207_/S VGND VPWR _4204_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5184_ _5184_/A _6352_/B VGND VPWR _5185_/S VGND VPWR sky130_fd_sc_hd__nand2_1
X_4135_ _4135_/A0 _5492_/A1 _4138_/S VGND VPWR _4135_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_63_csclk _6447_/CLK VGND VPWR _7011_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4066_ _4117_/A0 _5540_/A1 hold37/X VGND VPWR _4066_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_113_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6739_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4968_ _4627_/A _5041_/A _4789_/X VGND VPWR _5021_/B VGND VPWR sky130_fd_sc_hd__o21a_1
X_6707_ _6707_/CLK _6707_/D fanout445/X VGND VPWR _6707_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3919_ _6522_/Q input89/X _3921_/S VGND VPWR _3919_/X VGND VPWR sky130_fd_sc_hd__mux2_2
XFILLER_20_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4899_ _4899_/A _4899_/B _4877_/A VGND VPWR _5118_/A VGND VPWR sky130_fd_sc_hd__nor3b_1
XFILLER_177_494 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6638_ _7150_/CLK _6638_/D fanout487/X VGND VPWR _6638_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_137_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6569_ _6653_/CLK _6569_/D fanout454/X VGND VPWR _6569_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_767 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VPWR _7058_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_121_704 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_659 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_553 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5940_ _5964_/A _5981_/A _5981_/C VGND VPWR _5940_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_92_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5871_ _6717_/Q _5642_/X _5666_/X _6632_/Q VGND VPWR _5871_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4822_ _5084_/B _4942_/A VGND VPWR _5092_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_33_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4753_ _4753_/A _4753_/B _4753_/C VGND VPWR _5062_/C VGND VPWR sky130_fd_sc_hd__nand3_1
X_3704_ _6666_/Q _4268_/A _4316_/A _6706_/Q _3703_/X VGND VPWR _3709_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4684_ _4482_/A _4672_/A _4626_/Y _4230_/B VGND VPWR _4964_/A VGND VPWR sky130_fd_sc_hd__o31a_1
X_6423_ _7049_/CLK _6423_/D fanout457/X VGND VPWR _6423_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_147_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3635_ _7074_/Q _5532_/A _4202_/A _6607_/Q VGND VPWR _3635_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_127_380 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6354_ hold836/X _6354_/A1 _6357_/S VGND VPWR _6354_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3566_ _3573_/A hold66/X VGND VPWR _4316_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_115_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5305_ _5305_/A0 _5545_/A1 _5309_/S VGND VPWR _5305_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_103_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6285_ _6634_/Q _5946_/X _5955_/X _6554_/Q VGND VPWR _6285_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3497_ _3554_/A _3571_/B VGND VPWR _4220_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5236_ hold908/X _5548_/A1 _5237_/S VGND VPWR _5236_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_69_651 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5167_ _5167_/A0 _5524_/A1 _5170_/S VGND VPWR _5167_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4118_ _6400_/B _4118_/B _6352_/B VGND VPWR _4126_/S VGND VPWR sky130_fd_sc_hd__and3b_4
XFILLER_110_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5098_ _4810_/A _4582_/Y _4616_/Y _4626_/Y _4658_/C VGND VPWR _5099_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_83_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_518 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4049_ hold539/X _6357_/A1 _4049_/S VGND VPWR _4049_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_751 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_77 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold8 hold8/A VGND VPWR hold8/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_632 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_570 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire350 _3661_/Y VGND VPWR _3700_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_144_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire372 _3554_/A VGND VPWR _3374_/A VGND VPWR sky130_fd_sc_hd__buf_12
Xhold408 _5295_/X VGND VPWR _6860_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 _7073_/Q VGND VPWR hold419/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _7085_/Q _5541_/A hold76/A _7045_/Q VGND VPWR _3420_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_143_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3351_ _3586_/A _3573_/A VGND VPWR _5427_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6070_ _7050_/Q _5971_/A _5979_/X _6989_/Q VGND VPWR _6070_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3282_ hold47/X _3313_/A VGND VPWR _3586_/A VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold1108 _4023_/X VGND VPWR _6462_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5021_ _5021_/A _5021_/B _5021_/C _5021_/D VGND VPWR _5021_/X VGND VPWR sky130_fd_sc_hd__and4_1
Xhold1119 _7036_/Q VGND VPWR _5493_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6972_ _7080_/CLK _6972_/D fanout479/X VGND VPWR _6972_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_53_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5923_ _6608_/Q _5648_/X _5910_/X _5922_/X VGND VPWR _5923_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_179_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5854_ _6706_/Q _5638_/X _5654_/X _6676_/Q _5853_/X VGND VPWR _5862_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4805_ _4690_/A _4741_/A _4601_/B _4791_/X _4804_/X VGND VPWR _4805_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_5785_ _6904_/Q _5621_/X _5645_/X _7032_/Q _5784_/X VGND VPWR _5785_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_166_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4736_ _5010_/B _4644_/B _4735_/X _4921_/A VGND VPWR _4737_/B VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_162_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4667_ _4739_/B _4733_/B _4747_/B VGND VPWR _4668_/C VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_107_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6406_ _3945_/A1 _6406_/D _6362_/X VGND VPWR _6406_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_134_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold920 _6816_/Q VGND VPWR hold920/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ _6989_/Q _5436_/A _5463_/A _7013_/Q VGND VPWR _3618_/X VGND VPWR sky130_fd_sc_hd__a22o_2
Xhold931 _5380_/X VGND VPWR _6936_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4598_ _4642_/A _5043_/A VGND VPWR _4598_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold942 _6603_/Q VGND VPWR hold942/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_606 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold953 _4130_/X VGND VPWR _6542_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _6674_/Q VGND VPWR hold964/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6337_ _6336_/X _6337_/A1 _6346_/S VGND VPWR _7145_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold975 _4243_/X VGND VPWR _6634_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ _6822_/Q _5247_/A hold49/A _7030_/Q VGND VPWR _3549_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_1_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold986 _7178_/A VGND VPWR hold986/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold997 _7184_/A VGND VPWR hold997/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6268_ _6703_/Q _5971_/A _5979_/X _6473_/Q VGND VPWR _6268_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_88_267 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5219_ hold660/X _5513_/A1 hold18/X VGND VPWR _5219_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6199_ _6690_/Q _5954_/X _5976_/D _6619_/Q _6180_/X VGND VPWR _6200_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_151_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_573 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_61 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_434 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_226 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5570_ _7093_/Q _7092_/Q VGND VPWR _5658_/B VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_191_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4521_ _4584_/A _4531_/B VGND VPWR _4522_/D VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold205 _3286_/X VGND VPWR _3347_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 _5544_/X VGND VPWR _7081_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4452_ _4753_/A _4454_/A VGND VPWR _4453_/B VGND VPWR sky130_fd_sc_hd__nand2b_4
Xhold227 _6669_/Q VGND VPWR hold227/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _4105_/X VGND VPWR _6520_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold249 _6955_/Q VGND VPWR hold249/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3403_ _6977_/Q _5418_/A _3381_/Y input33/X _3402_/X VGND VPWR _3408_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_171_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7171_ _3945_/A1 _7171_/D _6401_/X VGND VPWR _7171_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4383_ _4892_/A VGND VPWR _4462_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6122_ _6447_/Q _5601_/X _5959_/X _6967_/Q VGND VPWR _6122_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3334_ _3571_/A _3370_/A VGND VPWR _5238_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_58_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6053_ _6053_/A0 _6052_/X _6279_/S VGND VPWR _6053_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3265_ _7159_/Q _6415_/Q _3266_/B VGND VPWR _3265_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_5004_ _5004_/A _5004_/B _5074_/B _5071_/B VGND VPWR _5004_/Y VGND VPWR sky130_fd_sc_hd__nand4_1
X_3196_ _7005_/Q VGND VPWR _3196_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_451 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6955_ _7012_/CLK _6955_/D fanout458/X VGND VPWR _6955_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5906_ _5906_/A _5906_/B _5906_/C _5906_/D VGND VPWR _5906_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_62_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6886_ _6890_/CLK _6886_/D fanout476/X VGND VPWR _6886_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_167_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5837_ _6650_/Q _5646_/X _5667_/X _6555_/Q VGND VPWR _5837_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_179_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5768_ _6447_/Q _5614_/X _5766_/X _5767_/X VGND VPWR _5768_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_108_604 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_529 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4719_ _4469_/A _4639_/Y _4673_/B _4694_/Y VGND VPWR _4719_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_108_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5699_ _6868_/Q _5628_/X _5634_/X _6972_/Q _5698_/X VGND VPWR _5706_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_478 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold750 _7016_/Q VGND VPWR hold750/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold761 _4137_/X VGND VPWR _6548_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _6437_/Q VGND VPWR hold772/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _4314_/X VGND VPWR _6703_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _6686_/Q VGND VPWR hold794/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_161 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1450 _3313_/A VGND VPWR _3375_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _6733_/Q VGND VPWR _3449_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 _6576_/Q VGND VPWR _4170_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1483 _7125_/Q VGND VPWR _6178_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1494 _6571_/Q VGND VPWR _4165_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_443 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_98 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_318 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_194 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_432 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6740_ _6746_/CLK _6740_/D _3946_/B VGND VPWR _6740_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3952_ _6404_/Q _3952_/B VGND VPWR _3952_/X VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_189_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6671_ _6671_/CLK _6671_/D fanout468/X VGND VPWR _6671_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3883_ _7088_/Q _7089_/Q _6509_/Q _5608_/C VGND VPWR _3883_/X VGND VPWR sky130_fd_sc_hd__and4b_1
X_5622_ _7018_/Q _5619_/X _5621_/X _6898_/Q _5617_/X VGND VPWR _5641_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5553_ _6509_/Q _5552_/B _6508_/Q _3885_/Y VGND VPWR _5562_/D VGND VPWR sky130_fd_sc_hd__o31a_1
XFILLER_191_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_754 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4504_ _4969_/A _4984_/A _4965_/B VGND VPWR _4504_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_5484_ hold878/X _5484_/A1 hold50/X VGND VPWR _5484_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4435_ _4566_/A _4591_/A VGND VPWR _4482_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_132_437 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7154_ _7155_/CLK _7154_/D fanout449/X VGND VPWR _7154_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4366_ _4690_/A _4460_/A VGND VPWR _5010_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_113_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6105_ _7068_/Q _5934_/X _5975_/B _6871_/Q VGND VPWR _6105_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3317_ hold27/X hold84/X VGND VPWR _3714_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7085_ _7085_/CLK _7085_/D fanout483/X VGND VPWR _7085_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4297_ hold531/X _6357_/A1 _4297_/S VGND VPWR _4297_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6036_ _6892_/Q _5946_/X _5955_/X _6804_/Q VGND VPWR _6036_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3248_ _3248_/A1 _3249_/B _3247_/Y _7168_/Q VGND VPWR _3248_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_100_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_484 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3179_ _6508_/Q VGND VPWR _5610_/B VGND VPWR sky130_fd_sc_hd__clkinv_2
XPHY_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7026_/CLK _6938_/D fanout463/X VGND VPWR _6938_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XPHY_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6869_ _7085_/CLK _6869_/D fanout477/X VGND VPWR _6869_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_50_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold580 _6709_/Q VGND VPWR hold580/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 _5500_/X VGND VPWR _7042_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_88 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_492 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1280 _4021_/X VGND VPWR _6460_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 _6560_/Q VGND VPWR _4152_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_373 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_201 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_286 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4220_ _4220_/A _4322_/B VGND VPWR _4225_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_4151_ _4151_/A _4322_/B VGND VPWR _4156_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_95_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4082_ hold239/X _4081_/X _4084_/S VGND VPWR _4082_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_593 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4984_ _4984_/A _4984_/B VGND VPWR _4997_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_177_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6723_ _7150_/CLK _6723_/D _6307_/B VGND VPWR _6723_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3935_ _3222_/Y input2/X input1/X VGND VPWR _3935_/X VGND VPWR sky130_fd_sc_hd__mux2_4
X_6654_ _6654_/CLK hold61/X fanout454/X VGND VPWR _6654_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3866_ _3865_/X _3866_/A1 _3866_/S VGND VPWR _6407_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_137_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5605_ _5552_/Y _5567_/Y _5604_/Y _6509_/Q VGND VPWR _5606_/B VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_176_175 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6585_ _7137_/CLK _6585_/D VGND VPWR _6585_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3797_ _6882_/Q _5319_/A _4238_/A _6630_/Q VGND VPWR _3797_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_11_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_540 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5536_ _5536_/A0 _5545_/A1 _5540_/S VGND VPWR _5536_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5467_ _5467_/A0 _5545_/A1 _5471_/S VGND VPWR _5467_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4418_ _4556_/A _4563_/A VGND VPWR _4600_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_5398_ hold636/X _5521_/A1 _5399_/S VGND VPWR _5398_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7137_ _7137_/CLK _7137_/D VGND VPWR _7137_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_4349_ _4471_/B _4591_/A VGND VPWR _4911_/A VGND VPWR sky130_fd_sc_hd__and2b_2
XFILLER_86_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xfanout389 _4546_/Y VGND VPWR _4846_/B VGND VPWR sky130_fd_sc_hd__buf_6
X_7068_ _7078_/CLK _7068_/D fanout482/X VGND VPWR _7068_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_143_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_175 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6019_ _7064_/Q _5934_/X _5975_/B _6867_/Q _6018_/X VGND VPWR _6024_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_100_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_418 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_598 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_402 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_610 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3720_ _3720_/A _3720_/B _3720_/C _3720_/D VGND VPWR _3730_/B VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_9_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3651_ _3651_/A _3651_/B _3651_/C _3651_/D VGND VPWR _3651_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_158_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6370_ _6383_/A _6396_/B VGND VPWR _6370_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3582_ _3582_/A _3582_/B _3582_/C VGND VPWR _3582_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
XFILLER_127_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5321_ hold535/X _5543_/A1 _5327_/S VGND VPWR _5321_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5252_ hold188/X _5519_/A1 _5255_/S VGND VPWR _5252_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_727 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4203_ _4203_/A0 _5491_/A1 _4207_/S VGND VPWR _4203_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5183_ hold17/X _5183_/B VGND VPWR _5183_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_4134_ _4134_/A0 _5491_/A1 _4138_/S VGND VPWR _4134_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4065_ _4065_/A0 _4064_/X _4067_/S VGND VPWR _4065_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4967_ _4967_/A _4967_/B VGND VPWR _5066_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_3918_ _6523_/Q input91/X _3921_/S VGND VPWR _3918_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_6706_ _6709_/CLK _6706_/D fanout445/X VGND VPWR _6706_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4898_ _4359_/Y _4892_/B _4877_/C VGND VPWR _4899_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_149_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6637_ _7150_/CLK _6637_/D fanout487/X VGND VPWR _6637_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3849_ _3849_/A1 _3851_/C _3848_/X _3292_/X VGND VPWR _6413_/D VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_20_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_465 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6568_ _6755_/CLK _6568_/D fanout445/X VGND VPWR _6568_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_98_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5519_ hold178/X _5519_/A1 hold87/A VGND VPWR _5519_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6499_ _6755_/CLK _6499_/D _6360_/A VGND VPWR _6499_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_133_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_145 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_540 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_476 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_565 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_90 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5870_ _6477_/Q _5630_/X _5867_/X _5868_/X _5869_/X VGND VPWR _5870_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_61_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4821_ _4542_/A _4562_/Y _4518_/B VGND VPWR _4821_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_61_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4752_ _4413_/Y _4672_/B _4619_/Y _4626_/Y VGND VPWR _4995_/A VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_147_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3703_ _6461_/Q _4020_/A _4014_/A _6456_/Q VGND VPWR _3703_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_119_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4683_ _4424_/Y _4430_/Y _4504_/X _4682_/Y _4920_/B VGND VPWR _4683_/X VGND VPWR
+ sky130_fd_sc_hd__o41a_1
X_6422_ _6749_/CLK _6422_/D fanout449/X VGND VPWR _6422_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3634_ _6973_/Q _5418_/A _5364_/A _6925_/Q _3633_/X VGND VPWR _3638_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_2
X_6353_ _6353_/A0 _6353_/A1 _6357_/S VGND VPWR _6353_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3565_ _3565_/A _3565_/B _3565_/C VGND VPWR _3581_/C VGND VPWR sky130_fd_sc_hd__nor3_1
X_5304_ hold966/X _5484_/A1 _5309_/S VGND VPWR _5304_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6284_ _6689_/Q _5961_/X _6282_/X _6283_/X VGND VPWR _6289_/A VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_0_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3496_ _6757_/Q _5182_/S _4310_/A _6704_/Q _3494_/X VGND VPWR _3504_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_130_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5235_ hold511/X _5538_/A1 _5237_/S VGND VPWR _5235_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5166_ _5166_/A hold17/X VGND VPWR _5170_/S VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_68_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4117_ _4117_/A0 hold22/X hold38/X VGND VPWR hold39/A VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_549 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5097_ _5115_/A _5087_/Y _5096_/X _5078_/X VGND VPWR _6724_/D VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_83_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4048_ hold774/X _6356_/A1 _4049_/S VGND VPWR _4048_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5999_ _6802_/Q _5955_/X _5975_/B _6866_/Q _5983_/X VGND VPWR _6000_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XPHY_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput290 _6437_/Q VGND VPWR pll_trim[3] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_58_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold9 hold9/A VGND VPWR hold9/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_74_110 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_644 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_224 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_270 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_112 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire351 _3651_/Y VGND VPWR _3700_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_62_csclk _6447_/CLK VGND VPWR _6963_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_156_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold409 _7057_/Q VGND VPWR hold409/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3350_ hold48/X _3543_/A VGND VPWR _5409_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_97_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_77_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6746_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_3281_ hold83/X hold64/X VGND VPWR _3313_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_151_192 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5020_ _5021_/A _5021_/B _5021_/D VGND VPWR _5135_/A VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1109 _6965_/Q VGND VPWR _5413_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_493 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6971_ _7080_/CLK _6971_/D fanout480/X VGND VPWR _6971_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_5922_ _6649_/Q _5621_/X _5654_/X _6679_/Q _5921_/X VGND VPWR _5922_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_15_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6712_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5853_ _7152_/Q _5625_/X _5666_/X _6631_/Q VGND VPWR _5853_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_167_708 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4804_ _4804_/A _4804_/B _4804_/C VGND VPWR _4804_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_5784_ _6944_/Q _5632_/X _5664_/X _6928_/Q VGND VPWR _5784_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_9_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4735_ _4735_/A _4735_/B _4747_/C VGND VPWR _4735_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_119_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4666_ _4441_/A _4400_/B _4665_/X VGND VPWR _4733_/B VGND VPWR sky130_fd_sc_hd__o21ai_1
X_6405_ _3945_/A1 _6405_/D _6361_/X VGND VPWR _6405_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3617_ _6949_/Q _3781_/A2 _4280_/A _6678_/Q _3616_/X VGND VPWR _3620_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold910 _7045_/Q VGND VPWR hold910/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _5245_/X VGND VPWR _6816_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _4735_/B _4735_/A VGND VPWR _4747_/B VGND VPWR sky130_fd_sc_hd__and2b_1
Xhold932 _6904_/Q VGND VPWR hold932/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _4201_/X VGND VPWR _6603_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 _6707_/Q VGND VPWR hold954/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _6642_/Q _6336_/A2 _6336_/B1 _6350_/A2 _6335_/X VGND VPWR _6336_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3548_ input24/X _3367_/Y _5463_/A _7014_/Q _3547_/X VGND VPWR _3552_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold965 _4279_/X VGND VPWR _6674_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _6599_/Q VGND VPWR hold976/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _4084_/X VGND VPWR _6505_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _4059_/X VGND VPWR _6493_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ _6563_/Q _5953_/X _5960_/X _6673_/Q _6266_/X VGND VPWR _6267_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3479_ _6807_/Q _5229_/A _5301_/A _6871_/Q _3478_/X VGND VPWR _3484_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5218_ hold139/X hold99/X hold18/X VGND VPWR _5218_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_88_279 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6198_ _6555_/Q _5971_/B _5949_/X _6675_/Q _6197_/X VGND VPWR _6200_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5149_ _5149_/A0 _5491_/A1 _5153_/S VGND VPWR _5149_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_151_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_699 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_410 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_487 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_719 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4520_ _4724_/A _4953_/A VGND VPWR _4522_/C VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_172_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4451_ _4753_/A _4495_/A VGND VPWR _4496_/B VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_172_744 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold206 _3370_/Y VGND VPWR _5454_/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 _6941_/Q VGND VPWR hold217/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _4273_/X VGND VPWR _6669_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold239 _6504_/Q VGND VPWR hold239/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ _6961_/Q _5400_/A _5256_/A _6833_/Q VGND VPWR _3402_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_7170_ _3927_/A1 _7170_/D _6400_/X VGND VPWR _7170_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4382_ _4359_/B _4382_/B VGND VPWR _4892_/A VGND VPWR sky130_fd_sc_hd__nand2b_2
XFILLER_124_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6121_ _7031_/Q _5944_/X _5975_/A _6847_/Q _6120_/X VGND VPWR _6125_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3333_ hold85/X hold75/X VGND VPWR _5445_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_112_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6052_ _7120_/Q _6051_/X _6303_/S VGND VPWR _6052_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3264_ _6485_/Q _3264_/B VGND VPWR _3266_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_39_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5003_ _5003_/A _5003_/B _5003_/C VGND VPWR _5071_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_3195_ _7013_/Q VGND VPWR _3195_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_463 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6954_ _7012_/CLK _6954_/D fanout458/X VGND VPWR _6954_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5905_ _6548_/Q _5905_/A2 _5666_/X _6633_/Q _5904_/X VGND VPWR _5906_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6885_ _6969_/CLK _6885_/D fanout475/X VGND VPWR _6885_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_22_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5836_ _6715_/Q _5642_/X _5666_/X _6630_/Q VGND VPWR _5836_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_167_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5767_ _6999_/Q _5643_/X _5664_/X _6927_/Q VGND VPWR _5767_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4718_ _4645_/Y _4690_/Y _4716_/Y _4717_/X VGND VPWR _4721_/B VGND VPWR sky130_fd_sc_hd__o211a_1
X_5698_ _6980_/Q _5624_/X _5654_/X _6932_/Q VGND VPWR _5698_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4649_ _4612_/Y _4613_/Y _4616_/Y _4609_/Y _4621_/X VGND VPWR _4660_/A VGND VPWR
+ sky130_fd_sc_hd__o221a_1
Xhold740 _6708_/Q VGND VPWR hold740/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _5470_/X VGND VPWR _7016_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _6817_/Q VGND VPWR hold762/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold773 _3994_/X VGND VPWR _6437_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _6421_/Q VGND VPWR hold784/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _6320_/B _6319_/B VGND VPWR _6319_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold795 _4294_/X VGND VPWR _6686_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1440 _6591_/Q VGND VPWR _4188_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 _3814_/B VGND VPWR _3376_/B VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1462 _6721_/Q VGND VPWR _4885_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1473 _6572_/Q VGND VPWR _4166_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1484 _6154_/X VGND VPWR _7125_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1495 _6589_/Q VGND VPWR _4185_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_541 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3951_ input85/X _3251_/A _6404_/Q VGND VPWR _3951_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_6670_ _6671_/CLK _6670_/D fanout468/X VGND VPWR _6670_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_149_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3882_ _7090_/Q _7091_/Q VGND VPWR _5608_/C VGND VPWR sky130_fd_sc_hd__nor2_1
X_5621_ _5664_/A _5666_/B _5660_/C VGND VPWR _5621_/X VGND VPWR sky130_fd_sc_hd__and3b_4
X_5552_ _6509_/Q _5552_/B VGND VPWR _5552_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_4503_ _4582_/B _4881_/B VGND VPWR _4925_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_129_295 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5483_ hold588/X _5543_/A1 hold50/X VGND VPWR _5483_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4434_ _4566_/A _4434_/B VGND VPWR _4984_/A VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_104_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_736 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7153_ _7155_/CLK _7153_/D fanout449/X VGND VPWR _7153_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4365_ _4556_/A _4563_/A VGND VPWR _4460_/A VGND VPWR sky130_fd_sc_hd__nand2b_4
XFILLER_113_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6104_ _6103_/Y _6102_/X _6279_/S _6104_/B2 VGND VPWR _7123_/D VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3316_ hold27/X hold84/X VGND VPWR _5161_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_113_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7084_ _7086_/CLK hold43/X fanout482/X VGND VPWR _7084_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4296_ hold724/X _6356_/A1 _4297_/S VGND VPWR _4296_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_140_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6035_ _6940_/Q _5961_/X _6031_/X _6034_/X VGND VPWR _6040_/A VGND VPWR sky130_fd_sc_hd__a211o_1
X_3247_ _3249_/B _3250_/A VGND VPWR _3247_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_86_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_400 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3178_ _5552_/B VGND VPWR _3178_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6937_ _7086_/CLK _6937_/D fanout483/X VGND VPWR _6937_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6868_ _6882_/CLK _6868_/D fanout475/X VGND VPWR _6868_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_313 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5819_ _6793_/Q _5652_/Y _5811_/X _5818_/X _6303_/S VGND VPWR _5819_/X VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_6799_ _6888_/CLK _6799_/D fanout474/X VGND VPWR _6799_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_182_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold570 _6987_/Q VGND VPWR hold570/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _4321_/X VGND VPWR _6709_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _6953_/Q VGND VPWR hold592/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_614 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1270 _4239_/X VGND VPWR _6630_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1281 _6650_/Q VGND VPWR _4251_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 _4152_/X VGND VPWR _6560_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_363 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_700 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_563 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_574 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_127 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4150_ hold192/X _5519_/A1 _4150_/S VGND VPWR _4150_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4081_ _4125_/A0 hold99/X _4118_/B VGND VPWR _4081_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_666 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4983_ _5066_/A _4983_/B _4983_/C VGND VPWR _4985_/D VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_189_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6722_ _7150_/CLK _6722_/D fanout487/X VGND VPWR _6722_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3934_ _3221_/Y _7157_/Q _6400_/B VGND VPWR _3934_/X VGND VPWR sky130_fd_sc_hd__mux2_2
X_6653_ _6653_/CLK _6653_/D _6401_/A VGND VPWR _6653_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3865_ _3167_/Y _3251_/A _6488_/Q VGND VPWR _3865_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5604_ _5608_/C _5604_/B VGND VPWR _5604_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_118_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6584_ _7137_/CLK _6584_/D VGND VPWR _6584_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3796_ _6914_/Q _5355_/A _5541_/A _7079_/Q _3795_/X VGND VPWR _3796_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_733 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5535_ hold419/X _5544_/A1 _5540_/S VGND VPWR _5535_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5466_ hold353/X _5526_/A1 _5471_/S VGND VPWR _5466_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_427 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4417_ _4459_/B _4456_/A VGND VPWR _4542_/B VGND VPWR sky130_fd_sc_hd__nand2_4
X_5397_ hold786/X _5538_/A1 _5399_/S VGND VPWR _5397_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_683 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7136_ _7140_/CLK _7136_/D VGND VPWR _7136_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_4348_ _4376_/A _4376_/B VGND VPWR _4471_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_101_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_709 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7067_ _7067_/CLK _7067_/D fanout477/X VGND VPWR _7067_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4279_ hold964/X _5546_/A1 _4279_/S VGND VPWR _4279_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_46_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6018_ _7048_/Q _5971_/A _5979_/X _6987_/Q VGND VPWR _6018_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_55_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_74 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_699 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3650_ _6892_/Q _5328_/A _3981_/A _6428_/Q _3649_/X VGND VPWR _3651_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_530 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3581_ _3581_/A _3581_/B _3581_/C _3581_/D VGND VPWR _3582_/C VGND VPWR sky130_fd_sc_hd__and4_2
X_5320_ _5320_/A0 _5473_/A1 _5327_/S VGND VPWR _5320_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_127_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_213 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5251_ _5251_/A0 _5545_/A1 _5255_/S VGND VPWR _5251_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4202_ _4202_/A _6352_/B VGND VPWR _4207_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_130_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5182_ hold990/X _5524_/A1 _5182_/S VGND VPWR _5182_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4133_ _4133_/A _6352_/B VGND VPWR _4138_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_68_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4064_ hold900/X _5548_/A1 hold37/X VGND VPWR _4064_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4966_ _5088_/A _5114_/A _5088_/C VGND VPWR _5008_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_177_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6705_ _6707_/CLK _6705_/D fanout445/X VGND VPWR _6705_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3917_ _6487_/Q _3916_/Y _3829_/B VGND VPWR _7157_/D VGND VPWR sky130_fd_sc_hd__o21a_2
X_4897_ _4900_/B _4911_/C VGND VPWR _4899_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_149_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6636_ _7150_/CLK _6636_/D fanout487/X VGND VPWR _6636_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3848_ _3866_/S _3845_/S _3847_/X _3860_/B VGND VPWR _3848_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_164_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6567_ _6653_/CLK _6567_/D _6401_/A VGND VPWR _6567_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3779_ _6426_/Q _3981_/A _6352_/A _7151_/Q _3778_/X VGND VPWR _3782_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5518_ hold323/X _5518_/A1 hold87/A VGND VPWR _5518_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6498_ _6735_/CLK _6498_/D _3946_/B VGND VPWR _6498_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_145_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5449_ hold219/X _5494_/A1 _5453_/S VGND VPWR _5449_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_333 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7119_ _7126_/CLK _7119_/D fanout466/X VGND VPWR _7119_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_101_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_358 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VPWR _6347_/A1 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_63_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_602 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_552 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_488 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_330 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_577 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_96 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4820_ _4542_/A _4902_/A _4456_/Y _4562_/Y VGND VPWR _4820_/X VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_61_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4751_ _4581_/B _4948_/C _4611_/Y _4639_/Y VGND VPWR _4768_/B VGND VPWR sky130_fd_sc_hd__o22a_1
XFILLER_193_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3702_ _3701_/X _3702_/A1 _3829_/B VGND VPWR _6729_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_4682_ _4682_/A _4682_/B _4682_/C VGND VPWR _4682_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_119_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6421_ _6749_/CLK _6421_/D fanout449/X VGND VPWR _6421_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3633_ _6957_/Q _5400_/A _4008_/A _6453_/Q VGND VPWR _3633_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_146_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6352_ _6352_/A _6352_/B VGND VPWR _6357_/S VGND VPWR sky130_fd_sc_hd__and2_2
X_3564_ _6998_/Q _5445_/A _5238_/A _6814_/Q _3563_/X VGND VPWR _3565_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5303_ hold551/X _5543_/A1 _5309_/S VGND VPWR _5303_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6283_ _6479_/Q _5940_/X _5967_/X _6608_/Q _6281_/X VGND VPWR _6283_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3495_ hold74/X _3814_/B VGND VPWR _4310_/A VGND VPWR sky130_fd_sc_hd__nor2_2
X_5234_ hold451/X _5528_/A1 _5237_/S VGND VPWR _5234_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5165_ _5165_/A0 _5524_/A1 _5165_/S VGND VPWR _5165_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4116_ hold900/X _5548_/A1 hold38/X VGND VPWR _4116_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5096_ _5122_/A _5096_/B _5096_/C VGND VPWR _5096_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_84_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4047_ hold934/X _6355_/A1 _4049_/S VGND VPWR _4047_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_542 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5998_ _6858_/Q _5943_/X _5952_/X _6954_/Q _5997_/X VGND VPWR _6000_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4949_ _4542_/A _4456_/Y _4948_/X _4946_/X VGND VPWR _4963_/A VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_33_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6619_ _6712_/CLK _6619_/D fanout470/X VGND VPWR _6619_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_165_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_352 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_374 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput280 _6420_/Q VGND VPWR pll_trim[18] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput291 _6438_/Q VGND VPWR pll_trim[4] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_87_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_715 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_282 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_472 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_124 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire352 _3611_/Y VGND VPWR _3640_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3280_ hold63/X _6723_/Q _3975_/S VGND VPWR hold64/A VGND VPWR sky130_fd_sc_hd__mux2_8
XFILLER_151_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_623 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_336 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6970_ _7063_/CLK _6970_/D fanout463/X VGND VPWR _6970_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5921_ _6464_/Q _5624_/X _5634_/X _6454_/Q _5911_/Y VGND VPWR _5921_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5852_ _5852_/A _5852_/B _5852_/C VGND VPWR _5852_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_61_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_726 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4803_ _5088_/A _5088_/C _4803_/C VGND VPWR _4804_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_21_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5783_ _6808_/Q _5660_/X _5667_/X _6816_/Q VGND VPWR _5783_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_166_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4734_ _4735_/A _4735_/B VGND VPWR _4740_/A VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_9_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_433 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4665_ _4563_/A _4642_/A _4441_/B _4739_/A VGND VPWR _4665_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_135_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6404_ _3927_/A1 _6404_/D _6360_/X VGND VPWR _6404_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_190_734 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold900 _6530_/Q VGND VPWR hold900/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ _6478_/Q _4038_/A _6352_/A _7154_/Q VGND VPWR _3616_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold911 _5503_/X VGND VPWR _7045_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 _6848_/Q VGND VPWR hold922/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4596_ _4627_/B _4562_/Y _4595_/A _4633_/B VGND VPWR _4735_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_1
Xhold933 _5344_/X VGND VPWR _6904_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _6554_/Q VGND VPWR hold944/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _6644_/Q _6335_/A2 _6335_/B1 _6643_/Q VGND VPWR _6335_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold955 _4319_/X VGND VPWR _6707_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3547_ _7051_/Q _5505_/A _4322_/A _6714_/Q VGND VPWR _3547_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold966 _6868_/Q VGND VPWR hold966/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _4197_/X VGND VPWR _6599_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold988 _6420_/Q VGND VPWR hold988/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 _6578_/Q VGND VPWR hold999/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _6653_/Q _5973_/A _5948_/X _6698_/Q _6265_/X VGND VPWR _6266_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3478_ _6959_/Q _5400_/A hold29/A hold56/A VGND VPWR _3478_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5217_ hold683/X _5469_/A1 hold18/X VGND VPWR _5217_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1600 _6535_/Q VGND VPWR hold243/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6197_ _7034_/Q _5601_/X _5959_/X _6715_/Q VGND VPWR _6197_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_192_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_472 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5148_ _5148_/A _6352_/B VGND VPWR _5153_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_57_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5079_ _4902_/A _4456_/Y _4689_/B _4691_/A _4872_/A VGND VPWR _5080_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_380 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_670 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_444 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_330 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_396 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_486 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_681 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_730 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_723 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_262 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4450_ _4902_/A _4948_/B _4442_/Y VGND VPWR _4450_/Y VGND VPWR sky130_fd_sc_hd__o21ai_1
XFILLER_156_296 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold207 _5461_/S VGND VPWR _5462_/S VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_447 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold218 _5386_/X VGND VPWR _6941_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _6679_/Q VGND VPWR hold229/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ _7062_/Q hold86/A _3981_/A _6433_/Q _3400_/X VGND VPWR _3408_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4381_ _4739_/A _4492_/D VGND VPWR _4381_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_6120_ hold56/A _5937_/X _5975_/D _6887_/Q VGND VPWR _6120_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3332_ _3347_/A hold73/X VGND VPWR hold74/A VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_124_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_344 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6051_ _6040_/Y _6050_/X _6788_/Q _6226_/B VGND VPWR _6051_/X VGND VPWR sky130_fd_sc_hd__o2bb2a_1
X_3263_ _3834_/B2 _3262_/Y _3261_/X VGND VPWR _7159_/D VGND VPWR sky130_fd_sc_hd__a21bo_1
XFILLER_98_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5002_ _5002_/A _5002_/B _5002_/C VGND VPWR _5074_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_3194_ _7021_/Q VGND VPWR _3194_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_53_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_486 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6953_ _6953_/CLK _6953_/D fanout460/X VGND VPWR _6953_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_53_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5904_ _6463_/Q _5624_/X _5664_/X _6668_/Q VGND VPWR _5904_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_34_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6884_ _6884_/CLK _6884_/D fanout477/X VGND VPWR _6884_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5835_ _6705_/Q _5638_/X _5834_/X VGND VPWR _5835_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_167_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5766_ _6823_/Q _5818_/A2 _5814_/B1 _6911_/Q VGND VPWR _5766_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4717_ _4482_/A _4672_/A _4902_/A _4476_/Y _4609_/Y VGND VPWR _4717_/X VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_175_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5697_ _6988_/Q _5627_/X _5635_/X _6828_/Q VGND VPWR _5697_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_30_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4648_ _4556_/A _4563_/A _4689_/B _5062_/A _4647_/X VGND VPWR _4648_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
XFILLER_123_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold730 _6607_/Q VGND VPWR hold730/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _4320_/X VGND VPWR _6708_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ _4579_/A _4579_/B VGND VPWR _4948_/D VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold752 _6521_/Q VGND VPWR hold752/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _5246_/X VGND VPWR _6817_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _6483_/Q VGND VPWR hold774/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6320_/B _6318_/B VGND VPWR _6318_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold785 _3972_/X VGND VPWR _6421_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _6476_/Q VGND VPWR hold796/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6249_ _7036_/Q _5601_/X _5959_/X _6717_/Q _6248_/X VGND VPWR _6250_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_420 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1430 _7136_/Q VGND VPWR _6311_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1441 _7134_/Q VGND VPWR _6309_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _3976_/X VGND VPWR _6423_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1463 _3303_/Y VGND VPWR hold27/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1474 _7139_/Q VGND VPWR _6314_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 _7129_/Q VGND VPWR _6278_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_61_csclk _6447_/CLK VGND VPWR _7017_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold1496 _6639_/Q VGND VPWR _3881_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_189_108 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_372 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_76_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6707_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_71_66 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_631 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_csclk clkbuf_3_5_0_csclk/X VGND VPWR _6629_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_136_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_431 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_401 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold90 hold90/A VGND VPWR hold90/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7080_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_91_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3950_ _3950_/A VGND VPWR _3950_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_90_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3881_ _6644_/Q _3962_/B _3881_/B1 VGND VPWR _6644_/D VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_149_528 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5620_ _7092_/Q _7093_/Q VGND VPWR _5660_/C VGND VPWR sky130_fd_sc_hd__and2b_2
X_5551_ _6506_/Q _6763_/Q _3177_/Y _5551_/B1 _5550_/Y VGND VPWR _7087_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_157_572 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4502_ _4896_/B _4462_/B _4496_/B _4900_/A _4465_/B VGND VPWR _4502_/X VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_184_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5482_ _5482_/A0 hold666/X hold50/X VGND VPWR _5482_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_609 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4433_ _4607_/A _4881_/A VGND VPWR _4691_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_104_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7152_ _7155_/CLK _7152_/D fanout449/X VGND VPWR _7152_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_116_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4364_ _4556_/A _4441_/A VGND VPWR _4690_/B VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_113_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6103_ _6507_/Q _7122_/Q _6103_/B1 VGND VPWR _6103_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_112_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3315_ hold83/X hold64/X VGND VPWR hold84/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_59_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7083_ _7083_/CLK _7083_/D fanout485/X VGND VPWR _7083_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4295_ hold958/X _6355_/A1 _4297_/S VGND VPWR _4295_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6034_ _7012_/Q _5940_/X _5967_/X _6852_/Q _6030_/X VGND VPWR _6034_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3246_ _7167_/Q _3253_/S VGND VPWR _3250_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_67_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3177_ _6509_/Q VGND VPWR _3177_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_132_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_445 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7069_/CLK _6936_/D fanout482/X VGND VPWR _6936_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XPHY_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6867_ _7067_/CLK _6867_/D fanout477/X VGND VPWR _6867_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5818_ _6825_/Q _5818_/A2 _5812_/X _5815_/X _5817_/X VGND VPWR _5818_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_4
X_6798_ _7049_/CLK _6798_/D fanout457/X VGND VPWR _6798_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_136_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5749_ _6846_/Q _5902_/A2 _5905_/A2 _6798_/Q _5739_/X VGND VPWR _5749_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_69 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold560 _6843_/Q VGND VPWR hold560/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 _5438_/X VGND VPWR _6987_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold582 _6474_/Q VGND VPWR hold582/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold593 _5399_/X VGND VPWR _6953_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1260 _4087_/X VGND VPWR _6510_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _6685_/Q VGND VPWR _4293_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _4251_/X VGND VPWR _6650_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1293 _6715_/Q VGND VPWR _4329_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_122 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_712 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_737 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_439 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4080_ hold405/X _4079_/X _4084_/S VGND VPWR _4080_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4982_ _4902_/B _4673_/A _4969_/Y _4689_/B VGND VPWR _4982_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_6721_ _3937_/A1 _6721_/D fanout487/X VGND VPWR _6721_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_51_459 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3933_ _6498_/Q input3/X input1/X VGND VPWR _3933_/X VGND VPWR sky130_fd_sc_hd__mux2_4
X_6652_ _6654_/CLK _6652_/D fanout454/X VGND VPWR _6652_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3864_ _3866_/A1 _3863_/Y _3862_/X VGND VPWR _6408_/D VGND VPWR sky130_fd_sc_hd__a21o_1
X_5603_ _6508_/Q _5601_/X _5602_/Y _7102_/Q VGND VPWR _7102_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_6583_ _7137_/CLK _6583_/D VGND VPWR _6583_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_3795_ _6460_/Q _4020_/A _4008_/A _6450_/Q VGND VPWR _3795_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_191_125 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_745 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_211 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5534_ hold261/X _5534_/A1 _5540_/S VGND VPWR _5534_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5465_ hold275/X _5465_/A1 _5471_/S VGND VPWR _5465_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4416_ _4551_/A _4549_/B VGND VPWR _4456_/A VGND VPWR sky130_fd_sc_hd__and2_2
X_5396_ hold445/X _5528_/A1 _5399_/S VGND VPWR _5396_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7135_ _7140_/CLK _7135_/D VGND VPWR _7135_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_113_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4347_ _4702_/B _4564_/A _4347_/C VGND VPWR _4376_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_99_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7066_ _7069_/CLK _7066_/D fanout477/X VGND VPWR _7066_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4278_ hold481/X _5518_/A1 _4279_/S VGND VPWR _4278_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6017_ _6819_/Q _5953_/X _5960_/X _7072_/Q _6016_/X VGND VPWR _6017_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3229_ _4563_/A VGND VPWR _4441_/A VGND VPWR sky130_fd_sc_hd__inv_6
XFILLER_39_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VPWR _3942_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_70_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6919_ _6999_/CLK _6919_/D fanout465/X VGND VPWR _6919_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_23_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_334 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_689 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_520 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_692 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold390 _4254_/X VGND VPWR _6653_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_770 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_483 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1090 _5233_/X VGND VPWR _6805_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_409 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3580_ _3580_/A _3580_/B _3580_/C _3580_/D VGND VPWR _3581_/D VGND VPWR sky130_fd_sc_hd__nor4_2
XFILLER_127_542 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5250_ _5250_/A0 _5484_/A1 _5255_/S VGND VPWR _5250_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4201_ hold942/X _5546_/A1 _4201_/S VGND VPWR _4201_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_301 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5181_ hold255/X _5465_/A1 _5181_/S VGND VPWR _5181_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4132_ hold608/X _6357_/A1 _4132_/S VGND VPWR _4132_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_68_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4063_ hold792/X _4062_/X _4067_/S VGND VPWR _4063_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4965_ _4984_/A _4965_/B _5051_/A VGND VPWR _5069_/B VGND VPWR sky130_fd_sc_hd__nand3_1
X_6704_ _6704_/CLK _6704_/D fanout450/X VGND VPWR _6704_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3916_ _6486_/Q _6489_/Q VGND VPWR _3916_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_189_291 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_442 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4896_ _4896_/A _4896_/B VGND VPWR _4911_/C VGND VPWR sky130_fd_sc_hd__and2_1
X_6635_ _7150_/CLK _6635_/D fanout487/X VGND VPWR _6635_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3847_ _6412_/Q hold70/A _3854_/S hold32/A VGND VPWR _3847_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_164_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6566_ _6755_/CLK _6566_/D fanout445/X VGND VPWR _6566_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3778_ _6906_/Q _5346_/A _4310_/A _6700_/Q VGND VPWR _3778_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_152_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5517_ hold409/X _5544_/A1 hold87/A VGND VPWR _5517_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_133_512 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6497_ _6990_/CLK _6497_/D fanout479/X VGND VPWR _7188_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5448_ hold385/X _5526_/A1 _5453_/S VGND VPWR _5448_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_154_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5379_ hold694/X _5469_/A1 _5381_/S VGND VPWR _5379_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7118_ _7130_/CLK _7118_/D fanout447/X VGND VPWR _7118_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_86_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_529 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7049_ _7049_/CLK _7049_/D fanout456/X VGND VPWR _7049_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_170_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_206 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_78 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_102 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_597 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_383 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_353 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_396 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_70 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_743 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4750_ _4542_/D _4672_/B _4626_/Y _4628_/Y VGND VPWR _4769_/A VGND VPWR sky130_fd_sc_hd__o22a_1
X_3701_ _3700_/Y _3764_/A1 _3829_/A VGND VPWR _3701_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4681_ _5010_/B _4686_/B VGND VPWR _4681_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_186_283 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6420_ _6749_/CLK _6420_/D fanout457/X VGND VPWR _6420_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
X_3632_ _6941_/Q _5382_/A _3358_/Y input14/X _3631_/X VGND VPWR _3638_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6351_ _6641_/Q _6351_/A2 _5006_/A _6350_/X VGND VPWR _6351_/X VGND VPWR sky130_fd_sc_hd__o31a_1
X_3563_ _6966_/Q _5409_/A _4139_/A _6554_/Q VGND VPWR _3563_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_5302_ _5302_/A0 _5473_/A1 _5309_/S VGND VPWR _5302_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6282_ _7155_/Q _5958_/X _5978_/X _6484_/Q VGND VPWR _6282_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_103_707 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3494_ _6613_/Q _4208_/A _4157_/A _6569_/Q VGND VPWR _3494_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_5233_ _5233_/A0 _5545_/A1 _5237_/S VGND VPWR _5233_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_526 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_opt_3_0_csclk _6888_/CLK VGND VPWR clkbuf_opt_3_0_csclk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5164_ _5171_/B _5164_/B hold17/X VGND VPWR _5164_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_4115_ _4115_/A0 hold42/X hold38/X VGND VPWR hold55/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_5095_ _5122_/C _5126_/B _5142_/B VGND VPWR _5096_/C VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_84_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4046_ hold848/X _6354_/A1 _4049_/S VGND VPWR _4046_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_17_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_554 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5997_ _7002_/Q _5958_/X _5975_/D _6882_/Q VGND VPWR _5997_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XPHY_229 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4948_ _4948_/A _4948_/B _4948_/C _4948_/D VGND VPWR _4948_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_4879_ _4902_/B _4613_/Y _4877_/X _4878_/X _4529_/Y VGND VPWR _4880_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_138_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6618_ _6655_/CLK _6618_/D fanout469/X VGND VPWR _6618_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6549_ _6674_/CLK _6549_/D _6383_/A VGND VPWR _6549_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_161_640 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_545 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_386 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_526 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _6744_/Q VGND VPWR pll_sel[2] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput281 _6421_/Q VGND VPWR pll_trim[19] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput292 _6439_/Q VGND VPWR pll_trim[5] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_58_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_757 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_294 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_242 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xwire353 _3604_/Y VGND VPWR _3640_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_139_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire364 _6225_/Y VGND VPWR _6226_/D VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_109_361 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_320 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_397 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_462 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_348 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5920_ _6559_/Q _5667_/X _5915_/X _5916_/X _5919_/X VGND VPWR _5920_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_515 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5851_ _6696_/Q _5637_/X _5848_/X _5850_/X VGND VPWR _5852_/C VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_21_204 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4802_ _4689_/A _4631_/Y _4645_/Y _4846_/B VGND VPWR _4803_/C VGND VPWR sky130_fd_sc_hd__o22a_1
X_5782_ _6992_/Q _5627_/X _5637_/X _6952_/Q _5781_/X VGND VPWR _5787_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4733_ _4739_/B _4733_/B VGND VPWR _4747_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_174_220 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4664_ _4664_/A _4664_/B VGND VPWR _4928_/A VGND VPWR sky130_fd_sc_hd__nor2_1
X_6403_ _3927_/A1 _6403_/D _6359_/X VGND VPWR _6403_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_135_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3615_ _7042_/Q hold76/A _5182_/S _6758_/Q _3614_/X VGND VPWR _3620_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold901 _4116_/X VGND VPWR _6530_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _4595_/A _4595_/B VGND VPWR _4735_/A VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold912 _6853_/Q VGND VPWR hold912/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _5281_/X VGND VPWR _6848_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold934 _6482_/Q VGND VPWR hold934/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6333_/X _6334_/A1 _6346_/S VGND VPWR _7144_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold945 _4144_/X VGND VPWR _6554_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3546_ _3546_/A hold75/X VGND VPWR _4322_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_89_705 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold956 _6697_/Q VGND VPWR hold956/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _5304_/X VGND VPWR _6868_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _6454_/Q VGND VPWR hold978/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _3970_/X VGND VPWR _6420_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6648_/Q _5976_/C _5971_/D _6568_/Q VGND VPWR _6265_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3477_ _6999_/Q _5445_/A _5211_/A _6791_/Q _3459_/X VGND VPWR _3484_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5216_ hold118/X hold60/X hold18/X VGND VPWR _5216_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6196_ _6455_/Q _5944_/X _5975_/A _6599_/Q _6195_/X VGND VPWR _6200_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1601 _7132_/Q VGND VPWR _6306_/B2 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_315 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_484 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5147_ hold884/X _6354_/A1 _5147_/S VGND VPWR _5147_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5078_ _6724_/Q _4229_/X _5103_/B _5077_/Y _5067_/Y VGND VPWR _5078_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4029_ hold870/X _5493_/A1 hold68/X VGND VPWR _4029_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_71_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_743 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_456 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_447 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_342 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_631 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_524 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_170 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_693 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_389 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_292 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_404 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold208 _5458_/X VGND VPWR _7005_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _6997_/Q VGND VPWR hold219/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _7070_/Q _5523_/A _5319_/A _6889_/Q VGND VPWR _3400_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4380_ _4739_/A _4492_/D VGND VPWR _4896_/B VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_125_684 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3331_ _3379_/A hold36/X VGND VPWR _3331_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6050_ _6043_/X _6045_/X _6050_/C _6301_/C VGND VPWR _6050_/X VGND VPWR sky130_fd_sc_hd__and4bb_1
XFILLER_112_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3262_ _6416_/Q _3837_/A _3262_/C VGND VPWR _3262_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
XFILLER_85_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5001_ _5001_/A _5001_/B _5076_/B VGND VPWR _5004_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_3193_ _7029_/Q VGND VPWR _3193_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6952_ _6969_/CLK _6952_/D fanout475/X VGND VPWR _6952_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5903_ _6617_/Q _5628_/X _5661_/X _6622_/Q _5902_/X VGND VPWR _5906_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6883_ _7067_/CLK _6883_/D fanout477/X VGND VPWR _6883_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_5834_ _7151_/Q _5625_/X _5661_/X _6619_/Q VGND VPWR _5834_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_61_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5765_ _6967_/Q _5642_/X _5666_/X _6895_/Q VGND VPWR _5765_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4716_ _4716_/A _4965_/B _4969_/B VGND VPWR _4716_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
X_5696_ _6940_/Q _5632_/X _5638_/X _6956_/Q _5694_/X VGND VPWR _5711_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_724 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4647_ _4846_/B _4673_/A _4611_/Y _4628_/Y VGND VPWR _4647_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_107_128 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold720 _6517_/Q VGND VPWR hold720/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 _4206_/X VGND VPWR _6607_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ _4947_/B _4902_/A _4846_/B _4672_/A VGND VPWR _4578_/X VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold742 _6537_/Q VGND VPWR hold742/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 _4106_/X VGND VPWR _6521_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ _6317_/A VGND VPWR _6317_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xhold764 _6815_/Q VGND VPWR hold764/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ _3562_/A _3573_/B VGND VPWR _4151_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold775 _4048_/X VGND VPWR _6483_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _6951_/Q VGND VPWR hold786/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _4040_/X VGND VPWR _6476_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6248_ _6557_/Q _5971_/B _5949_/X _6677_/Q VGND VPWR _6248_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_39_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6179_ _6179_/A0 _6178_/X _6304_/S VGND VPWR _7126_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_69_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1420 _6596_/Q VGND VPWR hold1420/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1431 _6587_/Q VGND VPWR _4183_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1442 _6432_/Q VGND VPWR hold151/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _6947_/Q VGND VPWR _5393_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _6727_/Q VGND VPWR _3830_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _6590_/Q VGND VPWR _4186_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1486 _6254_/X VGND VPWR _7129_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_115 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1497 _6583_/Q VGND VPWR _4179_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_384 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_518 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_579 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_359 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_264 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_286 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_662 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_527 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_443 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_70 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold80 hold80/A VGND VPWR hold80/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A VGND VPWR hold91/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_643 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3880_ _6643_/Q _3962_/B _3880_/B1 VGND VPWR _6643_/D VGND VPWR sky130_fd_sc_hd__a21o_1
X_5550_ _6506_/Q _3177_/Y _3883_/X VGND VPWR _5550_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_191_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4501_ _4782_/A _5051_/B VGND VPWR _4535_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_157_584 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5481_ hold49/X _5505_/B VGND VPWR hold50/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_172_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4432_ _4460_/A _4632_/B VGND VPWR _4969_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_132_429 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7151_ _7155_/CLK _7151_/D fanout450/X VGND VPWR _7151_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_4363_ _4556_/A _4690_/A VGND VPWR _4817_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_98_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6102_ _6089_/Y _6100_/X _6101_/Y _5552_/B VGND VPWR _6102_/X VGND VPWR sky130_fd_sc_hd__a211o_1
X_3314_ hold36/X _3546_/A VGND VPWR _4118_/B VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_113_665 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7082_ _7082_/CLK _7082_/D fanout479/X VGND VPWR _7082_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_98_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4294_ hold794/X _6354_/A1 _4297_/S VGND VPWR _4294_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6033_ _7081_/Q _5976_/B _5971_/C _7041_/Q VGND VPWR _6049_/B VGND VPWR sky130_fd_sc_hd__a22o_1
X_3245_ _3875_/B _3244_/Y _3249_/B VGND VPWR _3253_/S VGND VPWR sky130_fd_sc_hd__a21oi_1
X_3176_ _3176_/A VGND VPWR _3176_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_27_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_457 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_608 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6935_ _6997_/CLK _6935_/D fanout465/X VGND VPWR _6935_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_41_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6866_ _6908_/CLK _6866_/D fanout475/X VGND VPWR _6866_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
XFILLER_22_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_186 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5817_ _6841_/Q _5657_/X _5660_/X _6809_/Q _5816_/X VGND VPWR _5817_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6797_ _7012_/CLK _6797_/D fanout458/X VGND VPWR _6797_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_41_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5748_ _5748_/A _5748_/B _5748_/C _5748_/D VGND VPWR _5748_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_5679_ _6843_/Q _5902_/A2 _5814_/B1 _6907_/Q _5678_/X VGND VPWR _5679_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold550 _5330_/X VGND VPWR _6891_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _5276_/X VGND VPWR _6843_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold572 _6907_/Q VGND VPWR hold572/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _4037_/X VGND VPWR _6474_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _7019_/Q VGND VPWR hold594/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1250 _5524_/X VGND VPWR _7063_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 _6680_/Q VGND VPWR _4287_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _4293_/X VGND VPWR _6685_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 _6735_/Q VGND VPWR _5146_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1294 _4329_/X VGND VPWR _6715_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_543 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_362 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput170 wb_we_i VGND VPWR _6320_/B VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_36_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_619 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4981_ _4981_/A _4981_/B _4981_/C _4981_/D VGND VPWR _4983_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_17_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6720_ _3937_/A1 _6720_/D fanout487/X VGND VPWR _6720_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3932_ _3931_/X _3953_/B _6403_/Q VGND VPWR _3932_/X VGND VPWR sky130_fd_sc_hd__mux2_4
XFILLER_31_140 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6651_ _6668_/CLK _6651_/D fanout452/X VGND VPWR _6651_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3863_ hold24/A _3860_/B _3866_/S VGND VPWR _3863_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_149_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5602_ _5602_/A _5602_/B VGND VPWR _5602_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_31_195 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6582_ _6709_/CLK _6582_/D _6360_/A VGND VPWR _6582_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3794_ _3794_/A _3794_/B _3794_/C VGND VPWR _3828_/A VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_192_627 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5533_ _5533_/A0 hold667/X _5540_/S VGND VPWR _5533_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_340 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_csclk _6447_/CLK VGND VPWR _7054_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5464_ _5464_/A0 _5524_/A1 _5471_/S VGND VPWR _5464_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_502 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4415_ _4415_/A _4415_/B VGND VPWR _4549_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_132_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5395_ _5395_/A0 _5545_/A1 _5399_/S VGND VPWR _5395_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7134_ _7137_/CLK _7134_/D VGND VPWR _7134_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
X_4346_ _4564_/A _4347_/C _4702_/B VGND VPWR _4376_/A VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_59_516 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6704_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_7065_ _7065_/CLK _7065_/D fanout465/X VGND VPWR _7065_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xfanout359 _6301_/C VGND VPWR _6226_/B VGND VPWR sky130_fd_sc_hd__buf_12
X_4277_ hold612/X _5544_/A1 _4279_/S VGND VPWR _4277_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6016_ _6907_/Q _5973_/A _5948_/X _6947_/Q _6015_/X VGND VPWR _6016_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3228_ _6921_/Q VGND VPWR _3228_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_39_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_435 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6918_ _7081_/CLK _6918_/D fanout478/X VGND VPWR _6918_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6849_ _6865_/CLK _6849_/D fanout464/X VGND VPWR _6849_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_10_302 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VPWR _6990_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_184_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_259 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold380 _5442_/X VGND VPWR _6991_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_451 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold391 _6809_/Q VGND VPWR hold391/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_495 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1080 _5242_/X VGND VPWR _6813_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_541 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1091 _7074_/Q VGND VPWR _5536_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_454 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_554 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4200_ hold501/X _5518_/A1 _4201_/S VGND VPWR _4200_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5180_ hold129/X hold99/X _5181_/S VGND VPWR _5180_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4131_ hold758/X _6356_/A1 _4132_/S VGND VPWR _4131_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_421 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_432 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_357 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4062_ _4115_/A0 _5538_/A1 hold37/X VGND VPWR _4062_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_95_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_316 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4964_ _4964_/A _4964_/B _4964_/C VGND VPWR _5005_/B VGND VPWR sky130_fd_sc_hd__and3_1
X_6703_ _6704_/CLK _6703_/D fanout450/X VGND VPWR _6703_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_32_460 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3915_ _3954_/A _3962_/B _3908_/Y _6635_/Q VGND VPWR _6640_/D VGND VPWR sky130_fd_sc_hd__a22o_1
X_4895_ _5084_/D _4895_/B _5029_/B _5085_/A VGND VPWR _4918_/A VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_149_134 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6634_ _6659_/CLK _6634_/D _6383_/A VGND VPWR _6634_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3846_ _3845_/X _3846_/A1 _3866_/S VGND VPWR _6414_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_158_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6565_ _6755_/CLK _6565_/D _6360_/A VGND VPWR _6565_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3777_ _6970_/Q _5418_/A _3358_/Y input11/X _3776_/X VGND VPWR _3782_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_159 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5516_ hold600/X _5543_/A1 hold87/X VGND VPWR _5516_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6496_ _6990_/CLK _6496_/D fanout479/X VGND VPWR _7187_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_5447_ hold259/X _5465_/A1 _5453_/S VGND VPWR _5447_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_105_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5378_ hold477/X _5528_/A1 _5381_/S VGND VPWR _5378_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_160_398 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7117_ _7130_/CLK _7117_/D fanout447/X VGND VPWR _7117_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4329_ _4329_/A0 _6353_/A1 _4333_/S VGND VPWR _4329_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_86_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7048_ _7067_/CLK _7048_/D fanout485/X VGND VPWR _7048_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_15_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_218 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_498 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_114 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_395 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_563 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3700_ _3700_/A _3700_/B _3700_/C VGND VPWR _3700_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_4680_ _4773_/A _4737_/A VGND VPWR _4774_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_159_476 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_627 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3631_ _6703_/Q _4310_/A _4133_/A _6548_/Q VGND VPWR _3631_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_146_137 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6350_ _3910_/A _6350_/A2 _6317_/A _6349_/X _6320_/B VGND VPWR _6350_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_351 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3562_ _3562_/A _3562_/B VGND VPWR _4139_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_127_362 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5301_ _5301_/A _5505_/B VGND VPWR _5309_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_6281_ _6613_/Q _5943_/X _5981_/X _6659_/Q VGND VPWR _6281_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3493_ _3571_/A hold66/X VGND VPWR _4157_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5232_ hold850/X _5484_/A1 _5237_/S VGND VPWR _5232_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_170_674 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_110 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5163_ hold852/X _6354_/A1 _5163_/S VGND VPWR _5163_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_603 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4114_ hold812/X _5546_/A1 hold38/X VGND VPWR _4114_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_56_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5094_ _4948_/C _4946_/X _5058_/A _5093_/X _4818_/X VGND VPWR _5142_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_4045_ _4045_/A0 _5491_/A1 _4049_/S VGND VPWR _4045_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_714 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_566 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5996_ _7079_/Q _5976_/B _5975_/C _6834_/Q _5995_/X VGND VPWR _6000_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4947_ _4947_/A _4947_/B _4947_/C VGND VPWR _5043_/B VGND VPWR sky130_fd_sc_hd__nand3_2
X_4878_ _5083_/A _5029_/A _4878_/C VGND VPWR _4878_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_6617_ _6769_/CLK _6617_/D fanout469/X VGND VPWR _6617_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_20_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3829_ _3829_/A _3829_/B VGND VPWR _3829_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_146_660 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_276 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6548_ _6735_/CLK _6548_/D fanout445/X VGND VPWR _6548_/Q VGND VPWR sky130_fd_sc_hd__dfstp_4
XFILLER_192_287 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6479_ _6707_/CLK _6479_/D _3946_/B VGND VPWR _6479_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_161_652 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput260 _6750_/Q VGND VPWR pll_bypass VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput271 _6434_/Q VGND VPWR pll_trim[0] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_121_538 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput282 _6435_/Q VGND VPWR pll_trim[1] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_181_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput293 _6440_/Q VGND VPWR pll_trim[6] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_87_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_669 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_240 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_485 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xwire354 _3504_/Y VGND VPWR _3582_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire365 _6200_/Y VGND VPWR _6201_/B VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_99_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_373 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_86 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_544 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5850_ _6566_/Q _5635_/X _5661_/X _6620_/Q _5849_/X VGND VPWR _5850_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4801_ _4673_/B _4700_/Y _4707_/Y _4799_/X _4800_/X VGND VPWR _4804_/B VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_61_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5781_ _6848_/Q _5902_/A2 _5654_/X _6936_/Q VGND VPWR _5781_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_21_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4732_ _4428_/Y _4611_/Y _4500_/A VGND VPWR _5114_/B VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_187_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_424 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4663_ _4716_/A _4686_/B VGND VPWR _4663_/Y VGND VPWR sky130_fd_sc_hd__nand2_2
X_6402_ _3927_/A1 _6402_/D _6358_/X VGND VPWR _6402_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3614_ _6745_/Q _5154_/A _3585_/Y input95/X VGND VPWR _3614_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4594_ _4563_/A _4661_/A _4441_/B _4631_/D VGND VPWR _4595_/B VGND VPWR sky130_fd_sc_hd__a31o_1
Xhold902 _6719_/Q VGND VPWR hold902/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 _5287_/X VGND VPWR _6853_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold924 _6968_/Q VGND VPWR hold924/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _6642_/Q _6333_/A2 _6333_/B1 _6350_/A2 _6332_/X VGND VPWR _6333_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3545_ _6958_/Q _5400_/A _4127_/A _6544_/Q _3544_/X VGND VPWR _3552_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold935 _4047_/X VGND VPWR _6482_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _6564_/Q VGND VPWR hold946/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _4307_/X VGND VPWR _6697_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold968 _6477_/Q VGND VPWR hold968/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6264_ _6264_/A _6264_/B _6264_/C VGND VPWR _6276_/C VGND VPWR sky130_fd_sc_hd__nor3_1
Xhold979 _4013_/X VGND VPWR _6454_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3476_ _6879_/Q _5310_/A hold49/A _7031_/Q _3475_/X VGND VPWR _3485_/B VGND VPWR
+ sky130_fd_sc_hd__a221oi_1
X_5215_ hold225/X _5494_/A1 hold18/X VGND VPWR _5215_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_130_335 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6195_ _6465_/Q _5937_/X _5975_/D _6625_/Q VGND VPWR _6195_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold1602 _7123_/Q VGND VPWR _6128_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5146_ _5146_/A0 _5491_/A1 _5147_/S VGND VPWR _5146_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_111_571 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_327 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5077_ _5077_/A _5103_/C _5077_/C VGND VPWR _5077_/Y VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_84_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4028_ _4028_/A0 _5492_/A1 hold68/X VGND VPWR _4028_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_588 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5979_ _5979_/A _5981_/A _5979_/C VGND VPWR _5979_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_40_569 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_711 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_76 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_693 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_630 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_216 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_687 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_335 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_536 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_711 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_210 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold209 _6758_/Q VGND VPWR hold209/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_166_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3330_ _3543_/A _3373_/B VGND VPWR _5391_/A VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_125_696 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_481 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3261_ _6417_/Q _6415_/Q _6485_/Q _3164_/Y VGND VPWR _3261_/X VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_98_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5000_ _4948_/C _4582_/Y _4941_/D _4991_/X VGND VPWR _5076_/B VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_22_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3192_ _6445_/Q VGND VPWR _3192_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_636 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6951_ _6951_/CLK _6951_/D fanout474/X VGND VPWR _6951_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_19_371 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5902_ _6602_/Q _5902_/A2 _5634_/X _6453_/Q VGND VPWR _5902_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6882_ _6882_/CLK _6882_/D fanout475/X VGND VPWR _6882_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_5833_ _6560_/Q _5631_/X _5830_/X _5832_/X VGND VPWR _5833_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_14_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5764_ _7015_/Q _5630_/X _5761_/X _5762_/X _5763_/X VGND VPWR _5764_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_1
XFILLER_147_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4715_ _4469_/A _4714_/X _4713_/X _5084_/C _5062_/B VGND VPWR _4722_/C VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
XFILLER_30_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5695_ _7020_/Q _5619_/X _5663_/X _6860_/Q VGND VPWR _5695_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4646_ _4646_/A _4707_/C VGND VPWR _4646_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_190_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_544 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold710 _6959_/Q VGND VPWR hold710/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _4101_/X VGND VPWR _6517_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _4672_/A _4902_/A VGND VPWR _4723_/B VGND VPWR sky130_fd_sc_hd__nor2_1
Xhold732 _7188_/A VGND VPWR hold732/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_408 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold743 _4124_/X VGND VPWR _6537_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _6745_/Q VGND VPWR hold754/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _6320_/B _6316_/A2 _6640_/Q VGND VPWR _6317_/A VGND VPWR sky130_fd_sc_hd__a21bo_1
XFILLER_89_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold765 _5244_/X VGND VPWR _6815_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3528_ _6438_/Q _3372_/Y hold76/A _7043_/Q _3527_/X VGND VPWR _3538_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold776 _6478_/Q VGND VPWR hold776/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _5397_/X VGND VPWR _6951_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 _6886_/Q VGND VPWR hold798/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ _6457_/Q _5944_/X _5975_/A _6601_/Q _6246_/X VGND VPWR _6250_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3459_ _6799_/Q _3326_/Y _4102_/A _7200_/A VGND VPWR _3459_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_69_271 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1410 _6424_/Q VGND VPWR _3978_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6178_ _6178_/A0 _6177_/X _6303_/S VGND VPWR _6178_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold1421 _6598_/Q VGND VPWR hold1421/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 _6574_/Q VGND VPWR _4168_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1443 _3988_/X VGND VPWR _6432_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _5113_/X _5129_/B _5129_/C _5129_/D VGND VPWR _6725_/D VGND VPWR sky130_fd_sc_hd__nand4b_1
Xhold1454 _6730_/Q VGND VPWR _3642_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _6433_/Q VGND VPWR hold557/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1476 _6597_/Q VGND VPWR _4194_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1487 _6414_/Q VGND VPWR _3846_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 _6486_/Q VGND VPWR _3911_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_80_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_744 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_61 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_688 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_400 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_539 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_495 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold70 hold70/A VGND VPWR hold70/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold81 hold81/A VGND VPWR hold81/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A VGND VPWR hold92/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_380 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_580 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4500_ _4500_/A _4689_/A VGND VPWR _4500_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_184_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5480_ _5480_/A0 hold22/X hold30/X VGND VPWR hold31/A VGND VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_1 _7157_/D VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
X_4431_ _4753_/A _4460_/A VGND VPWR _4881_/A VGND VPWR sky130_fd_sc_hd__nor2_2
XFILLER_6_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_7150_ _7150_/CLK _7150_/D _6307_/B VGND VPWR _7150_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4362_ _4911_/A _4489_/A VGND VPWR _4500_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_6101_ _6790_/Q _6226_/B VGND VPWR _6101_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
X_3313_ _3313_/A _3454_/A VGND VPWR _3546_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_7081_ _7081_/CLK _7081_/D fanout485/X VGND VPWR _7081_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4293_ _4293_/A0 _5491_/A1 _4297_/S VGND VPWR _4293_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6032_ _7057_/Q _5954_/X _5976_/D _6876_/Q VGND VPWR _6049_/A VGND VPWR sky130_fd_sc_hd__a22o_1
X_3244_ _3875_/C _3260_/S VGND VPWR _3244_/Y VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_67_753 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3175_ _7089_/Q VGND VPWR _3886_/B VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_82_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_200 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_233 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_244 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_469 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6934_ _7081_/CLK _6934_/D fanout478/X VGND VPWR _6934_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6865_ _6865_/CLK _6865_/D fanout465/X VGND VPWR _6865_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_22_344 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5816_ _7025_/Q _5619_/X _5663_/X _6865_/Q VGND VPWR _5816_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6796_ _7011_/CLK _6796_/D fanout456/X VGND VPWR _6796_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_22_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5747_ _6822_/Q _5818_/A2 _5814_/B1 _6910_/Q _5746_/X VGND VPWR _5748_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_175_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5678_ _6899_/Q _5621_/X _5818_/A2 _6819_/Q VGND VPWR _5678_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4629_ _4716_/A _4975_/A _4698_/C VGND VPWR _5099_/B VGND VPWR sky130_fd_sc_hd__nand3_2
XFILLER_151_739 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold540 _4049_/X VGND VPWR _6484_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _6867_/Q VGND VPWR hold551/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold562 _6582_/Q VGND VPWR hold562/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _5348_/X VGND VPWR _6907_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _7009_/Q VGND VPWR hold584/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _5474_/X VGND VPWR _7019_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_517 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_165 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_64 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_742 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1240 _5515_/X VGND VPWR _7055_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_572 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1251 _6625_/Q VGND VPWR _4233_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1262 _4287_/X VGND VPWR _6680_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1273 _6705_/Q VGND VPWR _4317_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 _5146_/X VGND VPWR _6735_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 _6604_/Q VGND VPWR _4203_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_417 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_697 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_319 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_585 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_374 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_587 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_471 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_493 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_771 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_625 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_230 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput160 wb_dat_i[6] VGND VPWR _6342_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4980_ _4619_/Y _4970_/Y _4975_/Y _4644_/Y _5062_/A VGND VPWR _4981_/D VGND VPWR
+ sky130_fd_sc_hd__o221a_1
XFILLER_51_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3931_ _3930_/X input38/X _6405_/Q VGND VPWR _3931_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6650_ _6668_/CLK _6650_/D fanout452/X VGND VPWR _6650_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_3862_ _3167_/Y _3866_/S _3860_/B hold24/A VGND VPWR _3862_/X VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_176_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5601_ _5968_/A _5964_/A _5981_/A VGND VPWR _5601_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_6581_ _6709_/CLK _6581_/D fanout445/X VGND VPWR _6581_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3793_ _3793_/A _3793_/B _3793_/C _3793_/D VGND VPWR _3794_/C VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_118_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5532_ _5532_/A _5541_/B VGND VPWR _5540_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_191_149 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_csclk _6601_/CLK VGND VPWR _6659_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_5463_ _5463_/A hold17/X VGND VPWR _5471_/S VGND VPWR sky130_fd_sc_hd__and2_4
X_4414_ _4459_/B _4579_/A VGND VPWR _4542_/A VGND VPWR sky130_fd_sc_hd__nand2_8
X_5394_ hold363/X _5526_/A1 _5399_/S VGND VPWR _5394_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_132_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7133_ _7137_/CLK _7133_/D VGND VPWR _7133_/Q VGND VPWR sky130_fd_sc_hd__dfxtp_1
XFILLER_113_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4345_ _4631_/D _4633_/B _4661_/A _4357_/B VGND VPWR _4347_/C VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_59_528 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7064_ _7067_/CLK _7064_/D fanout477/X VGND VPWR _7064_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4276_ hold421/X _5534_/A1 _4279_/S VGND VPWR _4276_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_100_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3227_ _6792_/Q VGND VPWR _3227_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_6015_ _6899_/Q _5976_/C _5971_/D _6827_/Q VGND VPWR _6015_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_82_575 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6917_ _7085_/CLK _6917_/D fanout477/X VGND VPWR _6917_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_23_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6848_ _7069_/CLK _6848_/D fanout482/X VGND VPWR _6848_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6779_ _6969_/CLK _6779_/D fanout473/X VGND VPWR _6779_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_10_347 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_547 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold370 _5268_/X VGND VPWR _6836_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _6796_/Q VGND VPWR hold381/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _5237_/X VGND VPWR _6809_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_314 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_339 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1070 _5377_/X VGND VPWR _6933_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 _7082_/Q VGND VPWR _5545_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 _5536_/X VGND VPWR _7074_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_553 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_214 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_466 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_739 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4130_ hold952/X _6355_/A1 _4132_/S VGND VPWR _4130_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_96_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_444 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4061_ _4061_/A0 _4060_/X _4067_/S VGND VPWR _4061_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_328 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_350 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4963_ _4963_/A _4963_/B VGND VPWR _4963_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_6702_ _7155_/CLK _6702_/D fanout450/X VGND VPWR _6702_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3914_ _3837_/B _3875_/X _3875_/B _6488_/Q VGND VPWR _6487_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_1
X_4894_ _4689_/A _4631_/Y _5034_/B _4518_/C VGND VPWR _5085_/A VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_149_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_146 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6633_ _6659_/CLK _6633_/D fanout469/X VGND VPWR _6633_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3845_ _3288_/Y hold33/A _3845_/S VGND VPWR _3845_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_105 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6564_ _6674_/CLK _6564_/D _6383_/A VGND VPWR _6564_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_138_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3776_ _6994_/Q _5445_/A _3367_/Y input20/X VGND VPWR _3776_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_118_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5515_ _5515_/A0 hold667/X hold87/A VGND VPWR _5515_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6495_ _6990_/CLK _6495_/D fanout478/X VGND VPWR _7186_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_105_205 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5446_ _5446_/A0 _5524_/A1 _5453_/S VGND VPWR _5446_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_172_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5377_ _5377_/A0 _5545_/A1 _5381_/S VGND VPWR _5377_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7116_ _7130_/CLK _7116_/D fanout447/X VGND VPWR _7116_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_59_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4328_ _4328_/A _5490_/B VGND VPWR _4333_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_87_656 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7047_ _7049_/CLK _7047_/D fanout457/X VGND VPWR _7047_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4259_ hold642/X _5544_/A1 _4261_/S VGND VPWR _4259_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_266 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_126 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_138 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_95 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_100 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_199 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_288 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_709 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_409 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_411 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_422 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6747_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_147_639 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3630_ _6789_/Q _5211_/A _4044_/A _6483_/Q _3629_/X VGND VPWR _3638_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3561_ _6934_/Q _5373_/A _5154_/A _6746_/Q _3560_/X VGND VPWR _3565_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5300_ hold606/X _5513_/A1 _5300_/S VGND VPWR _5300_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6280_ _6664_/Q _5976_/B _5971_/C _6714_/Q VGND VPWR _6280_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3492_ _3562_/A _3814_/B VGND VPWR _4208_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_5231_ hold537/X _5543_/A1 _5237_/S VGND VPWR _5231_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_142_377 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_686 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5162_ _5162_/A0 _6353_/A1 _5163_/S VGND VPWR _5162_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_12_csclk _6601_/CLK VGND VPWR _6671_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4113_ hold692/X _5509_/A1 hold38/X VGND VPWR _4113_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5093_ _4672_/B _4496_/Y _4456_/Y VGND VPWR _5093_/X VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_84_615 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4044_ _4044_/A _6352_/B VGND VPWR _4049_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_83_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7081_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_52_501 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5995_ _7055_/Q _5954_/X _5976_/C _6898_/Q VGND VPWR _5995_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_52_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4946_ _4947_/A _4947_/B _4947_/C VGND VPWR _4946_/X VGND VPWR sky130_fd_sc_hd__and3_2
XFILLER_33_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4877_ _4877_/A _4877_/B _4877_/C _4877_/D VGND VPWR _4877_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_6616_ _6655_/CLK _6616_/D fanout469/X VGND VPWR _6616_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3828_ _3828_/A _3828_/B VGND VPWR _3828_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_6547_ _6654_/CLK _6547_/D fanout454/X VGND VPWR _6547_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_192_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_3759_ input72/X _3331_/Y _4238_/A _6631_/Q _3758_/X VGND VPWR _3760_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_672 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_160 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6478_ _6704_/CLK _6478_/D fanout448/X VGND VPWR _6478_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_145_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_664 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5429_ hold299/X _5465_/A1 _5435_/S VGND VPWR _5429_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput250 _3944_/Y VGND VPWR pad_flash_csb_oeb VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput261 _6736_/Q VGND VPWR pll_dco_ena VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput272 _6428_/Q VGND VPWR pll_trim[10] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput283 _6422_/Q VGND VPWR pll_trim[20] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_58_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xoutput294 _6441_/Q VGND VPWR pll_trim[7] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_181_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_506 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_628 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_200 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_497 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xwire355 _3467_/Y VGND VPWR _3486_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_99_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xwire366 _6049_/Y VGND VPWR _6050_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_266 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_65 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_1_wb_clk_i/A VGND VPWR clkbuf_2_3_0_wb_clk_i/A VGND
+ VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_151_130 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_344 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_82 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4800_ _4902_/B _4673_/A _4616_/Y VGND VPWR _4800_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_5780_ _6832_/Q _5635_/X _5928_/A2 _6840_/Q _5779_/X VGND VPWR _5787_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4731_ _4538_/X _4683_/X _4730_/X _5006_/A _4731_/B2 VGND VPWR _6720_/D VGND VPWR
+ sky130_fd_sc_hd__o32a_1
XFILLER_30_740 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4662_ _4686_/B VGND VPWR _4662_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_147_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6401_ _6401_/A _6401_/B VGND VPWR _6401_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3613_ _6965_/Q _5409_/A _3367_/Y input23/X _3612_/X VGND VPWR _3620_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4593_ _4920_/B VGND VPWR _4593_/Y VGND VPWR sky130_fd_sc_hd__inv_2
Xhold903 _4333_/X VGND VPWR _6719_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 _6845_/Q VGND VPWR hold914/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6332_ _6644_/Q _6332_/A2 _6332_/B1 _6643_/Q VGND VPWR _6332_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold925 _5416_/X VGND VPWR _6968_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ _6878_/Q _5310_/A _4328_/A _6719_/Q VGND VPWR _3544_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold936 _6606_/Q VGND VPWR hold936/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _4156_/X VGND VPWR _6564_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _6687_/Q VGND VPWR hold958/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold969 _4041_/X VGND VPWR _6477_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _6463_/Q _5945_/X _5975_/C _6581_/Q _6262_/X VGND VPWR _6264_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3475_ _6919_/Q _5355_/A _5238_/A _6815_/Q _3474_/X VGND VPWR _3475_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_142_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_325 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5214_ _5214_/A0 hold6/X hold18/X VGND VPWR _5214_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6194_ _6680_/Q _5934_/X _5975_/B _6614_/Q _6193_/X VGND VPWR _6200_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_604 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1603 _7126_/Q VGND VPWR _6203_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5145_ _5145_/A _6352_/B VGND VPWR _5147_/S VGND VPWR sky130_fd_sc_hd__and2_1
XFILLER_151_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5076_/A _5076_/B _5076_/C VGND VPWR _5077_/C VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_44_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4027_ _4027_/A0 _6353_/A1 hold68/X VGND VPWR _4027_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_16 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_342 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5978_ _5978_/A _5981_/A _5979_/C VGND VPWR _5978_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4929_ _4673_/A _4613_/Y _4772_/A _4928_/Y VGND VPWR _5002_/C VGND VPWR sky130_fd_sc_hd__o211a_1
XFILLER_166_723 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_773 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xmgmt_gpio_9_buff_inst _3927_/X VGND VPWR mgmt_gpio_out[9] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_69_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_697 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_629 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_681 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_523 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_303 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_436 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_575 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_236 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_491 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_247 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_601 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3260_ _3251_/A _3260_/A1 _3260_/S VGND VPWR _7160_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_140_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3191_ _7042_/Q VGND VPWR _3191_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_78_261 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_272 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_732 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_648 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_242 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_158 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6950_ _7067_/CLK _6950_/D fanout476/X VGND VPWR _6950_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_19_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5901_ _6607_/Q _5648_/X _5663_/X _6612_/Q _5900_/X VGND VPWR _5906_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_6881_ _7070_/CLK _6881_/D fanout473/X VGND VPWR _6881_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_5832_ _6645_/Q _5621_/X _5648_/X _6604_/Q _5831_/X VGND VPWR _5832_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5763_ _6951_/Q _5637_/X _5645_/X _7031_/Q VGND VPWR _5763_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4714_ _4633_/B _4627_/A _4479_/Y _4619_/Y _4645_/Y VGND VPWR _4714_/X VGND VPWR
+ sky130_fd_sc_hd__o311a_1
X_5694_ _7004_/Q _5625_/X _5661_/X _6876_/Q VGND VPWR _5694_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_4645_ _4716_/A _4645_/B VGND VPWR _4645_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_147_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_597 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_214 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold700 _6977_/Q VGND VPWR hold700/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_556 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold711 _5406_/X VGND VPWR _6959_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4576_ _4965_/B _4576_/B VGND VPWR _4576_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold722 _6800_/Q VGND VPWR hold722/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 _4067_/X VGND VPWR _6497_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 _6449_/Q VGND VPWR hold744/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _3410_/Y _6315_/A1 _6315_/S VGND VPWR _7140_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_190_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold755 _5158_/X VGND VPWR _6745_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ _6942_/Q _5382_/A _5211_/A _6790_/Q VGND VPWR _3527_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_163 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold766 _6782_/Q VGND VPWR hold766/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 _4042_/X VGND VPWR _6478_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_548 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold788 _6887_/Q VGND VPWR hold788/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 _5324_/X VGND VPWR _6886_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6467_/Q _5937_/X _5975_/D _6627_/Q VGND VPWR _6246_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3458_ input17/X _3358_/Y _3372_/Y _6439_/Q VGND VPWR _3458_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_76_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6177_ _6793_/Q _6226_/B _6176_/X VGND VPWR _6177_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
Xhold1400 _7031_/Q VGND VPWR _5487_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3389_ _6929_/Q _5364_/A _3365_/Y input10/X _3386_/X VGND VPWR _3392_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1411 _7173_/A VGND VPWR _5173_/B1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 _6585_/Q VGND VPWR hold1422/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1433 _7140_/Q VGND VPWR _6315_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5128_ _5142_/A _5126_/X _5142_/C _5123_/Y VGND VPWR _5129_/C VGND VPWR sky130_fd_sc_hd__a31o_1
XFILLER_57_445 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1444 _6624_/Q VGND VPWR _3963_/S VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _3642_/X VGND VPWR _6730_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1466 _3989_/X VGND VPWR _6433_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_478 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1477 _6734_/Q VGND VPWR _3413_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1488 _6636_/Q VGND VPWR _6641_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5059_ _5058_/X _5122_/A VGND VPWR _5059_/X VGND VPWR sky130_fd_sc_hd__and2b_1
XFILLER_55_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1499 _3911_/X VGND VPWR _6486_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_684 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_172 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_548 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_391 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_222 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_756 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_412 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold60 hold60/A VGND VPWR hold60/X VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_29_93 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold71 hold71/A VGND VPWR hold71/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_467 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold82 hold82/A VGND VPWR hold82/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_489 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold93 hold93/A VGND VPWR hold93/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_139 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_312 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_155 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_166 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_345 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_177 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_356 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4430_ _5068_/A VGND VPWR _4430_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XANTENNA_2 _5190_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_567 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_461 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_589 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4361_ _4911_/A _4489_/A VGND VPWR _4685_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_6100_ _6092_/X _6094_/X _6100_/C _6301_/C VGND VPWR _6100_/X VGND VPWR sky130_fd_sc_hd__and4bb_2
X_3312_ hold26/X hold46/X VGND VPWR _3454_/A VGND VPWR sky130_fd_sc_hd__and2b_4
XFILLER_140_431 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7080_ _7080_/CLK _7080_/D fanout479/X VGND VPWR _7080_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_4292_ _4292_/A _5490_/B VGND VPWR _4297_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_58_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6031_ _7004_/Q _5958_/X _5978_/X _6996_/Q VGND VPWR _6031_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3243_ _6487_/Q _3837_/C VGND VPWR _3260_/S VGND VPWR sky130_fd_sc_hd__nand2_8
XFILLER_100_317 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_328 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3174_ _6763_/Q VGND VPWR _3174_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6933_ _7082_/CLK _6933_/D fanout483/X VGND VPWR _6933_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6864_ _6951_/CLK _6864_/D fanout474/X VGND VPWR _6864_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
X_5815_ _6817_/Q _5667_/X _5813_/X _5814_/X VGND VPWR _5815_/X VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_22_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6795_ _6963_/CLK _6795_/D fanout456/X VGND VPWR _6795_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_5746_ _6998_/Q _5643_/X _5652_/B _6918_/Q _5651_/Y VGND VPWR _5746_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_41_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_553 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5677_ _6795_/Q _5905_/A2 _5660_/X _6803_/Q VGND VPWR _5677_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_135_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4628_ _4661_/A _4716_/A _4653_/B VGND VPWR _4628_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
XFILLER_190_331 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold530 _4207_/X VGND VPWR _6608_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _6875_/Q VGND VPWR hold541/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _5088_/B _4559_/B _4721_/A VGND VPWR _4559_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_89_312 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold552 _5303_/X VGND VPWR _6867_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold563 _4177_/X VGND VPWR _6582_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_634 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold574 _6439_/Q VGND VPWR hold574/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold585 _5462_/X VGND VPWR _7009_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold596 _6562_/Q VGND VPWR hold596/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_144 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6229_ _6229_/A0 _6228_/X _6279_/S VGND VPWR _7128_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_66_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold1230 _5497_/X VGND VPWR _7039_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_551 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1241 _6710_/Q VGND VPWR _4323_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _4233_/X VGND VPWR _6625_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_584 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1263 _6480_/Q VGND VPWR _4045_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _4317_/X VGND VPWR _6705_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 _6609_/Q VGND VPWR _4209_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 _4203_/X VGND VPWR _6604_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_103 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_637 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_186 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_331 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_83 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_72 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_280 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_dat_i[26] VGND VPWR _6330_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VPWR _6345_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_651 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3930_ _6499_/Q _6734_/Q _6400_/B VGND VPWR _3930_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_44_470 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_183 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3861_ _3861_/A _3861_/B VGND VPWR _6409_/D VGND VPWR sky130_fd_sc_hd__xnor2_1
XFILLER_189_486 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5600_ _5600_/A _7102_/Q VGND VPWR _5981_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_6580_ _6677_/CLK _6580_/D fanout452/X VGND VPWR _6580_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3792_ _6442_/Q _3999_/A _5182_/S _7087_/Q _3791_/X VGND VPWR _3793_/D VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_607 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5531_ hold176/X hold22/X _5531_/S VGND VPWR _5531_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_145_501 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_203 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5462_ hold584/X _5513_/A1 _5462_/S VGND VPWR _5462_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_4413_ _4549_/A _4579_/A VGND VPWR _4413_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
X_5393_ _5393_/A0 hold13/X _5399_/S VGND VPWR hold10/A VGND VPWR sky130_fd_sc_hd__mux2_1
X_7132_ _7150_/CLK _7132_/D fanout487/X VGND VPWR _7132_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_141_740 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4344_ _4631_/D _4661_/A _4357_/B VGND VPWR _4352_/B VGND VPWR sky130_fd_sc_hd__nand3_1
XFILLER_125_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_304 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_164 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7063_ _7063_/CLK _7063_/D fanout463/X VGND VPWR _7063_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_101_626 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4275_ _4275_/A0 hold667/X _4279_/S VGND VPWR _4275_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6014_ _6014_/A _6014_/B _6014_/C VGND VPWR _6014_/Y VGND VPWR sky130_fd_sc_hd__nor3_1
X_3226_ _6919_/Q VGND VPWR _3226_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_100_136 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6916_ _7081_/CLK _6916_/D fanout478/X VGND VPWR _6916_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_70_749 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_654 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_626 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6847_ _6951_/CLK _6847_/D fanout474/X VGND VPWR _6847_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_167_147 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6778_ _6969_/CLK _6778_/D fanout473/X VGND VPWR _6778_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_106 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_670 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5729_ _7021_/Q _5619_/X _5663_/X _6861_/Q VGND VPWR _5729_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_108_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
Xhold360 _5178_/X VGND VPWR _6759_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _7065_/Q VGND VPWR hold371/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _5223_/X VGND VPWR _6796_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _7180_/A VGND VPWR hold393/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1060 _5341_/X VGND VPWR _6901_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _6821_/Q VGND VPWR _5251_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1082 _5545_/X VGND VPWR _7082_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 _6748_/Q VGND VPWR _5162_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _4102_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_60_226 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_401 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_440 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_142 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_473 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_629 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_386 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_570 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_635 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4060_ hold812/X _5546_/A1 hold37/X VGND VPWR _4060_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_110_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_307 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_573 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_489 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_392 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_362 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_470 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4962_ _4950_/X _4962_/B _4962_/C VGND VPWR _4963_/B VGND VPWR sky130_fd_sc_hd__and3b_1
XFILLER_51_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6701_ _7155_/CLK _6701_/D fanout449/X VGND VPWR _6701_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3913_ _3164_/Y _3165_/Y _3868_/S _3867_/B _6488_/Q VGND VPWR _6488_/D VGND VPWR
+ sky130_fd_sc_hd__a32o_1
X_4893_ _4893_/A VGND VPWR _5034_/B VGND VPWR sky130_fd_sc_hd__inv_2
X_6632_ _6632_/CLK _6632_/D fanout454/X VGND VPWR _6632_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3844_ hold32/A _6412_/Q hold70/A _3854_/S VGND VPWR _3845_/S VGND VPWR sky130_fd_sc_hd__nand4_1
XFILLER_149_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6563_ _6674_/CLK _6563_/D _6383_/A VGND VPWR _6563_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_192_426 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3775_ _6922_/Q _5364_/A _5274_/A _6842_/Q _3774_/X VGND VPWR _3782_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5514_ hold86/X _5541_/B VGND VPWR hold87/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_118_545 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6494_ _7079_/CLK _6494_/D fanout478/X VGND VPWR _7185_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_589 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5445_ _5445_/A hold17/X VGND VPWR _5453_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_105_217 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_695 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5376_ hold864/X _5484_/A1 _5381_/S VGND VPWR _5376_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_120_209 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_613 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7115_ _7130_/CLK _7115_/D fanout447/X VGND VPWR _7115_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4327_ hold826/X _5546_/A1 _4327_/S VGND VPWR _4327_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7046_ _7086_/CLK _7046_/D fanout483/X VGND VPWR _7046_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_4258_ hold427/X _5534_/A1 _4261_/S VGND VPWR _4258_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_28_713 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_178 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3209_ _6901_/Q VGND VPWR _3209_/Y VGND VPWR sky130_fd_sc_hd__inv_2
X_4189_ _3762_/Y _4189_/A1 _4195_/S VGND VPWR _6592_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_245 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_256 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_513 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_738 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_456 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_628 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_459 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_85 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold190 _6830_/Q VGND VPWR hold190/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_581 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_721 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_668 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_csclk _6601_/CLK VGND VPWR _6769_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_61_535 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_94 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_473 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_81 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3560_ _6674_/Q _4274_/A _4133_/A _6549_/Q VGND VPWR _3560_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_155_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_515 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_683 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3491_ input56/X _5193_/A _5274_/A _6846_/Q _3490_/X VGND VPWR _3504_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5230_ _5230_/A0 _5473_/A1 _5237_/S VGND VPWR _5230_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5161_ _5161_/A _5190_/B hold16/X VGND VPWR _5163_/S VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_96_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4112_ _4112_/A0 hold6/X hold38/A VGND VPWR _4112_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5092_ _5092_/A _5092_/B _5092_/C VGND VPWR _5126_/B VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_110_275 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_498 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4043_ hold533/X _6357_/A1 _4043_/S VGND VPWR _4043_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_513 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5994_ _7063_/Q _5934_/X _5973_/A _6906_/Q _5993_/X VGND VPWR _6000_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4945_ _4930_/X _4944_/X _5069_/A VGND VPWR _4945_/Y VGND VPWR sky130_fd_sc_hd__a21boi_1
X_4876_ _4623_/Y _4700_/Y _4864_/X _4875_/X _4523_/Y VGND VPWR _4877_/D VGND VPWR
+ sky130_fd_sc_hd__o2111a_1
X_6615_ _7036_/CLK _6615_/D fanout455/X VGND VPWR _6615_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3827_ _3798_/X _3827_/B _3827_/C _3827_/D VGND VPWR _3828_/B VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_192_223 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6546_ _6677_/CLK _6546_/D fanout452/X VGND VPWR _6546_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_3758_ _6891_/Q _5328_/A _5541_/A _7080_/Q VGND VPWR _3758_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_180_407 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_150 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6477_ _6707_/CLK _6477_/D fanout450/X VGND VPWR _6477_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
X_3689_ _6948_/Q _5391_/A _5400_/A _6956_/Q VGND VPWR _3689_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_106_559 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5428_ _5428_/A0 _5524_/A1 _5435_/S VGND VPWR _5428_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput240 _3919_/X VGND VPWR mgmt_gpio_out[36] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput251 _3951_/X VGND VPWR pad_flash_io0_do VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput262 _6737_/Q VGND VPWR pll_div[0] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput273 _6429_/Q VGND VPWR pll_trim[11] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput284 _6423_/Q VGND VPWR pll_trim[21] VGND VPWR sky130_fd_sc_hd__buf_12
X_5359_ _5359_/A0 _5545_/A1 _5363_/S VGND VPWR _5359_/X VGND VPWR sky130_fd_sc_hd__mux2_1
Xoutput295 _6426_/Q VGND VPWR pll_trim[8] VGND VPWR sky130_fd_sc_hd__buf_12
XFILLER_160_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_605 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_7029_ _7082_/CLK _7029_/D fanout483/X VGND VPWR _7029_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_59_189 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_351 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_58 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_598 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_343 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_579 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_231 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_754 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_253 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_79 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_404 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_713 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_403 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_640 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire356 _3446_/Y VGND VPWR _3447_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_139_73 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xwire367 _5748_/Y VGND VPWR wire367/X VGND VPWR sky130_fd_sc_hd__clkbuf_2
XFILLER_137_673 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_356 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_142 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_389 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_608 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_576 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_181 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_568 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_20 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4730_ _5039_/A _4589_/Y _4729_/X VGND VPWR _4730_/X VGND VPWR sky130_fd_sc_hd__a21o_1
X_4661_ _4661_/A _4661_/B VGND VPWR _4686_/B VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_187_595 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_746 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6400_ _6400_/A _6400_/B VGND VPWR _6400_/X VGND VPWR sky130_fd_sc_hd__and2_1
X_3612_ _6445_/Q _3999_/A _4322_/A _6713_/Q VGND VPWR _3612_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_4592_ _4565_/X _4601_/A _6643_/Q VGND VPWR _4920_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_174_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold904 _6781_/Q VGND VPWR hold904/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6331_ _6330_/X _6331_/A1 _6346_/S VGND VPWR _7143_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3543_ _3543_/A _3577_/B VGND VPWR _4328_/A VGND VPWR sky130_fd_sc_hd__nor2_4
Xhold915 _5278_/X VGND VPWR _6845_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _7085_/Q VGND VPWR hold926/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _4205_/X VGND VPWR _6606_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 _6472_/Q VGND VPWR hold948/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 _4295_/X VGND VPWR _6687_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6668_/Q _5938_/X _5952_/X _6708_/Q VGND VPWR _6262_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3474_ _6927_/Q _5364_/A _3999_/A _6447_/Q _3473_/X VGND VPWR _3474_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_2
XFILLER_143_698 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5213_ hold251/X _5465_/A1 hold18/X VGND VPWR _5213_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6193_ _6700_/Q _5971_/A _5979_/X _6470_/Q VGND VPWR _6193_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_142_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_741 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5144_ _5123_/A _5142_/Y _5143_/Y _5136_/X VGND VPWR _6726_/D VGND VPWR sky130_fd_sc_hd__a211o_1
XFILLER_28_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5075_ _4428_/Y _4456_/Y _4846_/B _4689_/B _4768_/A VGND VPWR _5076_/C VGND VPWR
+ sky130_fd_sc_hd__o221a_1
X_4026_ hold67/X _5490_/B VGND VPWR hold68/A VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_71_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5977_ _5977_/A _5977_/B _5977_/C VGND VPWR _6301_/C VGND VPWR sky130_fd_sc_hd__nand3_4
X_4928_ _4928_/A _4984_/B VGND VPWR _4928_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_21_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_735 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_212 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4859_ _4947_/C _4689_/A _4500_/A VGND VPWR _5023_/C VGND VPWR sky130_fd_sc_hd__a21o_1
XFILLER_176_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_109 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_673 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_161 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6529_ _6990_/CLK hold55/X fanout478/X VGND VPWR _6529_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_161_484 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_623 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VPWR _7155_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_56_693 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_359 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_csclk _6601_/CLK VGND VPWR _6674_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_184_521 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_723 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_278 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_26_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7051_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_140_613 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3190_ _7050_/Q VGND VPWR _3190_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_38_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_284 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_221 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_254 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_90 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5900_ _6468_/Q _5619_/X _5652_/B _5899_/Y VGND VPWR _5900_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_81_449 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6880_ _7069_/CLK _6880_/D fanout482/X VGND VPWR _6880_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_179_315 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5831_ _6614_/Q _5628_/X _5910_/B1 _6625_/Q VGND VPWR _5831_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_34_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_348 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5762_ _6943_/Q _5632_/X _5638_/X _6959_/Q _5759_/X VGND VPWR _5762_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4713_ _5041_/B _4576_/Y _4712_/X _4711_/X VGND VPWR _4713_/X VGND VPWR sky130_fd_sc_hd__a31o_1
X_5693_ _5713_/A0 _5692_/X _6279_/S VGND VPWR _5693_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_175_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_768 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4644_ _4716_/A _4644_/B VGND VPWR _4644_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_162_226 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold701 _5426_/X VGND VPWR _6977_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4574_/A _4574_/B _4551_/A VGND VPWR _4575_/Y VGND VPWR sky130_fd_sc_hd__a21oi_1
Xhold712 _6943_/Q VGND VPWR hold712/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 _5227_/X VGND VPWR _6800_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _6581_/Q VGND VPWR hold734/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _3447_/Y _6314_/A1 _6315_/S VGND VPWR _7139_/D VGND VPWR sky130_fd_sc_hd__mux2_1
X_3526_ _6798_/Q _3326_/Y _3981_/A _6430_/Q _3525_/X VGND VPWR _3538_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_505 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold745 _4007_/X VGND VPWR _6449_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 _6458_/Q VGND VPWR hold756/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _5207_/X VGND VPWR _6782_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _6473_/Q VGND VPWR hold778/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6245_ _6682_/Q _5934_/X _5975_/B _6616_/Q _6244_/X VGND VPWR _6250_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold789 _5325_/X VGND VPWR _6887_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3457_ input8/X _3365_/Y _3367_/Y input25/X VGND VPWR _3457_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_103_337 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6176_ _6168_/X _6226_/B _6176_/C _6176_/D VGND VPWR _6176_/X VGND VPWR sky130_fd_sc_hd__and4b_2
X_3388_ input60/X _5193_/A _3326_/Y _6801_/Q _3385_/X VGND VPWR _3392_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold1401 _6881_/Q VGND VPWR _5318_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 _6576_/Q VGND VPWR hold1412/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _4948_/B _5042_/Y _5043_/Y _4948_/D VGND VPWR _5142_/C VGND VPWR sky130_fd_sc_hd__o22a_1
Xhold1423 _6590_/Q VGND VPWR hold1423/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _7135_/Q VGND VPWR _6310_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1445 _3965_/X VGND VPWR hold665/A VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 _6728_/Q VGND VPWR _3764_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1467 _6440_/Q VGND VPWR _3997_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5058_/A _5122_/B _5058_/C _5058_/D VGND VPWR _5058_/X VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_55_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1478 _6596_/Q VGND VPWR _4193_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1489 _7122_/Q VGND VPWR _6078_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4009_ _4009_/A0 _6353_/A1 _4013_/S VGND VPWR _4009_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_332 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_641 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_354 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_702 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_379 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_234 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_657 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_690 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold50 hold50/A VGND VPWR hold50/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_152_51 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold61 hold61/A VGND VPWR hold61/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_243 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold72 hold72/A VGND VPWR hold72/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VPWR hold83/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A VGND VPWR hold94/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_63_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_630 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_123 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_324 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_360 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_368 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_371 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_429 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _5346_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4360_ _4359_/Y _4360_/B _4379_/B VGND VPWR _4489_/A VGND VPWR sky130_fd_sc_hd__and3b_2
X_3311_ hold34/X _3323_/B _3311_/C VGND VPWR hold35/A VGND VPWR sky130_fd_sc_hd__nand3_2
X_4291_ hold186/X _5519_/A1 _4291_/S VGND VPWR _4291_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_193_91 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_443 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6030_ _6860_/Q _5943_/X _5981_/X _6916_/Q VGND VPWR _6030_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_3242_ _6488_/Q _6485_/Q VGND VPWR _3837_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_79_571 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3173_ _6813_/Q VGND VPWR _3173_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_66_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_107 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_725 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6932_ _7067_/CLK _6932_/D fanout476/X VGND VPWR _6932_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_47_490 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_192 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6863_ _6865_/CLK _6863_/D fanout465/X VGND VPWR _6863_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_35_685 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_156 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5814_ _6449_/Q _5614_/X _5814_/B1 _6913_/Q VGND VPWR _5814_/X VGND VPWR sky130_fd_sc_hd__a22o_1
X_6794_ _7006_/CLK _6794_/D fanout458/X VGND VPWR _6794_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_167_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_508 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_510 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5745_ hold79/A _5614_/X _5664_/X _6926_/Q _5738_/X VGND VPWR _5748_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_565 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5676_ _6443_/Q _5614_/X _5625_/X _7003_/Q _5675_/X VGND VPWR _5681_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4627_ _4627_/A _4627_/B VGND VPWR _4703_/B VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_163_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_343 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold520 _4289_/X VGND VPWR _6682_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold531 _6689_/Q VGND VPWR hold531/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _4563_/A _4484_/Y _5088_/C VGND VPWR _4721_/A VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_150_207 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold542 _5312_/X VGND VPWR _6875_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _6746_/Q VGND VPWR hold553/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _6741_/Q VGND VPWR hold564/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold575 _3996_/X VGND VPWR _6439_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ _6484_/Q _4044_/A _4250_/A _6654_/Q _3508_/X VGND VPWR _3523_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
Xhold586 _6438_/Q VGND VPWR hold586/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4489_/A _4489_/B VGND VPWR _4490_/B VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold597 _4154_/X VGND VPWR _6562_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_134 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_668 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6228_ _7127_/Q _6227_/X _6303_/S VGND VPWR _6228_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_106_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6159_ _7009_/Q _5958_/X _5978_/X _7001_/Q VGND VPWR _6159_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold1220 _5506_/X VGND VPWR _7047_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_59 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1231 _7071_/Q VGND VPWR _5533_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 _4323_/X VGND VPWR _6710_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1253 _6778_/Q VGND VPWR _5203_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _4045_/X VGND VPWR _6480_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold1275 _6695_/Q VGND VPWR _4305_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_596 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_298 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1286 _4209_/X VGND VPWR _6609_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1297 hold1589/X VGND VPWR _4119_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_184 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_534 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_387 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_305 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput140 wb_dat_i[17] VGND VPWR _6326_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_dat_i[27] VGND VPWR _6332_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_243 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xinput162 wb_dat_i[8] VGND VPWR _6324_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3860_ hold81/A _3860_/B VGND VPWR _3861_/B VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_32_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3791_ _6750_/Q _3355_/X _5164_/B _3365_/Y input34/X VGND VPWR _3791_/X VGND VPWR
+ sky130_fd_sc_hd__a32o_1
XPHY_190 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5530_ hold938/X _5548_/A1 _5531_/S VGND VPWR _5530_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_8_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5461_ hold164/X hold99/X _5461_/S VGND VPWR _5461_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7200_ _7200_/A VGND VPWR _7200_/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4412_ _4551_/A _4959_/A VGND VPWR _4579_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_5392_ _5392_/A0 _5524_/A1 _5399_/S VGND VPWR _5392_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_7131_ _7131_/CLK _7131_/D fanout459/X VGND VPWR _7131_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4343_ _4556_/A _4563_/A _4753_/A _4607_/A VGND VPWR _4357_/B VGND VPWR sky130_fd_sc_hd__o211a_2
XFILLER_141_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_7062_ _7086_/CLK _7062_/D fanout483/X VGND VPWR _7062_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4274_ _4274_/A _4322_/B VGND VPWR _4279_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_98_176 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_638 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6013_ _6979_/Q _5945_/X _5975_/C _6835_/Q _6012_/X VGND VPWR _6014_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3225_ _6659_/Q VGND VPWR _3225_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_27_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_213 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_382 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6915_ _6981_/CLK _6915_/D fanout463/X VGND VPWR _6915_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_35_471 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6846_ _7051_/CLK _6846_/D fanout476/X VGND VPWR _6846_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_22_132 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_441 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_666 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_6777_ _6777_/CLK _6777_/D fanout483/X VGND VPWR _7196_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_22_187 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3989_ hold557/X _5513_/A1 _3989_/S VGND VPWR _3989_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_148_340 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5728_ _6973_/Q _5634_/X _5722_/X _5723_/X _5727_/X VGND VPWR _5728_/X VGND VPWR
+ sky130_fd_sc_hd__a2111o_2
XFILLER_6_309 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_682 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_310 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5659_ _6834_/Q _5928_/A2 _5910_/B1 _6882_/Q VGND VPWR _5659_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_108_248 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_557 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_663 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold350 _4078_/X VGND VPWR _6502_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold361 _6628_/Q VGND VPWR hold361/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_559 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold372 _5526_/X VGND VPWR _7065_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _6523_/Q VGND VPWR hold383/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _4095_/X VGND VPWR _6514_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_273 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1050 _5277_/X VGND VPWR _6844_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 _6938_/Q VGND VPWR _5383_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _5251_/X VGND VPWR _6821_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_97 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1083 _7029_/Q VGND VPWR _5485_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_57 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1094 _5162_/X VGND VPWR _6748_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_201 _5614_/X VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_73_588 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_655 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_413 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_485 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_496 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_752 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_582 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_80 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_585 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_511 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_92 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_747 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_728 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_374 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4961_ _4957_/Y _5046_/B _5088_/D _5039_/D VGND VPWR _4962_/C VGND VPWR sky130_fd_sc_hd__and4b_1
XFILLER_17_482 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6700_ _6704_/CLK _6700_/D fanout449/X VGND VPWR _6700_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_51_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3912_ _3912_/A1 _6485_/Q _3875_/B _3912_/B1 VGND VPWR _6489_/D VGND VPWR sky130_fd_sc_hd__a31o_1
X_4892_ _4892_/A _4892_/B VGND VPWR _4893_/A VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_149_104 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6631_ _6632_/CLK _6631_/D fanout454/X VGND VPWR _6631_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3843_ hold62/A hold81/A hold24/A hold44/A VGND VPWR _3854_/S VGND VPWR sky130_fd_sc_hd__and4_1
XFILLER_177_468 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6562_ _6674_/CLK _6562_/D _6383_/A VGND VPWR _6562_/Q VGND VPWR sky130_fd_sc_hd__dfstp_2
X_3774_ _6818_/Q _5247_/A _4298_/A _6690_/Q VGND VPWR _3774_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_192_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5513_ hold650/X _5513_/A1 _5513_/S VGND VPWR _5513_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6493_ _6527_/CLK _6493_/D fanout484/X VGND VPWR _7184_/A VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_118_557 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_505 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5444_ hold685/X _5513_/A1 _5444_/S VGND VPWR _5444_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_133_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_441 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5375_ hold295/X _5465_/A1 _5381_/S VGND VPWR _5375_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_99_463 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7114_ _7130_/CLK _7114_/D fanout448/X VGND VPWR _7114_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_59_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4326_ hold303/X _5518_/A1 _4327_/S VGND VPWR _4326_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7045_ _7085_/CLK _7045_/D fanout485/X VGND VPWR _7045_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4257_ _4257_/A0 hold667/X _4261_/S VGND VPWR _4257_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_3208_ _6909_/Q VGND VPWR _3208_/Y VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4188_ _3828_/Y _4188_/A1 _4195_/S VGND VPWR _6591_/D VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_55_522 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_393 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_603 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6829_ _6967_/CLK _6829_/D fanout474/X VGND VPWR _6829_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_11_647 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_658 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_682 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_170 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_685 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_75 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_68 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_763 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold180 _6862_/Q VGND VPWR hold180/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _5261_/X VGND VPWR _6830_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_636 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_124 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_744 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_533 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_246 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_385 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_700 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_435 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_755 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_71 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_129 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_298 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_652 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_600 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_3490_ _6902_/Q _5337_/A _4232_/A _6629_/Q VGND VPWR _3490_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_527 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_162 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_695 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5160_ hold545/X _5469_/A1 _5160_/S VGND VPWR _5160_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_722 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_4111_ hold622/X _5543_/A1 hold38/X VGND VPWR _4111_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5091_ _4584_/A _5043_/B _5090_/Y VGND VPWR _5092_/C VGND VPWR sky130_fd_sc_hd__a21oi_1
XFILLER_110_232 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4042_ hold776/X _6356_/A1 _4043_/S VGND VPWR _4042_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_661 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_525 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5993_ _6978_/Q _5945_/X _5978_/X _6994_/Q VGND VPWR _5993_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_24_249 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_290 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4944_ _4944_/A _4944_/B _4944_/C VGND VPWR _4944_/X VGND VPWR sky130_fd_sc_hd__and3_1
X_4875_ _4875_/A _5034_/A _4875_/C VGND VPWR _4875_/X VGND VPWR sky130_fd_sc_hd__and3_1
XFILLER_177_254 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6614_ _7036_/CLK _6614_/D fanout455/X VGND VPWR _6614_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_165_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3826_ _3826_/A _3826_/B _3826_/C _3826_/D VGND VPWR _3826_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_20_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_129 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_235 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_490 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6545_ _6709_/CLK _6545_/D fanout445/X VGND VPWR _6545_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_2
XFILLER_146_641 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_3757_ input21/X _3367_/Y _4038_/A _6476_/Q _3756_/X VGND VPWR _3760_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_365 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6476_ _6746_/CLK _6476_/D _3946_/B VGND VPWR _6476_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
X_3688_ _3688_/A _3688_/B _3688_/C VGND VPWR _3699_/C VGND VPWR sky130_fd_sc_hd__nor3_1
Xoutput230 _7192_/X VGND VPWR mgmt_gpio_out[27] VGND VPWR sky130_fd_sc_hd__buf_12
X_5427_ _5427_/A hold17/X VGND VPWR _5435_/S VGND VPWR sky130_fd_sc_hd__and2_4
Xoutput241 _3918_/X VGND VPWR mgmt_gpio_out[37] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput252 _3948_/A VGND VPWR pad_flash_io0_ieb VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput263 _6738_/Q VGND VPWR pll_div[1] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput274 _6430_/Q VGND VPWR pll_trim[12] VGND VPWR sky130_fd_sc_hd__buf_12
Xoutput285 _6424_/Q VGND VPWR pll_trim[22] VGND VPWR sky130_fd_sc_hd__buf_12
X_5358_ hold874/X _5484_/A1 _5363_/S VGND VPWR _5358_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_59_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xoutput296 _6427_/Q VGND VPWR pll_trim[9] VGND VPWR sky130_fd_sc_hd__buf_12
X_4309_ hold578/X _6357_/A1 _4309_/S VGND VPWR _4309_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_5289_ hold702/X _5469_/A1 _5291_/S VGND VPWR _5289_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7080_/CLK _7028_/D fanout479/X VGND VPWR _7028_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_28_511 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_706 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_363 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_694 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_766 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_725 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_416 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_415 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_438 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_437 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xwire346 _3538_/Y VGND VPWR _3581_/A VGND VPWR sky130_fd_sc_hd__clkbuf_2
Xwire357 _3408_/Y VGND VPWR wire357/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_137_652 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xwire379 _5976_/Y VGND VPWR _5977_/C VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_152_611 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_173 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_655 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_154 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_62 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_95 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_197 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_60 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_414 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_341 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_32 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_405 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4660_ _4660_/A _4660_/B _4660_/C _4660_/D VGND VPWR _4660_/X VGND VPWR sky130_fd_sc_hd__and4_1
X_3611_ _3611_/A _3611_/B _3611_/C _3611_/D VGND VPWR _3611_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
X_4591_ _4591_/A _4664_/B VGND VPWR _4601_/A VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_190_717 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_6330_ _6644_/Q _6330_/A2 _6330_/B1 _6643_/Q _6329_/X VGND VPWR _6330_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_611 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold905 _5206_/X VGND VPWR _6781_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3542_ _3546_/A _3714_/B VGND VPWR _4127_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_128_696 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold916 _6861_/Q VGND VPWR hold916/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _5548_/X VGND VPWR _7085_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _7069_/Q VGND VPWR hold938/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 _4035_/X VGND VPWR _6472_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6261_ _6453_/Q _5947_/X _5965_/X _6548_/Q _6260_/X VGND VPWR _6264_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_3473_ _7007_/Q _3370_/Y _5182_/S _3450_/X VGND VPWR _3473_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_88_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_519 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5212_ _5212_/A0 _5524_/A1 hold18/X VGND VPWR _5212_/X VGND VPWR sky130_fd_sc_hd__mux2_1
X_6192_ _6560_/Q _5953_/X _5960_/X _6670_/Q _6191_/X VGND VPWR _6192_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_5143_ _5143_/A _5143_/B VGND VPWR _5143_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
XFILLER_57_617 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5074_ _5074_/A _5074_/B _5074_/C VGND VPWR _5103_/C VGND VPWR sky130_fd_sc_hd__and3_1
X_4025_ hold213/X hold60/X _4025_/S VGND VPWR _4025_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_84_458 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_650 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_182 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5976_ _5981_/A _5976_/B _5976_/C _5976_/D VGND VPWR _5976_/Y VGND VPWR sky130_fd_sc_hd__nor4_1
XFILLER_12_208 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_219 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4927_ _4542_/B _4562_/Y _4771_/A VGND VPWR _4995_/B VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_21_764 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4482_/B _4694_/Y _4529_/Y VGND VPWR _4858_/X VGND VPWR sky130_fd_sc_hd__o21a_1
XFILLER_119_630 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3809_ _6930_/Q _5373_/A _4151_/A _6560_/Q _3808_/X VGND VPWR _3817_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_285 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4789_ _4672_/A _4620_/Y _4701_/Y _4710_/Y VGND VPWR _4789_/X VGND VPWR sky130_fd_sc_hd__o22a_1
X_6528_ _7079_/CLK _6528_/D fanout478/X VGND VPWR _6528_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_7_csclk clkbuf_3_1_0_csclk/X VGND VPWR _7038_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_6459_ _6704_/CLK _6459_/D fanout448/X VGND VPWR _6459_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_134_677 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_349 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_657 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_679 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_653 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_569 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_405 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_500 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_449 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_757 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_121 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_506 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_625 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_70 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_617 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_296 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_650 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_277 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5830_ _6480_/Q _5643_/X _5664_/X _6665_/Q VGND VPWR _5830_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_34_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5761_ _6847_/Q _5902_/A2 _5905_/A2 _6799_/Q _5760_/X VGND VPWR _5761_/X VGND VPWR
+ sky130_fd_sc_hd__a221o_1
X_4712_ _4691_/A _4673_/B _4710_/Y VGND VPWR _4712_/X VGND VPWR sky130_fd_sc_hd__o21a_1
X_5692_ _7106_/Q _5691_/X _6303_/S VGND VPWR _5692_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_175_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4643_ _4653_/C _4661_/B VGND VPWR _4643_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
X_4574_ _4574_/A _4574_/B VGND VPWR _4574_/Y VGND VPWR sky130_fd_sc_hd__nand2_1
Xhold702 _6855_/Q VGND VPWR hold702/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _5388_/X VGND VPWR _6943_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_430 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
Xhold724 _6688_/Q VGND VPWR hold724/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ _3486_/Y _6313_/A1 _6315_/S VGND VPWR _7138_/D VGND VPWR sky130_fd_sc_hd__mux2_1
Xhold735 _4176_/X VGND VPWR _6581_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3525_ input16/X _3358_/Y _4202_/A _6608_/Q VGND VPWR _3525_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xhold746 _6825_/Q VGND VPWR hold746/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_517 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold757 _4018_/X VGND VPWR _6458_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold768 _7154_/Q VGND VPWR hold768/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _4036_/X VGND VPWR _6473_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _6702_/Q _5971_/A _5979_/X _6472_/Q VGND VPWR _6244_/X VGND VPWR sky130_fd_sc_hd__a22o_2
X_3456_ _6991_/Q _5436_/A hold76/A _7044_/Q VGND VPWR _3456_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_115_198 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_6175_ _6175_/A _6175_/B _6175_/C _6175_/D VGND VPWR _6176_/D VGND VPWR sky130_fd_sc_hd__nor4_1
X_3387_ _7001_/Q _5445_/A _5373_/A _6937_/Q _3382_/X VGND VPWR _3392_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_561 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1402 _6468_/Q VGND VPWR _4030_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _6577_/Q VGND VPWR hold1413/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _5126_/A _5126_/B _5126_/C VGND VPWR _5126_/X VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1424 _7139_/Q VGND VPWR hold1424/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold1435 _6570_/Q VGND VPWR _4164_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _7133_/Q VGND VPWR _6308_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1457 _3764_/X VGND VPWR _6728_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _6577_/Q VGND VPWR _4171_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _5057_/A _5057_/B _5057_/C VGND VPWR _5126_/A VGND VPWR sky130_fd_sc_hd__and3_1
Xhold1479 _6585_/Q VGND VPWR _4181_/A1 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_288 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_4008_ _4008_/A _4322_/B VGND VPWR _4013_/S VGND VPWR sky130_fd_sc_hd__and2_2
XFILLER_37_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_653 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_185 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A _5981_/A VGND VPWR _5959_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_185_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_714 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_561 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_555 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_237 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_669 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VPWR hold40/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A VGND VPWR hold51/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A VGND VPWR hold62/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_63 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold73 hold73/A VGND VPWR hold73/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_255 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold84 hold84/A VGND VPWR hold84/X VGND VPWR sky130_fd_sc_hd__buf_6
XFILLER_152_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold95 hold95/A VGND VPWR hold95/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_300 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_299 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_543 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_257 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_599 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 _5310_/A VGND VPWR VPWR VGND sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_603 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_474 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3310_ _3374_/A _3370_/A VGND VPWR _5310_/A VGND VPWR sky130_fd_sc_hd__nor2_8
X_4290_ hold377/X _5518_/A1 _4291_/S VGND VPWR _4290_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_98_336 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_281 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_135 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3241_ _7169_/Q _7168_/Q VGND VPWR _3875_/C VGND VPWR sky130_fd_sc_hd__nor2_1
XFILLER_140_455 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_701 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_477 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_3172_ _6485_/Q VGND VPWR _3867_/A VGND VPWR sky130_fd_sc_hd__inv_2
XFILLER_79_583 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_244 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_119 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_737 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6931_ _6963_/CLK _6931_/D fanout458/X VGND VPWR _6931_/Q VGND VPWR sky130_fd_sc_hd__dfstp_1
XFILLER_81_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_642 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6862_ _7079_/CLK _6862_/D fanout480/X VGND VPWR _6862_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_4
XFILLER_179_113 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_601 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
X_5813_ _6969_/Q _5642_/X _5666_/X _6897_/Q VGND VPWR _5813_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_62_494 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_645 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6793_ _7053_/CLK _6793_/D fanout459/X VGND VPWR _6793_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_179_179 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_5744_ _6854_/Q _5648_/X _5666_/X _6894_/Q _5743_/X VGND VPWR _5748_/B VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_533 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_5675_ _6995_/Q _5643_/X _5645_/X _7027_/Q VGND VPWR _5675_/X VGND VPWR sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VPWR _6749_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
X_4626_ _4753_/B _4626_/B VGND VPWR _4626_/Y VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold510 _4242_/X VGND VPWR _6633_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_355 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
X_4557_ _4557_/A VGND VPWR _4967_/A VGND VPWR sky130_fd_sc_hd__inv_2
Xhold521 _6984_/Q VGND VPWR hold521/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _4297_/X VGND VPWR _6689_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_377 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold543 _7064_/Q VGND VPWR hold543/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _5159_/X VGND VPWR _6746_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _5153_/X VGND VPWR _6741_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _7006_/Q _3370_/Y _4292_/A _6689_/Q VGND VPWR _3508_/X VGND VPWR sky130_fd_sc_hd__a22o_2
XFILLER_103_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold576 _6961_/Q VGND VPWR hold576/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _4600_/B _4611_/B VGND VPWR _4672_/B VGND VPWR sky130_fd_sc_hd__nand2_8
Xhold587 _3995_/X VGND VPWR _6438_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_444 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xhold598 _7050_/Q VGND VPWR hold598/X VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6541_/Q _6226_/B _6226_/X VGND VPWR _6227_/X VGND VPWR sky130_fd_sc_hd__o21ba_1
X_3439_ _6920_/Q _5355_/A _5247_/A _6824_/Q _3438_/X VGND VPWR _3446_/A VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XFILLER_103_157 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_701 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
X_6158_ _6865_/Q _5943_/X _5981_/X _6921_/Q VGND VPWR _6158_/X VGND VPWR sky130_fd_sc_hd__a22o_1
XFILLER_112_691 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xhold1210 _5221_/X VGND VPWR _6794_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1221 _6986_/Q VGND VPWR _5437_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk _6601_/CLK VGND VPWR _6655_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
Xhold1232 _5533_/X VGND VPWR _7071_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _6655_/Q VGND VPWR _4257_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _5135_/A _5109_/B _5135_/B VGND VPWR _5109_/Y VGND VPWR sky130_fd_sc_hd__nand3_2
Xhold1254 _5203_/X VGND VPWR _6778_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
X_6089_ _6089_/A _6089_/B _6089_/C VGND VPWR _6089_/Y VGND VPWR sky130_fd_sc_hd__nor3_2
XFILLER_45_417 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xhold1265 _6614_/Q VGND VPWR _4215_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _4305_/X VGND VPWR _6695_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _6450_/Q VGND VPWR _4009_/A0 VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 _4119_/X VGND VPWR _6532_/D VGND VPWR sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_82_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_99 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_csclk clkbuf_3_7_0_csclk/X VGND VPWR _7067_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_196 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_329 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_166 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_546 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_430 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_260 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VPWR _4337_/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_dat_i[18] VGND VPWR _6329_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_dat_i[28] VGND VPWR _6335_/A2 VGND VPWR sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VPWR _6326_/B1 VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_748 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_439 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_225 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_578 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_141 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_433 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_308 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_667 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_628 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_499 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_3790_ _6986_/Q _5436_/A _5145_/A _6735_/Q _3789_/X VGND VPWR _3793_/C VGND VPWR
+ sky130_fd_sc_hd__a221o_1
XPHY_180 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_5460_ hold648/X _5469_/A1 _5462_/S VGND VPWR _5460_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_117_238 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_193 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
X_4411_ _4739_/A _4415_/A VGND VPWR _4959_/A VGND VPWR sky130_fd_sc_hd__and2_1
X_5391_ _5391_/A _5505_/B VGND VPWR _5399_/S VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_99_612 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_388 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7130_ _7130_/CLK _7130_/D fanout486/X VGND VPWR _7130_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
XFILLER_141_720 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_100 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_4342_ _4556_/A _4563_/A VGND VPWR _4753_/B VGND VPWR sky130_fd_sc_hd__nor2_8
XFILLER_99_656 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_241 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_7061_ _7082_/CLK _7061_/D fanout483/X VGND VPWR _7061_/Q VGND VPWR sky130_fd_sc_hd__dfrtp_1
X_4273_ hold227/X hold60/X _4273_/S VGND VPWR _4273_/X VGND VPWR sky130_fd_sc_hd__mux2_1
XFILLER_140_263 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
X_6012_ _6923_/Q _5938_/X _5952_/X _6955_/Q VGND VPWR _6012_/X VGND VPWR sky130_fd_sc_hd__a22o_1
.ends

.subckt buff_flash_clkrst VPWR in_n[0] in_n[10] in_n[11] in_n[1] in_n[2] in_n[3] in_n[4]
+ in_n[5] in_n[6] in_n[7] in_n[8] in_n[9] in_s[0] in_s[1] in_s[2] out_n[0] out_n[1]
+ out_n[2] out_s[0] out_s[10] out_s[11] out_s[1] out_s[2] out_s[3] out_s[4] out_s[5]
+ out_s[6] out_s[7] out_s[8] out_s[9] VGND
XBUF\[10\] in_n[7] VGND VPWR out_s[7] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XBUF\[5\] in_n[2] VGND VPWR out_s[2] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_3_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XBUF\[3\] in_n[0] VGND VPWR out_s[0] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_1_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XBUF\[1\] in_s[1] VGND VPWR out_n[1] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XBUF\[13\] in_n[10] VGND VPWR out_s[10] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XPHY_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XBUF\[8\] in_n[5] VGND VPWR out_s[5] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_1_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_3
XBUF\[6\] in_n[3] VGND VPWR out_s[3] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_1_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XBUF\[11\] in_n[8] VGND VPWR out_s[8] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_4_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XBUF\[4\] in_n[1] VGND VPWR out_s[1] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_2_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XBUF\[2\] in_s[2] VGND VPWR out_n[2] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_2_67 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XBUF\[0\] in_s[0] VGND VPWR out_n[0] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_70 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
XBUF\[9\] in_n[6] VGND VPWR out_s[6] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_2_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XBUF\[14\] in_n[11] VGND VPWR out_s[11] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XFILLER_3_42 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
XBUF\[12\] in_n[9] VGND VPWR out_s[9] VGND VPWR sky130_fd_sc_hd__clkbuf_8
XBUF\[7\] in_n[4] VGND VPWR out_s[4] VGND VPWR sky130_fd_sc_hd__clkbuf_8
.ends

.subckt caravan clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vccd vccd1 vccd2 vdda vdda1 vdda1_2 vdda2 vddio vddio_2 vssa vssa1 vssa1_2
+ vssa2 vssd vssd1 vssd2 vssio vssio_2
Xgpio_control_in_2\[0\] gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[10]
+ gpio_defaults_block_25/gpio_defaults[11] gpio_defaults_block_25/gpio_defaults[12]
+ gpio_defaults_block_25/gpio_defaults[1] gpio_defaults_block_25/gpio_defaults[2]
+ gpio_defaults_block_25/gpio_defaults[3] gpio_defaults_block_25/gpio_defaults[4]
+ gpio_defaults_block_25/gpio_defaults[5] gpio_defaults_block_25/gpio_defaults[6]
+ gpio_defaults_block_25/gpio_defaults[7] gpio_defaults_block_25/gpio_defaults[8]
+ gpio_defaults_block_25/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[7] padframe/mprj_io_one[0]
+ sigbuf/mgmt_io_out_buf[7] padframe/mprj_io_one[0] padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] gpio_control_in_2\[0\]/resetn
+ gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[0\]/serial_clock_out
+ gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out gpio_control_in_2\[0\]/serial_load
+ gpio_control_in_2\[0\]/serial_load_out mprj/io_in[14] mprj/io_oeb[14] mprj/io_out[14]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[0\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_11 soc/VPWR gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_defaults_block_33 soc/VPWR gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_defaults_block_12 soc/VPWR gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_defaults_block_34 soc/VPWR gpio_defaults_block_34/gpio_defaults[0] gpio_defaults_block_34/gpio_defaults[10]
+ gpio_defaults_block_34/gpio_defaults[11] gpio_defaults_block_34/gpio_defaults[12]
+ gpio_defaults_block_34/gpio_defaults[1] gpio_defaults_block_34/gpio_defaults[2]
+ gpio_defaults_block_34/gpio_defaults[3] gpio_defaults_block_34/gpio_defaults[4]
+ gpio_defaults_block_34/gpio_defaults[5] gpio_defaults_block_34/gpio_defaults[6]
+ gpio_defaults_block_34/gpio_defaults[7] gpio_defaults_block_34/gpio_defaults[8]
+ gpio_defaults_block_34/gpio_defaults[9] VSUBS gpio_defaults_block
Xpll soc/VPWR pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3] pll/div[4]
+ pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13]
+ pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18]
+ pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22]
+ pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3]
+ pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8]
+ pll/ext_trim[9] pll/osc pll/resetb pll/clockp[0] VSUBS digital_pll
Xpadframe clock padframe/clock_core padframe/por flash_clk flash_csb flash_io0 padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ieb_core padframe/flash_io0_oeb_core
+ flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ieb_core
+ padframe/flash_io1_oeb_core gpio soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad
+ soc/gpio_out_pad soc/gpio_outenb_pad vccd vdda vddio vddio_2 vssa vssd vssio vssio_2
+ mprj_io[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0] padframe/mprj_io_analog_sel[0]
+ padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2] padframe/mprj_io_holdover[0]
+ padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_inp_dis[0] padframe/mprj_io_oeb[0]
+ padframe/mprj_io_out[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_in[0] mprj/io_in_3v3[0] mprj/gpio_analog[3] mprj/gpio_noesd[3]
+ mprj_io[10] padframe/mprj_io_analog_en[10] padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10]
+ padframe/mprj_io_dm[30] padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10]
+ padframe/mprj_io_ib_mode_sel[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_out[10] padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10]
+ padframe/mprj_io_in[10] mprj/io_in_3v3[10] mprj/gpio_analog[4] mprj/gpio_noesd[4]
+ mprj_io[11] padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11]
+ padframe/mprj_io_dm[33] padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11]
+ padframe/mprj_io_ib_mode_sel[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_out[11] padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11]
+ padframe/mprj_io_in[11] mprj/io_in_3v3[11] mprj/gpio_analog[5] mprj/gpio_noesd[5]
+ mprj_io[12] padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12]
+ padframe/mprj_io_dm[36] padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12]
+ padframe/mprj_io_ib_mode_sel[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_out[12] padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12]
+ padframe/mprj_io_in[12] mprj/io_in_3v3[12] mprj/gpio_analog[6] mprj/gpio_noesd[6]
+ mprj_io[13] padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13]
+ padframe/mprj_io_dm[39] padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13]
+ padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_out[13] padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13]
+ padframe/mprj_io_in[13] mprj/io_in_3v3[13] mprj_io[1] padframe/mprj_io_analog_en[1]
+ padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3]
+ padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_oeb[1] padframe/mprj_io_out[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] padframe/mprj_io_in[1] mprj/io_in_3v3[1] mprj_io[2]
+ padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2] padframe/mprj_io_analog_sel[2]
+ padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8] padframe/mprj_io_holdover[2]
+ padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_inp_dis[2] padframe/mprj_io_oeb[2]
+ padframe/mprj_io_out[2] padframe/mprj_io_slow_sel[2] padframe/mprj_io_vtrip_sel[2]
+ padframe/mprj_io_in[2] mprj/io_in_3v3[2] mprj_io[3] padframe/mprj_io_analog_en[3]
+ padframe/mprj_io_analog_pol[3] padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[10]
+ padframe/mprj_io_dm[11] padframe/mprj_io_dm[9] padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_oeb[3] padframe/mprj_io_out[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] padframe/mprj_io_in[3] mprj/io_in_3v3[3] mprj_io[4]
+ padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4] padframe/mprj_io_analog_sel[4]
+ padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14] padframe/mprj_io_holdover[4]
+ padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_inp_dis[4] padframe/mprj_io_oeb[4]
+ padframe/mprj_io_out[4] padframe/mprj_io_slow_sel[4] padframe/mprj_io_vtrip_sel[4]
+ padframe/mprj_io_in[4] mprj/io_in_3v3[4] mprj_io[5] padframe/mprj_io_analog_en[5]
+ padframe/mprj_io_analog_pol[5] padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15]
+ padframe/mprj_io_dm[16] padframe/mprj_io_dm[17] padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_oeb[5] padframe/mprj_io_out[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] padframe/mprj_io_in[5] mprj/io_in_3v3[5] mprj_io[6]
+ padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6] padframe/mprj_io_analog_sel[6]
+ padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20] padframe/mprj_io_holdover[6]
+ padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_inp_dis[6] padframe/mprj_io_oeb[6]
+ padframe/mprj_io_out[6] padframe/mprj_io_slow_sel[6] padframe/mprj_io_vtrip_sel[6]
+ padframe/mprj_io_in[6] mprj/io_in_3v3[6] mprj/gpio_analog[0] mprj/gpio_noesd[0]
+ mprj_io[7] padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_inp_dis[7] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ padframe/mprj_io_in[7] mprj/io_in_3v3[7] mprj/gpio_analog[1] mprj/gpio_noesd[1]
+ mprj_io[8] padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_inp_dis[8] padframe/mprj_io_oeb[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ padframe/mprj_io_in[8] mprj/io_in_3v3[8] mprj/gpio_analog[2] mprj/gpio_noesd[2]
+ mprj_io[9] padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_inp_dis[9] padframe/mprj_io_oeb[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ padframe/mprj_io_in[9] mprj/io_in_3v3[9] mprj/gpio_analog[7] mprj/gpio_noesd[7]
+ mprj_io[25] padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14]
+ padframe/mprj_io_dm[42] padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14]
+ padframe/mprj_io_ib_mode_sel[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_out[14] padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14]
+ padframe/mprj_io_in[14] mprj/io_in_3v3[14] mprj/gpio_analog[17] mprj/gpio_noesd[17]
+ mprj_io[35] padframe/mprj_io_analog_en[24] padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24]
+ padframe/mprj_io_dm[72] padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24]
+ padframe/mprj_io_ib_mode_sel[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_out[24] padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24]
+ padframe/mprj_io_in[24] mprj/io_in_3v3[24] mprj_io[36] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_inp_dis[25] padframe/mprj_io_oeb[25] padframe/mprj_io_out[25] padframe/mprj_io_slow_sel[25]
+ padframe/mprj_io_vtrip_sel[25] padframe/mprj_io_in[25] mprj/io_in_3v3[25] mprj_io[37]
+ padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26]
+ padframe/mprj_io_dm[78] padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26]
+ padframe/mprj_io_ib_mode_sel[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_out[26] padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26]
+ padframe/mprj_io_in[26] mprj/io_in_3v3[26] mprj/gpio_analog[8] mprj/gpio_noesd[8]
+ mprj_io[26] padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15]
+ padframe/mprj_io_dm[45] padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_out[15] padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_in[15] mprj/io_in_3v3[15] mprj/gpio_analog[9] mprj/gpio_noesd[9]
+ mprj_io[27] padframe/mprj_io_analog_en[16] padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16]
+ padframe/mprj_io_dm[48] padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16]
+ padframe/mprj_io_ib_mode_sel[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_out[16] padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16]
+ padframe/mprj_io_in[16] mprj/io_in_3v3[16] mprj/gpio_analog[10] mprj/gpio_noesd[10]
+ mprj_io[28] padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17]
+ padframe/mprj_io_dm[51] padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17]
+ padframe/mprj_io_ib_mode_sel[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_out[17] padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17]
+ padframe/mprj_io_in[17] mprj/io_in_3v3[17] mprj/gpio_analog[11] mprj/gpio_noesd[11]
+ mprj_io[29] padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18]
+ padframe/mprj_io_dm[54] padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18]
+ padframe/mprj_io_ib_mode_sel[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_out[18] padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18]
+ padframe/mprj_io_in[18] mprj/io_in_3v3[18] mprj/gpio_analog[12] mprj/gpio_noesd[12]
+ mprj_io[30] padframe/mprj_io_analog_en[19] padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19]
+ padframe/mprj_io_dm[57] padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19]
+ padframe/mprj_io_ib_mode_sel[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_out[19] padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19]
+ padframe/mprj_io_in[19] mprj/io_in_3v3[19] mprj/gpio_analog[13] mprj/gpio_noesd[13]
+ mprj_io[31] padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20]
+ padframe/mprj_io_dm[60] padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20]
+ padframe/mprj_io_ib_mode_sel[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_out[20] padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20]
+ padframe/mprj_io_in[20] mprj/io_in_3v3[20] mprj/gpio_analog[14] mprj/gpio_noesd[14]
+ mprj_io[32] padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21]
+ padframe/mprj_io_dm[63] padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21]
+ padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_out[21] padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21]
+ padframe/mprj_io_in[21] mprj/io_in_3v3[21] mprj/gpio_analog[15] mprj/gpio_noesd[15]
+ mprj_io[33] padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22]
+ padframe/mprj_io_dm[66] padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22]
+ padframe/mprj_io_ib_mode_sel[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_out[22] padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22]
+ padframe/mprj_io_in[22] mprj/io_in_3v3[22] mprj/gpio_analog[16] mprj/gpio_noesd[16]
+ mprj_io[34] padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23]
+ padframe/mprj_io_dm[69] padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_out[23] padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_in[23] mprj/io_in_3v3[23] resetb rstb_level/A padframe/vdda mprj/io_analog[1]
+ mprj_io[15] mprj/io_analog[2] mprj_io[16] mprj/io_analog[3] mprj_io[17] mprj/io_analog[0]
+ mprj_io[14] mprj/io_clamp_high[0] mprj_io[18] vccd1 vdda1 vdda1_2 vssa1 vssa1_2
+ mprj/vccd1 mprj/vdda1 mprj/vssd1 vssd1 mprj/io_analog[7] mprj_io[21] mprj/io_analog[8]
+ mprj_io[22] mprj/io_analog[9] mprj_io[23] mprj/io_analog[10] mprj_io[24] mprj/io_analog[5]
+ mprj/io_clamp_high[1] mprj/io_clamp_low[1] mprj_io[19] mprj_io[20] vccd2 vdda2 vssa2
+ mprj/vccd2 mprj/vdda2 mprj/vssd2 vssd2 padframe/flash_csb_core padframe/flash_clk_oeb_core
+ padframe/flash_clk_core padframe/flash_csb_oeb_core padframe/mprj_io_one[0] padframe/mprj_io_one[1]
+ padframe/mprj_io_one[2] padframe/mprj_io_one[3] padframe/mprj_io_one[4] padframe/mprj_io_one[5]
+ padframe/mprj_io_one[6] padframe/mprj_io_one[7] padframe/mprj_io_one[8] padframe/mprj_io_one[9]
+ padframe/mprj_io_one[10] padframe/mprj_io_one[11] padframe/mprj_io_one[12] padframe/mprj_io_one[13]
+ padframe/mprj_io_one[14] padframe/mprj_io_one[15] padframe/mprj_io_one[16] padframe/mprj_io_one[17]
+ padframe/mprj_io_one[18] padframe/mprj_io_one[19] padframe/mprj_io_one[20] padframe/mprj_io_one[21]
+ padframe/mprj_io_one[22] padframe/mprj_io_one[23] padframe/mprj_io_one[24] padframe/mprj_io_one[25]
+ padframe/mprj_io_one[26] por/porb_h soc/gpio_mode1_pad padframe/vssa mprj/io_analog[6]
+ mprj/io_clamp_low[0] mprj/io_clamp_high[2] mprj/io_clamp_low[2] mprj/vssa2 por/vdd3v3
+ mprj/vssa1 VSUBS mprj/io_analog[4] soc/VPWR por/vss3v3 chip_io_alt
Xgpio_defaults_block_13 soc/VPWR gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_1a\[3\] gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] padframe/mprj_io_one[5] housekeeping/mgmt_gpio_out[5]
+ padframe/mprj_io_one[5] padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] soc/VPWR mprj/vccd1 gpio_control_in_1a\[3\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_35 soc/VPWR gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_bidir_2\[0\] gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[17] sigbuf/mgmt_io_oeb_buf[0]
+ sigbuf/mgmt_io_out_buf[17] padframe/mprj_io_one[24] padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] gpio_control_bidir_2\[0\]/resetn
+ gpio_control_in_2\[9\]/resetn gpio_control_bidir_2\[0\]/serial_clock gpio_control_in_2\[9\]/serial_clock
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_in_2\[9\]/serial_data_in gpio_control_bidir_2\[0\]/serial_load
+ gpio_control_in_2\[9\]/serial_load mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24]
+ soc/VPWR mprj/vccd1 gpio_control_bidir_2\[0\]/zero mprj/vssd1 VSUBS gpio_control_block
Xsoc VSUBS soc/VPWR soc/clk_in soc/clk_out soc/clk_in soc/resetn_in soc/debug_in soc/debug_mode
+ soc/debug_oeb soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do
+ soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di
+ soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb
+ soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad
+ soc/gpio_outenb_pad soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11]
+ soc/hk_dat_i[12] soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16]
+ soc/hk_dat_i[17] soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20]
+ soc/hk_dat_i[21] soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25]
+ soc/hk_dat_i[26] soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2]
+ soc/hk_dat_i[30] soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5]
+ soc/hk_dat_i[6] soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] soc/hk_stb_o soc/irq[0]
+ soc/irq[1] soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0] soc/la_iena[100]
+ soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105]
+ soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10]
+ soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114]
+ soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119]
+ soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123]
+ soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12]
+ soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17]
+ soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22]
+ soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27]
+ soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32]
+ soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37]
+ soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42]
+ soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47]
+ soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52]
+ soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57]
+ soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62]
+ soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67]
+ soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72]
+ soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77]
+ soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82]
+ soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87]
+ soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92]
+ soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97]
+ soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] soc/la_input[0] soc/la_input[100]
+ soc/la_input[101] soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105]
+ soc/la_input[106] soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10]
+ soc/la_input[110] soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114]
+ soc/la_input[115] soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119]
+ soc/la_input[11] soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123]
+ soc/la_input[124] soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12]
+ soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17]
+ soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21]
+ soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26]
+ soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30]
+ soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35]
+ soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3]
+ soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44]
+ soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49]
+ soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53]
+ soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58]
+ soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62]
+ soc/la_input[63] soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67]
+ soc/la_input[68] soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71]
+ soc/la_input[72] soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76]
+ soc/la_input[77] soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80]
+ soc/la_input[81] soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85]
+ soc/la_input[86] soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8]
+ soc/la_input[90] soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94]
+ soc/la_input[95] soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99]
+ soc/la_input[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102]
+ soc/la_output[103] soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107]
+ soc/la_output[108] soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111]
+ soc/la_output[112] soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116]
+ soc/la_output[117] soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120]
+ soc/la_output[121] soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125]
+ soc/la_output[126] soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14]
+ soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19]
+ soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23]
+ soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28]
+ soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32]
+ soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37]
+ soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41]
+ soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46]
+ soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50]
+ soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55]
+ soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5]
+ soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64]
+ soc/la_output[65] soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69]
+ soc/la_output[6] soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73]
+ soc/la_output[74] soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78]
+ soc/la_output[79] soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82]
+ soc/la_output[83] soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87]
+ soc/la_output[88] soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91]
+ soc/la_output[92] soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96]
+ soc/la_output[97] soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/mprj_ack_i
+ soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13]
+ soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18]
+ soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22]
+ soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27]
+ soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31]
+ soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7]
+ soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0] soc/mprj_dat_i[10]
+ soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15]
+ soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1]
+ soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24]
+ soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29]
+ soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4]
+ soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9]
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2]
+ soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_wb_iena soc/mprj_we_o por/por_l padframe/por
+ por/por_l soc/porb_h_out soc/qspi_enabled soc/resetn_in soc/resetn_out rstb_level/X
+ pll/resetb soc/ser_rx soc/ser_tx soc/serial_clock_in soc/serial_clock_out soc/serial_data_2_in
+ soc/serial_data_2_out soc/serial_load_in soc/serial_load_out soc/serial_resetn_in
+ soc/serial_resetn_out soc/spi_csb soc/spi_enabled soc/spi_sck soc/spi_sdi soc/spi_sdo
+ soc/spi_sdoenb soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1]
+ soc/user_irq_ena[2] mgmt_core_wrapper
Xgpio_defaults_block_25 soc/VPWR gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[10]
+ gpio_defaults_block_25/gpio_defaults[11] gpio_defaults_block_25/gpio_defaults[12]
+ gpio_defaults_block_25/gpio_defaults[1] gpio_defaults_block_25/gpio_defaults[2]
+ gpio_defaults_block_25/gpio_defaults[3] gpio_defaults_block_25/gpio_defaults[4]
+ gpio_defaults_block_25/gpio_defaults[5] gpio_defaults_block_25/gpio_defaults[6]
+ gpio_defaults_block_25/gpio_defaults[7] gpio_defaults_block_25/gpio_defaults[8]
+ gpio_defaults_block_25/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_2\[9\] gpio_defaults_block_34/gpio_defaults[0] gpio_defaults_block_34/gpio_defaults[10]
+ gpio_defaults_block_34/gpio_defaults[11] gpio_defaults_block_34/gpio_defaults[12]
+ gpio_defaults_block_34/gpio_defaults[1] gpio_defaults_block_34/gpio_defaults[2]
+ gpio_defaults_block_34/gpio_defaults[3] gpio_defaults_block_34/gpio_defaults[4]
+ gpio_defaults_block_34/gpio_defaults[5] gpio_defaults_block_34/gpio_defaults[6]
+ gpio_defaults_block_34/gpio_defaults[7] gpio_defaults_block_34/gpio_defaults[8]
+ gpio_defaults_block_34/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[16] padframe/mprj_io_one[9]
+ sigbuf/mgmt_io_out_buf[16] padframe/mprj_io_one[9] padframe/mprj_io_analog_en[23]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69]
+ padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[8\]/resetn gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load
+ gpio_control_in_2\[8\]/serial_load mprj/io_in[23] mprj/io_oeb[23] mprj/io_out[23]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[9\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_36 soc/VPWR gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_defaults_block_26 soc/VPWR gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_1\[4\] gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[5] padframe/mprj_io_one[12]
+ sigbuf/mgmt_io_out_buf[5] padframe/mprj_io_one[12] padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[5\]/resetn gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load
+ gpio_control_in_1\[5\]/serial_load mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12]
+ soc/VPWR mprj/vccd1 gpio_control_in_1\[4\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_37 soc/VPWR gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] VSUBS gpio_defaults_block
Xpor por/vdd3v3 soc/VPWR por/porb_h por/por_l por/porb_l VSUBS por/vss3v3 simple_por
Xgpio_defaults_block_27 soc/VPWR gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_1a\[1\] gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[3] padframe/mprj_io_one[3] housekeeping/mgmt_gpio_out[3]
+ padframe/mprj_io_one[3] padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[1\]/serial_data_in
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load gpio_control_in_1a\[2\]/serial_load
+ mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3] soc/VPWR mprj/vccd1 gpio_control_in_1a\[1\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xclock_ctrl clock_ctrl/core_clk pll/osc clock_ctrl/ext_clk_sel housekeeping/reset
+ pll/clockp[1] pll/clockp[0] pll/resetb housekeeping/wb_rstn_i clock_ctrl/sel2[0]
+ clock_ctrl/sel2[1] clock_ctrl/sel2[2] clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2]
+ clock_ctrl/user_clk VSUBS soc/VPWR caravel_clocking
Xgpio_defaults_block_28 soc/VPWR gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_2\[7\] gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[14] padframe/mprj_io_one[7]
+ sigbuf/mgmt_io_out_buf[14] padframe/mprj_io_one[7] padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63]
+ padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[6\]/resetn gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load
+ gpio_control_in_2\[6\]/serial_load mprj/io_in[21] mprj/io_oeb[21] mprj/io_out[21]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[7\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_29 soc/VPWR gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_1\[2\] gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[3] padframe/mprj_io_one[10]
+ sigbuf/mgmt_io_out_buf[3] padframe/mprj_io_one[10] padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[3\]/resetn gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load
+ gpio_control_in_1\[3\]/serial_load mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10]
+ soc/VPWR mprj/vccd1 gpio_control_in_1\[2\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1\[0\] gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[1] padframe/mprj_io_one[8] sigbuf/mgmt_io_out_buf[1] padframe/mprj_io_one[8]
+ padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8] padframe/mprj_io_inp_dis[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn gpio_control_in_1\[0\]/serial_clock
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load mprj/io_in[8]
+ mprj/io_oeb[8] mprj/io_out[8] soc/VPWR mprj/vccd1 gpio_control_in_1\[0\]/zero mprj/vssd1
+ VSUBS gpio_control_block
Xgpio_control_in_2\[5\] gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[12] padframe/mprj_io_one[5]
+ sigbuf/mgmt_io_out_buf[12] padframe/mprj_io_one[5] padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load
+ gpio_control_in_2\[4\]/serial_load mprj/io_in[19] mprj/io_oeb[19] mprj/io_out[19]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[5\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_0 soc/VPWR gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xspare_logic\[3\] spare_logic\[3\]/spare_xfq[0] spare_logic\[3\]/spare_xfq[1] spare_logic\[3\]/spare_xfqn[0]
+ spare_logic\[3\]/spare_xfqn[1] spare_logic\[3\]/spare_xi[0] spare_logic\[3\]/spare_xi[1]
+ spare_logic\[3\]/spare_xi[2] spare_logic\[3\]/spare_xi[3] spare_logic\[3\]/spare_xib
+ spare_logic\[3\]/spare_xmx[0] spare_logic\[3\]/spare_xmx[1] spare_logic\[3\]/spare_xna[0]
+ spare_logic\[3\]/spare_xna[1] spare_logic\[3\]/spare_xno[0] spare_logic\[3\]/spare_xno[1]
+ spare_logic\[3\]/spare_xz[0] spare_logic\[3\]/spare_xz[10] spare_logic\[3\]/spare_xz[11]
+ spare_logic\[3\]/spare_xz[12] spare_logic\[3\]/spare_xz[13] spare_logic\[3\]/spare_xz[14]
+ spare_logic\[3\]/spare_xz[15] spare_logic\[3\]/spare_xz[16] spare_logic\[3\]/spare_xz[17]
+ spare_logic\[3\]/spare_xz[18] spare_logic\[3\]/spare_xz[19] spare_logic\[3\]/spare_xz[1]
+ spare_logic\[3\]/spare_xz[20] spare_logic\[3\]/spare_xz[21] spare_logic\[3\]/spare_xz[22]
+ spare_logic\[3\]/spare_xz[23] spare_logic\[3\]/spare_xz[24] spare_logic\[3\]/spare_xz[25]
+ spare_logic\[3\]/spare_xz[26] spare_logic\[3\]/spare_xz[2] spare_logic\[3\]/spare_xz[3]
+ spare_logic\[3\]/spare_xz[4] spare_logic\[3\]/spare_xz[5] spare_logic\[3\]/spare_xz[6]
+ spare_logic\[3\]/spare_xz[7] spare_logic\[3\]/spare_xz[8] spare_logic\[3\]/spare_xz[9]
+ soc/VPWR VSUBS spare_logic_block
Xgpio_defaults_block_1 soc/VPWR gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ soc/VPWR VSUBS user_id_programming
Xgpio_control_in_2\[3\] gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[10] padframe/mprj_io_one[3]
+ sigbuf/mgmt_io_out_buf[10] padframe/mprj_io_one[3] padframe/mprj_io_analog_en[17]
+ padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51]
+ padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] gpio_control_in_2\[3\]/resetn
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[3\]/serial_load
+ gpio_control_in_2\[2\]/serial_load mprj/io_in[17] mprj/io_oeb[17] mprj/io_out[17]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[3\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_2 soc/VPWR gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_defaults_block_3 soc/VPWR gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_control_bidir_1\[0\] gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_out[0]
+ padframe/mprj_io_one[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0]
+ padframe/mprj_io_inp_dis[0] padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0]
+ padframe/mprj_io_vtrip_sel[0] soc/serial_resetn_in gpio_control_bidir_1\[1\]/resetn
+ soc/serial_clock_in gpio_control_bidir_1\[1\]/serial_clock housekeeping/serial_data_1
+ gpio_control_bidir_1\[1\]/serial_data_in soc/serial_load_in gpio_control_bidir_1\[1\]/serial_load
+ mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0] soc/VPWR mprj/vccd1 gpio_control_bidir_1\[0\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_5 soc/VPWR gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_defaults_block_4 soc/VPWR gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xspare_logic\[1\] spare_logic\[1\]/spare_xfq[0] spare_logic\[1\]/spare_xfq[1] spare_logic\[1\]/spare_xfqn[0]
+ spare_logic\[1\]/spare_xfqn[1] spare_logic\[1\]/spare_xi[0] spare_logic\[1\]/spare_xi[1]
+ spare_logic\[1\]/spare_xi[2] spare_logic\[1\]/spare_xi[3] spare_logic\[1\]/spare_xib
+ spare_logic\[1\]/spare_xmx[0] spare_logic\[1\]/spare_xmx[1] spare_logic\[1\]/spare_xna[0]
+ spare_logic\[1\]/spare_xna[1] spare_logic\[1\]/spare_xno[0] spare_logic\[1\]/spare_xno[1]
+ spare_logic\[1\]/spare_xz[0] spare_logic\[1\]/spare_xz[10] spare_logic\[1\]/spare_xz[11]
+ spare_logic\[1\]/spare_xz[12] spare_logic\[1\]/spare_xz[13] spare_logic\[1\]/spare_xz[14]
+ spare_logic\[1\]/spare_xz[15] spare_logic\[1\]/spare_xz[16] spare_logic\[1\]/spare_xz[17]
+ spare_logic\[1\]/spare_xz[18] spare_logic\[1\]/spare_xz[19] spare_logic\[1\]/spare_xz[1]
+ spare_logic\[1\]/spare_xz[20] spare_logic\[1\]/spare_xz[21] spare_logic\[1\]/spare_xz[22]
+ spare_logic\[1\]/spare_xz[23] spare_logic\[1\]/spare_xz[24] spare_logic\[1\]/spare_xz[25]
+ spare_logic\[1\]/spare_xz[26] spare_logic\[1\]/spare_xz[2] spare_logic\[1\]/spare_xz[3]
+ spare_logic\[1\]/spare_xz[4] spare_logic\[1\]/spare_xz[5] spare_logic\[1\]/spare_xz[6]
+ spare_logic\[1\]/spare_xz[7] spare_logic\[1\]/spare_xz[8] spare_logic\[1\]/spare_xz[9]
+ soc/VPWR VSUBS spare_logic_block
Xgpio_control_in_2\[1\] gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[8] padframe/mprj_io_one[1]
+ sigbuf/mgmt_io_out_buf[8] padframe/mprj_io_one[1] padframe/mprj_io_analog_en[15]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45]
+ padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] gpio_control_in_2\[1\]/resetn
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[1\]/serial_load
+ gpio_control_in_2\[0\]/serial_load mprj/io_in[15] mprj/io_oeb[15] mprj/io_out[15]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[1\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_6 soc/VPWR gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_defaults_block_7 soc/VPWR gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xsigbuf sigbuf/mgmt_io_in_unbuf[6] sigbuf/mgmt_io_out_buf[6] sigbuf/mgmt_io_in_unbuf[5]
+ sigbuf/mgmt_io_in_unbuf[4] sigbuf/mgmt_io_in_unbuf[3] sigbuf/mgmt_io_in_unbuf[2]
+ sigbuf/mgmt_io_in_unbuf[1] sigbuf/mgmt_io_in_unbuf[0] sigbuf/mgmt_io_out_buf[0]
+ sigbuf/mgmt_io_out_buf[1] sigbuf/mgmt_io_out_buf[2] sigbuf/mgmt_io_out_buf[3] sigbuf/mgmt_io_out_buf[4]
+ sigbuf/mgmt_io_out_buf[5] sigbuf/mgmt_io_out_unbuf[0] sigbuf/mgmt_io_out_unbuf[1]
+ sigbuf/mgmt_io_out_unbuf[2] sigbuf/mgmt_io_out_unbuf[3] sigbuf/mgmt_io_out_unbuf[4]
+ sigbuf/mgmt_io_out_unbuf[5] sigbuf/mgmt_io_out_unbuf[6] sigbuf/mgmt_io_in_buf[6]
+ sigbuf/mgmt_io_in_buf[5] sigbuf/mgmt_io_in_buf[4] sigbuf/mgmt_io_in_buf[3] sigbuf/mgmt_io_in_buf[2]
+ sigbuf/mgmt_io_in_buf[1] sigbuf/mgmt_io_in_buf[0] sigbuf/mgmt_io_out_buf[10] sigbuf/mgmt_io_out_buf[11]
+ sigbuf/mgmt_io_in_unbuf[11] sigbuf/mgmt_io_in_unbuf[10] sigbuf/mgmt_io_out_buf[12]
+ sigbuf/mgmt_io_out_buf[13] sigbuf/mgmt_io_out_buf[14] sigbuf/mgmt_io_out_buf[15]
+ sigbuf/mgmt_io_in_unbuf[15] sigbuf/mgmt_io_in_unbuf[14] sigbuf/mgmt_io_in_unbuf[13]
+ sigbuf/mgmt_io_in_unbuf[12] sigbuf/mgmt_io_out_buf[16] sigbuf/mgmt_io_out_buf[17]
+ sigbuf/mgmt_io_out_buf[18] sigbuf/mgmt_io_out_buf[19] sigbuf/mgmt_io_in_unbuf[19]
+ sigbuf/mgmt_io_in_unbuf[18] sigbuf/mgmt_io_in_unbuf[17] sigbuf/mgmt_io_in_unbuf[16]
+ sigbuf/mgmt_io_oeb_buf[0] sigbuf/mgmt_io_oeb_buf[1] sigbuf/mgmt_io_oeb_buf[2] sigbuf/mgmt_io_oeb_unbuf[2]
+ sigbuf/mgmt_io_oeb_unbuf[1] sigbuf/mgmt_io_oeb_unbuf[0] sigbuf/mgmt_io_in_buf[19]
+ sigbuf/mgmt_io_in_buf[18] sigbuf/mgmt_io_in_buf[17] sigbuf/mgmt_io_in_buf[16] sigbuf/mgmt_io_out_unbuf[16]
+ sigbuf/mgmt_io_out_unbuf[17] sigbuf/mgmt_io_out_unbuf[18] sigbuf/mgmt_io_out_unbuf[19]
+ sigbuf/mgmt_io_out_unbuf[15] sigbuf/mgmt_io_out_unbuf[14] sigbuf/mgmt_io_out_unbuf[13]
+ sigbuf/mgmt_io_out_unbuf[12] sigbuf/mgmt_io_out_unbuf[11] sigbuf/mgmt_io_out_unbuf[10]
+ sigbuf/mgmt_io_out_unbuf[9] sigbuf/mgmt_io_out_unbuf[8] sigbuf/mgmt_io_out_unbuf[7]
+ sigbuf/mgmt_io_in_buf[7] sigbuf/mgmt_io_in_buf[8] sigbuf/mgmt_io_in_buf[9] sigbuf/mgmt_io_in_buf[10]
+ sigbuf/mgmt_io_in_buf[11] sigbuf/mgmt_io_in_buf[12] sigbuf/mgmt_io_in_buf[13] sigbuf/mgmt_io_in_buf[14]
+ sigbuf/mgmt_io_in_buf[15] soc/VPWR sigbuf/mgmt_io_out_buf[9] sigbuf/mgmt_io_in_unbuf[9]
+ sigbuf/mgmt_io_out_buf[8] sigbuf/mgmt_io_in_unbuf[8] sigbuf/mgmt_io_out_buf[7] sigbuf/mgmt_io_in_unbuf[7]
+ VSUBS gpio_signal_buffering_alt
Xgpio_defaults_block_8 soc/VPWR gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_control_in_1a\[4\] gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] padframe/mprj_io_one[6] housekeeping/mgmt_gpio_out[6]
+ padframe/mprj_io_one[6] padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] soc/VPWR mprj/vccd1 gpio_control_in_1a\[4\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xmgmt_buffers soc/clk_out clock_ctrl/user_clk soc/resetn_out mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102]
+ mprj/la_data_out[103] mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106]
+ mprj/la_data_out[107] mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10]
+ mprj/la_data_out[110] mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113]
+ mprj/la_data_out[114] mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117]
+ mprj/la_data_out[118] mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120]
+ mprj/la_data_out[121] mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124]
+ mprj/la_data_out[125] mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[64] mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67]
+ mprj/la_data_out[68] mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70]
+ mprj/la_data_out[71] mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74]
+ mprj/la_data_out[75] mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78]
+ mprj/la_data_out[79] mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81]
+ mprj/la_data_out[82] mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85]
+ mprj/la_data_out[86] mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89]
+ mprj/la_data_out[8] mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92]
+ mprj/la_data_out[93] mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96]
+ mprj/la_data_out[97] mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103]
+ soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108]
+ soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112]
+ soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117]
+ soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121]
+ soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126]
+ soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15]
+ soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1]
+ soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24]
+ soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29]
+ soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33]
+ soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38]
+ soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42]
+ soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47]
+ soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51]
+ soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56]
+ soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60]
+ soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65]
+ soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6]
+ soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74]
+ soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79]
+ soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83]
+ soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88]
+ soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92]
+ soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97]
+ soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/la_iena[0] soc/la_iena[100]
+ soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105]
+ soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10]
+ soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114]
+ soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119]
+ soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123]
+ soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12]
+ soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17]
+ soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22]
+ soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27]
+ soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32]
+ soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37]
+ soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42]
+ soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47]
+ soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52]
+ soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57]
+ soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62]
+ soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67]
+ soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72]
+ soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77]
+ soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82]
+ soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87]
+ soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92]
+ soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97]
+ soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[100]
+ mprj/la_oenb[101] mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105]
+ mprj/la_oenb[106] mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10]
+ mprj/la_oenb[110] mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114]
+ mprj/la_oenb[115] mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119]
+ mprj/la_oenb[11] mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123]
+ mprj/la_oenb[124] mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67]
+ mprj/la_oenb[68] mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71]
+ mprj/la_oenb[72] mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76]
+ mprj/la_oenb[77] mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80]
+ mprj/la_oenb[81] mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85]
+ mprj/la_oenb[86] mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8]
+ mprj/la_oenb[90] mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94]
+ mprj/la_oenb[95] mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13]
+ mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18]
+ mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22]
+ mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27]
+ mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31]
+ mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7]
+ mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o mprj/wbs_cyc_i soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11] mprj/wbs_dat_o[12]
+ mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16] mprj/wbs_dat_o[17]
+ mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20] mprj/wbs_dat_o[21]
+ mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25] mprj/wbs_dat_o[26]
+ mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2] mprj/wbs_dat_o[30]
+ mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5] mprj/wbs_dat_o[6]
+ mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_wb_iena soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2]
+ mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i soc/mprj_we_o mprj/wbs_we_i housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1] soc/irq[2] mprj/user_irq[0]
+ mprj/user_irq[1] mprj/user_irq[2] soc/user_irq_ena[0] soc/user_irq_ena[1] soc/user_irq_ena[2]
+ mprj/wb_rst_i mprj/vccd1 mprj/vccd2 mprj/vdda1 mprj/vdda2 mprj/vssa2 mprj/vssa1
+ mprj/vssd2 VSUBS mprj/vssd1 soc/VPWR mgmt_protect
Xrstb_level rstb_level/A rstb_level/X por/vdd3v3 por/vss3v3 soc/VPWR VSUBS xres_buf
Xgpio_defaults_block_9 soc/VPWR gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ VSUBS gpio_defaults_block
Xgpio_control_bidir_2\[1\] gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[18] sigbuf/mgmt_io_oeb_buf[1]
+ sigbuf/mgmt_io_out_buf[18] padframe/mprj_io_one[25] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] gpio_control_bidir_2\[1\]/resetn
+ gpio_control_bidir_2\[0\]/resetn gpio_control_bidir_2\[1\]/serial_clock gpio_control_bidir_2\[0\]/serial_clock
+ gpio_control_bidir_2\[1\]/serial_data_in gpio_control_bidir_2\[0\]/serial_data_in
+ gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load mprj/io_in[25]
+ mprj/io_oeb[25] mprj/io_out[25] soc/VPWR mprj/vccd1 gpio_control_bidir_2\[1\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1\[5\] gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[6] padframe/mprj_io_one[13]
+ sigbuf/mgmt_io_out_buf[6] padframe/mprj_io_one[13] padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[5\]/resetn_out gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[5\]/serial_clock_out
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[5\]/serial_data_out gpio_control_in_1\[5\]/serial_load
+ gpio_control_in_1\[5\]/serial_load_out mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13]
+ soc/VPWR mprj/vccd1 gpio_control_in_1\[5\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1a\[2\] gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[4] padframe/mprj_io_one[4] housekeeping/mgmt_gpio_out[4]
+ padframe/mprj_io_one[4] padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[3\]/resetn
+ gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[2\]/serial_data_in
+ gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load gpio_control_in_1a\[3\]/serial_load
+ mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4] soc/VPWR mprj/vccd1 gpio_control_in_1a\[2\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_2\[8\] gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[15] padframe/mprj_io_one[8]
+ sigbuf/mgmt_io_out_buf[15] padframe/mprj_io_one[8] padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[7\]/resetn gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load
+ gpio_control_in_2\[7\]/serial_load mprj/io_in[22] mprj/io_oeb[22] mprj/io_out[22]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[8\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1\[3\] gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[4] padframe/mprj_io_one[11]
+ sigbuf/mgmt_io_out_buf[4] padframe/mprj_io_one[11] padframe/mprj_io_analog_en[11]
+ padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33]
+ padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[4\]/resetn gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load
+ gpio_control_in_1\[4\]/serial_load mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11]
+ soc/VPWR mprj/vccd1 gpio_control_in_1\[3\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1a\[0\] gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[2] padframe/mprj_io_one[2] housekeeping/mgmt_gpio_out[2]
+ padframe/mprj_io_one[2] padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] gpio_control_in_1a\[0\]/resetn gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load gpio_control_in_1a\[1\]/serial_load
+ mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2] soc/VPWR mprj/vccd1 gpio_control_in_1a\[0\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_2\[6\] gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[13] padframe/mprj_io_one[6]
+ sigbuf/mgmt_io_out_buf[13] padframe/mprj_io_one[6] padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[5\]/resetn gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load
+ gpio_control_in_2\[5\]/serial_load mprj/io_in[20] mprj/io_oeb[20] mprj/io_out[20]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[6\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_in_1\[1\] gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[2] padframe/mprj_io_one[9] sigbuf/mgmt_io_out_buf[2] padframe/mprj_io_one[9]
+ padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9] padframe/mprj_io_inp_dis[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn gpio_control_in_1\[1\]/serial_clock
+ gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[2\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load mprj/io_in[9]
+ mprj/io_oeb[9] mprj/io_out[9] soc/VPWR mprj/vccd1 gpio_control_in_1\[1\]/zero mprj/vssd1
+ VSUBS gpio_control_block
Xmprj mprj/gpio_analog[0] mprj/gpio_analog[10] mprj/gpio_analog[11] mprj/gpio_analog[12]
+ mprj/gpio_analog[13] mprj/gpio_analog[14] mprj/gpio_analog[15] mprj/gpio_analog[16]
+ mprj/gpio_analog[17] mprj/gpio_analog[1] mprj/gpio_analog[2] mprj/gpio_analog[3]
+ mprj/gpio_analog[4] mprj/gpio_analog[5] mprj/gpio_analog[6] mprj/gpio_analog[7]
+ mprj/gpio_analog[8] mprj/gpio_analog[9] mprj/gpio_noesd[0] mprj/gpio_noesd[10] mprj/gpio_noesd[11]
+ mprj/gpio_noesd[12] mprj/gpio_noesd[13] mprj/gpio_noesd[14] mprj/gpio_noesd[15]
+ mprj/gpio_noesd[16] mprj/gpio_noesd[17] mprj/gpio_noesd[1] mprj/gpio_noesd[2] mprj/gpio_noesd[3]
+ mprj/gpio_noesd[4] mprj/gpio_noesd[5] mprj/gpio_noesd[6] mprj/gpio_noesd[7] mprj/gpio_noesd[8]
+ mprj/gpio_noesd[9] mprj/io_analog[0] mprj/io_analog[10] mprj/io_analog[1] mprj/io_analog[2]
+ mprj/io_analog[3] mprj/io_analog[7] mprj/io_analog[8] mprj/io_analog[9] mprj/io_analog[4]
+ mprj/io_analog[5] mprj/io_analog[6] mprj/io_clamp_high[0] mprj/io_clamp_high[1]
+ mprj/io_clamp_high[2] mprj/io_clamp_low[0] mprj/io_clamp_low[1] mprj/io_clamp_low[2]
+ mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14]
+ mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1]
+ mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25]
+ mprj/io_in[26] mprj/io_in[2] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6]
+ mprj/io_in[7] mprj/io_in[8] mprj/io_in[9] mprj/io_in_3v3[0] mprj/io_in_3v3[10] mprj/io_in_3v3[11]
+ mprj/io_in_3v3[12] mprj/io_in_3v3[13] mprj/io_in_3v3[14] mprj/io_in_3v3[15] mprj/io_in_3v3[16]
+ mprj/io_in_3v3[17] mprj/io_in_3v3[18] mprj/io_in_3v3[19] mprj/io_in_3v3[1] mprj/io_in_3v3[20]
+ mprj/io_in_3v3[21] mprj/io_in_3v3[22] mprj/io_in_3v3[23] mprj/io_in_3v3[24] mprj/io_in_3v3[25]
+ mprj/io_in_3v3[26] mprj/io_in_3v3[2] mprj/io_in_3v3[3] mprj/io_in_3v3[4] mprj/io_in_3v3[5]
+ mprj/io_in_3v3[6] mprj/io_in_3v3[7] mprj/io_in_3v3[8] mprj/io_in_3v3[9] mprj/io_oeb[0]
+ mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12] mprj/io_oeb[13] mprj/io_oeb[14]
+ mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17] mprj/io_oeb[18] mprj/io_oeb[19]
+ mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22] mprj/io_oeb[23] mprj/io_oeb[24]
+ mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[2] mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5]
+ mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10]
+ mprj/io_out[11] mprj/io_out[12] mprj/io_out[13] mprj/io_out[14] mprj/io_out[15]
+ mprj/io_out[16] mprj/io_out[17] mprj/io_out[18] mprj/io_out[19] mprj/io_out[1] mprj/io_out[20]
+ mprj/io_out[21] mprj/io_out[22] mprj/io_out[23] mprj/io_out[24] mprj/io_out[25]
+ mprj/io_out[26] mprj/io_out[2] mprj/io_out[3] mprj/io_out[4] mprj/io_out[5] mprj/io_out[6]
+ mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[100]
+ mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103] mprj/la_data_out[104]
+ mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107] mprj/la_data_out[108]
+ mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110] mprj/la_data_out[111]
+ mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114] mprj/la_data_out[115]
+ mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118] mprj/la_data_out[119]
+ mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121] mprj/la_data_out[122]
+ mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125] mprj/la_data_out[126]
+ mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14]
+ mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18]
+ mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21]
+ mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25]
+ mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29]
+ mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32]
+ mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36]
+ mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3]
+ mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43]
+ mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47]
+ mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50]
+ mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54]
+ mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58]
+ mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61]
+ mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64] mprj/la_data_out[65]
+ mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68] mprj/la_data_out[69]
+ mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71] mprj/la_data_out[72]
+ mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75] mprj/la_data_out[76]
+ mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79] mprj/la_data_out[7]
+ mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82] mprj/la_data_out[83]
+ mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86] mprj/la_data_out[87]
+ mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8] mprj/la_data_out[90]
+ mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93] mprj/la_data_out[94]
+ mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97] mprj/la_data_out[98]
+ mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[100] mprj/la_oenb[101]
+ mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105] mprj/la_oenb[106]
+ mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10] mprj/la_oenb[110]
+ mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114] mprj/la_oenb[115]
+ mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119] mprj/la_oenb[11]
+ mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123] mprj/la_oenb[124]
+ mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12] mprj/la_oenb[13]
+ mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17] mprj/la_oenb[18]
+ mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21] mprj/la_oenb[22]
+ mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26] mprj/la_oenb[27]
+ mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30] mprj/la_oenb[31]
+ mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35] mprj/la_oenb[36]
+ mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3] mprj/la_oenb[40]
+ mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44] mprj/la_oenb[45]
+ mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49] mprj/la_oenb[4]
+ mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53] mprj/la_oenb[54]
+ mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58] mprj/la_oenb[59]
+ mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62] mprj/la_oenb[63]
+ mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67] mprj/la_oenb[68]
+ mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71] mprj/la_oenb[72]
+ mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76] mprj/la_oenb[77]
+ mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80] mprj/la_oenb[81]
+ mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85] mprj/la_oenb[86]
+ mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8] mprj/la_oenb[90]
+ mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94] mprj/la_oenb[95]
+ mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] mprj/vccd1 mprj/vccd2
+ mprj/vdda1 mprj/vdda2 mprj/vssa1 mprj/vssa2 mprj/vssd1 mprj/vssd2 mprj/wb_clk_i
+ mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11]
+ mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16]
+ mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20]
+ mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25]
+ mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2]
+ mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5]
+ mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i
+ user_analog_project_wrapper
Xgpio_control_in_2\[4\] gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[11] padframe/mprj_io_one[4]
+ sigbuf/mgmt_io_out_buf[11] padframe/mprj_io_one[4] padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[4\]/serial_load
+ gpio_control_in_2\[3\]/serial_load mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[4\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_control_bidir_1\[1\] gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_out[1]
+ padframe/mprj_io_one[1] padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5]
+ padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] gpio_control_bidir_1\[1\]/resetn gpio_control_in_1a\[0\]/resetn
+ gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock gpio_control_bidir_1\[1\]/serial_data_in
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load
+ mprj/io_in[1] mprj/io_oeb[1] mprj/io_out[1] soc/VPWR mprj/vccd1 gpio_control_bidir_1\[1\]/zero
+ mprj/vssd1 VSUBS gpio_control_block
Xspare_logic\[2\] spare_logic\[2\]/spare_xfq[0] spare_logic\[2\]/spare_xfq[1] spare_logic\[2\]/spare_xfqn[0]
+ spare_logic\[2\]/spare_xfqn[1] spare_logic\[2\]/spare_xi[0] spare_logic\[2\]/spare_xi[1]
+ spare_logic\[2\]/spare_xi[2] spare_logic\[2\]/spare_xi[3] spare_logic\[2\]/spare_xib
+ spare_logic\[2\]/spare_xmx[0] spare_logic\[2\]/spare_xmx[1] spare_logic\[2\]/spare_xna[0]
+ spare_logic\[2\]/spare_xna[1] spare_logic\[2\]/spare_xno[0] spare_logic\[2\]/spare_xno[1]
+ spare_logic\[2\]/spare_xz[0] spare_logic\[2\]/spare_xz[10] spare_logic\[2\]/spare_xz[11]
+ spare_logic\[2\]/spare_xz[12] spare_logic\[2\]/spare_xz[13] spare_logic\[2\]/spare_xz[14]
+ spare_logic\[2\]/spare_xz[15] spare_logic\[2\]/spare_xz[16] spare_logic\[2\]/spare_xz[17]
+ spare_logic\[2\]/spare_xz[18] spare_logic\[2\]/spare_xz[19] spare_logic\[2\]/spare_xz[1]
+ spare_logic\[2\]/spare_xz[20] spare_logic\[2\]/spare_xz[21] spare_logic\[2\]/spare_xz[22]
+ spare_logic\[2\]/spare_xz[23] spare_logic\[2\]/spare_xz[24] spare_logic\[2\]/spare_xz[25]
+ spare_logic\[2\]/spare_xz[26] spare_logic\[2\]/spare_xz[2] spare_logic\[2\]/spare_xz[3]
+ spare_logic\[2\]/spare_xz[4] spare_logic\[2\]/spare_xz[5] spare_logic\[2\]/spare_xz[6]
+ spare_logic\[2\]/spare_xz[7] spare_logic\[2\]/spare_xz[8] spare_logic\[2\]/spare_xz[9]
+ soc/VPWR VSUBS spare_logic_block
Xhousekeeping soc/VPWR soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out soc/irq[3]
+ soc/irq[4] soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ housekeeping/mgmt_gpio_in[0] sigbuf/mgmt_io_in_buf[3] sigbuf/mgmt_io_in_buf[4] sigbuf/mgmt_io_in_buf[5]
+ sigbuf/mgmt_io_in_buf[6] housekeeping/mgmt_gpio_in[14] housekeeping/mgmt_gpio_in[15]
+ housekeeping/mgmt_gpio_in[16] housekeeping/mgmt_gpio_in[17] housekeeping/mgmt_gpio_in[18]
+ housekeeping/mgmt_gpio_in[19] housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_in[20]
+ housekeeping/mgmt_gpio_in[21] housekeeping/mgmt_gpio_in[22] housekeeping/mgmt_gpio_in[23]
+ housekeeping/mgmt_gpio_in[24] sigbuf/mgmt_io_in_buf[7] sigbuf/mgmt_io_in_buf[8]
+ sigbuf/mgmt_io_in_buf[9] sigbuf/mgmt_io_in_buf[10] sigbuf/mgmt_io_in_buf[11] housekeeping/mgmt_gpio_in[2]
+ sigbuf/mgmt_io_in_buf[12] sigbuf/mgmt_io_in_buf[13] sigbuf/mgmt_io_in_buf[14] sigbuf/mgmt_io_in_buf[15]
+ sigbuf/mgmt_io_in_buf[16] sigbuf/mgmt_io_in_buf[17] sigbuf/mgmt_io_in_buf[18] sigbuf/mgmt_io_in_buf[19]
+ housekeeping/mgmt_gpio_in[3] housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5]
+ housekeeping/mgmt_gpio_in[6] sigbuf/mgmt_io_in_buf[0] sigbuf/mgmt_io_in_buf[1] sigbuf/mgmt_io_in_buf[2]
+ housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_oeb[10] housekeeping/mgmt_gpio_oeb[11]
+ housekeeping/mgmt_gpio_oeb[12] housekeeping/mgmt_gpio_oeb[13] housekeeping/mgmt_gpio_oeb[14]
+ housekeeping/mgmt_gpio_oeb[15] housekeeping/mgmt_gpio_oeb[16] housekeeping/mgmt_gpio_oeb[17]
+ housekeeping/mgmt_gpio_oeb[18] housekeeping/mgmt_gpio_oeb[19] housekeeping/mgmt_gpio_oeb[1]
+ housekeeping/mgmt_gpio_oeb[20] housekeeping/mgmt_gpio_oeb[21] housekeeping/mgmt_gpio_oeb[22]
+ housekeeping/mgmt_gpio_oeb[23] housekeeping/mgmt_gpio_oeb[24] housekeeping/mgmt_gpio_oeb[25]
+ housekeeping/mgmt_gpio_oeb[26] housekeeping/mgmt_gpio_oeb[27] housekeeping/mgmt_gpio_oeb[28]
+ housekeeping/mgmt_gpio_oeb[29] housekeeping/mgmt_gpio_oeb[2] housekeeping/mgmt_gpio_oeb[30]
+ housekeeping/mgmt_gpio_oeb[31] housekeeping/mgmt_gpio_oeb[32] housekeeping/mgmt_gpio_oeb[33]
+ housekeeping/mgmt_gpio_oeb[34] sigbuf/mgmt_io_oeb_unbuf[0] sigbuf/mgmt_io_oeb_unbuf[1]
+ sigbuf/mgmt_io_oeb_unbuf[2] housekeeping/mgmt_gpio_oeb[3] housekeeping/mgmt_gpio_oeb[4]
+ housekeeping/mgmt_gpio_oeb[5] housekeeping/mgmt_gpio_oeb[6] housekeeping/mgmt_gpio_oeb[7]
+ housekeeping/mgmt_gpio_oeb[8] housekeeping/mgmt_gpio_oeb[9] housekeeping/mgmt_gpio_out[0]
+ sigbuf/mgmt_io_out_unbuf[3] sigbuf/mgmt_io_out_unbuf[4] sigbuf/mgmt_io_out_unbuf[5]
+ sigbuf/mgmt_io_out_unbuf[6] housekeeping/mgmt_gpio_out[14] housekeeping/mgmt_gpio_out[15]
+ housekeeping/mgmt_gpio_out[16] housekeeping/mgmt_gpio_out[17] housekeeping/mgmt_gpio_out[18]
+ housekeeping/mgmt_gpio_out[19] housekeeping/mgmt_gpio_out[1] housekeeping/mgmt_gpio_out[20]
+ housekeeping/mgmt_gpio_out[21] housekeeping/mgmt_gpio_out[22] housekeeping/mgmt_gpio_out[23]
+ housekeeping/mgmt_gpio_out[24] sigbuf/mgmt_io_out_unbuf[7] sigbuf/mgmt_io_out_unbuf[8]
+ sigbuf/mgmt_io_out_unbuf[9] sigbuf/mgmt_io_out_unbuf[10] sigbuf/mgmt_io_out_unbuf[11]
+ housekeeping/mgmt_gpio_out[2] sigbuf/mgmt_io_out_unbuf[12] sigbuf/mgmt_io_out_unbuf[13]
+ sigbuf/mgmt_io_out_unbuf[14] sigbuf/mgmt_io_out_unbuf[15] sigbuf/mgmt_io_out_unbuf[16]
+ sigbuf/mgmt_io_out_unbuf[17] sigbuf/mgmt_io_out_unbuf[18] sigbuf/mgmt_io_out_unbuf[19]
+ housekeeping/mgmt_gpio_out[3] housekeeping/mgmt_gpio_out[4] housekeeping/mgmt_gpio_out[5]
+ housekeeping/mgmt_gpio_out[6] sigbuf/mgmt_io_out_unbuf[0] sigbuf/mgmt_io_out_unbuf[1]
+ sigbuf/mgmt_io_out_unbuf[2] housekeeping/pad_flash_clk flash_clkrst_buffers/in_n[7]
+ housekeeping/pad_flash_csb flash_clkrst_buffers/in_n[6] housekeeping/pad_flash_io0_di
+ flash_clkrst_buffers/in_n[1] flash_clkrst_buffers/in_n[3] flash_clkrst_buffers/in_n[5]
+ housekeeping/pad_flash_io1_di flash_clkrst_buffers/in_n[0] flash_clkrst_buffers/in_n[2]
+ flash_clkrst_buffers/in_n[4] clock_ctrl/sel2[0] clock_ctrl/sel2[1] clock_ctrl/sel2[2]
+ clock_ctrl/ext_clk_sel pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3] pll/div[4]
+ pll/enable clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2] pll/ext_trim[0]
+ pll/ext_trim[10] pll/ext_trim[11] pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14]
+ pll/ext_trim[15] pll/ext_trim[16] pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19]
+ pll/ext_trim[1] pll/ext_trim[20] pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23]
+ pll/ext_trim[24] pll/ext_trim[25] pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4]
+ pll/ext_trim[5] pll/ext_trim[6] pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9]
+ por/porb_l housekeeping/pwr_ctrl_out[0] housekeeping/pwr_ctrl_out[1] housekeeping/pwr_ctrl_out[2]
+ housekeeping/pwr_ctrl_out[3] soc/qspi_enabled housekeeping/reset soc/ser_rx soc/ser_tx
+ soc/serial_clock_in housekeeping/serial_data_1 soc/serial_data_2_in soc/serial_load_in
+ soc/serial_resetn_in soc/spi_csb soc/spi_enabled soc/spi_sck soc/spi_sdi soc/spi_sdo
+ soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di soc/flash_io0_do soc/flash_io0_oeb
+ soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb soc/flash_io2_di soc/flash_io2_do
+ soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do soc/flash_io3_oeb soc/trap soc/uart_enabled
+ clock_ctrl/user_clk housekeeping/usr1_vcc_pwrgood housekeeping/usr1_vdd_pwrgood
+ housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood soc/hk_ack_i soc/mprj_adr_o[0]
+ soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14]
+ soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19]
+ soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23]
+ soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28]
+ soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3]
+ soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8]
+ soc/mprj_adr_o[9] clock_ctrl/core_clk soc/hk_cyc_o soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11] soc/hk_dat_i[12] soc/hk_dat_i[13]
+ soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16] soc/hk_dat_i[17] soc/hk_dat_i[18]
+ soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20] soc/hk_dat_i[21] soc/hk_dat_i[22]
+ soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25] soc/hk_dat_i[26] soc/hk_dat_i[27]
+ soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2] soc/hk_dat_i[30] soc/hk_dat_i[31]
+ soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5] soc/hk_dat_i[6] soc/hk_dat_i[7]
+ soc/hk_dat_i[8] soc/hk_dat_i[9] housekeeping/wb_rstn_i soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o soc/mprj_we_o VSUBS housekeeping
Xgpio_control_in_2\[2\] gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[9] padframe/mprj_io_one[2]
+ sigbuf/mgmt_io_out_buf[9] padframe/mprj_io_one[2] padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] gpio_control_in_2\[2\]/resetn
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[2\]/serial_load
+ gpio_control_in_2\[1\]/serial_load mprj/io_in[16] mprj/io_oeb[16] mprj/io_out[16]
+ soc/VPWR mprj/vccd1 gpio_control_in_2\[2\]/zero mprj/vssd1 VSUBS gpio_control_block
Xgpio_defaults_block_30 soc/VPWR gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] VSUBS gpio_defaults_block
Xspare_logic\[0\] spare_logic\[0\]/spare_xfq[0] spare_logic\[0\]/spare_xfq[1] spare_logic\[0\]/spare_xfqn[0]
+ spare_logic\[0\]/spare_xfqn[1] spare_logic\[0\]/spare_xi[0] spare_logic\[0\]/spare_xi[1]
+ spare_logic\[0\]/spare_xi[2] spare_logic\[0\]/spare_xi[3] spare_logic\[0\]/spare_xib
+ spare_logic\[0\]/spare_xmx[0] spare_logic\[0\]/spare_xmx[1] spare_logic\[0\]/spare_xna[0]
+ spare_logic\[0\]/spare_xna[1] spare_logic\[0\]/spare_xno[0] spare_logic\[0\]/spare_xno[1]
+ spare_logic\[0\]/spare_xz[0] spare_logic\[0\]/spare_xz[10] spare_logic\[0\]/spare_xz[11]
+ spare_logic\[0\]/spare_xz[12] spare_logic\[0\]/spare_xz[13] spare_logic\[0\]/spare_xz[14]
+ spare_logic\[0\]/spare_xz[15] spare_logic\[0\]/spare_xz[16] spare_logic\[0\]/spare_xz[17]
+ spare_logic\[0\]/spare_xz[18] spare_logic\[0\]/spare_xz[19] spare_logic\[0\]/spare_xz[1]
+ spare_logic\[0\]/spare_xz[20] spare_logic\[0\]/spare_xz[21] spare_logic\[0\]/spare_xz[22]
+ spare_logic\[0\]/spare_xz[23] spare_logic\[0\]/spare_xz[24] spare_logic\[0\]/spare_xz[25]
+ spare_logic\[0\]/spare_xz[26] spare_logic\[0\]/spare_xz[2] spare_logic\[0\]/spare_xz[3]
+ spare_logic\[0\]/spare_xz[4] spare_logic\[0\]/spare_xz[5] spare_logic\[0\]/spare_xz[6]
+ spare_logic\[0\]/spare_xz[7] spare_logic\[0\]/spare_xz[8] spare_logic\[0\]/spare_xz[9]
+ soc/VPWR VSUBS spare_logic_block
Xflash_clkrst_buffers soc/VPWR flash_clkrst_buffers/in_n[0] housekeeping/wb_rstn_i
+ clock_ctrl/core_clk flash_clkrst_buffers/in_n[1] flash_clkrst_buffers/in_n[2] flash_clkrst_buffers/in_n[3]
+ flash_clkrst_buffers/in_n[4] flash_clkrst_buffers/in_n[5] flash_clkrst_buffers/in_n[6]
+ flash_clkrst_buffers/in_n[7] housekeeping/pad_flash_csb housekeeping/pad_flash_clk
+ padframe/flash_io0_di_core padframe/flash_io1_di_core padframe/clock_core housekeeping/pad_flash_io0_di
+ housekeeping/pad_flash_io1_di pll/osc padframe/flash_io1_do_core soc/resetn_in soc/clk_in
+ padframe/flash_io0_do_core padframe/flash_io1_ieb_core padframe/flash_io0_ieb_core
+ padframe/flash_io1_oeb_core padframe/flash_io0_oeb_core padframe/flash_csb_oeb_core
+ padframe/flash_clk_oeb_core padframe/flash_csb_core padframe/flash_clk_core VSUBS
+ buff_flash_clkrst
Xgpio_defaults_block_10 soc/VPWR gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_defaults_block_31 soc/VPWR gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_in_1a\[5\] gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[0] padframe/mprj_io_one[7] sigbuf/mgmt_io_out_buf[0] padframe/mprj_io_one[7]
+ padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7] padframe/mprj_io_inp_dis[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn gpio_control_in_1a\[5\]/serial_clock
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load mprj/io_in[7]
+ mprj/io_oeb[7] mprj/io_out[7] soc/VPWR mprj/vccd1 gpio_control_in_1a\[5\]/zero mprj/vssd1
+ VSUBS gpio_control_block
Xgpio_defaults_block_32 soc/VPWR gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] VSUBS gpio_defaults_block
Xgpio_control_bidir_2\[2\] gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[19] sigbuf/mgmt_io_oeb_buf[2]
+ sigbuf/mgmt_io_out_buf[19] padframe/mprj_io_one[26] padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] soc/serial_resetn_out
+ gpio_control_bidir_2\[1\]/resetn soc/serial_clock_out gpio_control_bidir_2\[1\]/serial_clock
+ soc/serial_data_2_out gpio_control_bidir_2\[1\]/serial_data_in soc/serial_load_out
+ gpio_control_bidir_2\[1\]/serial_load mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26]
+ soc/VPWR mprj/vccd1 gpio_control_bidir_2\[2\]/zero mprj/vssd1 VSUBS gpio_control_block
.ends

