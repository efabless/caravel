* NGSPICE file created from caravel_openframe.ext - technology: sky130A

.subckt sky130_fd_io__hvsbt_inv_x1 OUT VPWR VGND w_n46_415# a_119_118# SUB
X0 OUT a_119_118# VPWR w_n46_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X1 OUT a_119_118# VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X2 OUT a_119_118# VPWR w_n46_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__hvsbt_xor VPWR VGND IN0 IN1 OUT w_95_503# SUB
X0 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 OUT IN1 a_510_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X4 a_862_167# a_566_375# OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X7 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 VGND a_161_167# a_862_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X10 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 a_566_375# IN1 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X12 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X13 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X14 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 a_510_167# IN0 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X17 VGND IN0 a_161_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__hvsbt_nor IN0 a_239_144# a_295_118# w_0_415# SUB a_66_144# a_66_482#
X0 a_239_144# a_295_118# a_239_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X1 a_239_482# IN0 a_66_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X2 a_66_144# a_295_118# a_239_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.196 pd=1.96 as=0.098 ps=0.98 w=0.7 l=0.6
X3 a_239_144# IN0 a_66_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X4 a_239_144# a_295_118# a_239_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 a_239_482# IN0 a_66_482# w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__hvsbt_inv_x2 VPWR VGND IN OUT w_0_415# SUB
X0 VPWR IN OUT w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X1 OUT IN VPWR w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X2 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X3 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X4 VPWR IN OUT w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 OUT IN VPWR w_0_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_ls_octl OUT_H_N OUT_H IN RST_H SET_H HLD_H_N VPB a_992_934#
+ VCC_IO a_181_1305# a_n17_1379#
X0 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# a_181_1305# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# a_181_1305# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 a_181_1305# IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# a_181_1305# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# a_181_1305# a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# a_181_1305# a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__hvsbt_nand2 IN1 IN0 OUT VGND VPWR w_n42_415# SUB
X0 VPWR IN1 OUT w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X1 OUT IN0 VPWR w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X2 OUT IN1 a_239_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X3 a_239_144# IN0 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X4 VPWR IN1 OUT w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 OUT IN0 VPWR w_n42_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__hvsbt_xorv2 VPWR VGND IN0 IN1 OUT w_95_503# a_566_375# SUB a_742_141#
X0 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 OUT IN1 a_510_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X4 a_862_167# a_742_141# OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X5 VPWR IN1 a_862_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 a_566_375# IN1 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X7 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X8 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X9 VGND a_161_167# a_862_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X10 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 a_566_375# IN1 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X12 a_510_569# IN0 VPWR w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X13 VPWR IN0 a_161_167# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X14 a_862_569# a_161_167# OUT w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X15 OUT a_566_375# a_510_569# w_95_503# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X16 a_510_167# IN0 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X17 VGND IN0 a_161_167# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_octl DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] PUEN_2OR1_H
+ DM_H[1] PDEN_H_N[1] PDEN_H_N[0] SLOW SLOW_H VCC_IO sky130_fd_io__hvsbt_xorv2_0/a_742_141#
+ sky130_fd_io__hvsbt_nand2_0/VPWR sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__hvsbt_inv_x2_3/OUT
+ sky130_fd_io__hvsbt_nor_0/w_0_415# sky130_fd_io__hvsbt_nand2_0/VGND li_n9202_2336#
+ m1_n8913_3102# VPWR sky130_fd_io__hvsbt_nor_0/IN0 sky130_fd_io__hvsbt_nand2_0/IN0
+ sky130_fd_io__hvsbt_xorv2_0/a_566_375# sky130_fd_io__hvsbt_inv_x2_2/OUT sky130_fd_io__hvsbt_nand2_4/IN1
+ SLOW_H_N HLD_I_H_N VGND OD_H
Xsky130_fd_io__hvsbt_inv_x1_4 sky130_fd_io__hvsbt_inv_x2_2/IN VCC_IO VGND VCC_IO li_5323_4140#
+ VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_xor_0 VCC_IO VGND DM_H[2] DM_H[1] sky130_fd_io__hvsbt_xor_0/OUT
+ VCC_IO VGND sky130_fd_io__hvsbt_xor
Xsky130_fd_io__hvsbt_nor_0 sky130_fd_io__hvsbt_nor_0/IN0 sky130_fd_io__hvsbt_nand2_0/IN1
+ li_n9202_2336# sky130_fd_io__hvsbt_nor_0/w_0_415# VGND sky130_fd_io__hvsbt_nand2_0/VGND
+ sky130_fd_io__hvsbt_nand2_0/VPWR sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x2_0 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_0/IN PDEN_H_N[0]
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nor_1 DM_H_N[2] sky130_fd_io__hvsbt_nand2_3/IN0 DM_H_N[1] VCC_IO
+ VGND VGND VCC_IO sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x2_1 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_1/IN PDEN_H_N[1]
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nor_2 sky130_fd_io__hvsbt_nor_2/IN0 li_5323_4140# DM_H_N[1] VCC_IO
+ VGND VGND VCC_IO sky130_fd_io__hvsbt_nor
Xsky130_fd_io__com_ctl_ls_octl_0 SLOW_H_N SLOW_H SLOW OD_H VGND HLD_I_H_N VPWR m2_5755_2254#
+ VCC_IO VPWR VGND sky130_fd_io__com_ctl_ls_octl
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nand2_0/IN0
+ sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__hvsbt_nand2_0/VGND sky130_fd_io__hvsbt_nand2_0/VPWR
+ sky130_fd_io__hvsbt_nor_0/w_0_415# VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__hvsbt_nand2_2/OUT
+ PUEN_2OR1_H VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x2_2 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_2/IN sky130_fd_io__hvsbt_inv_x2_2/OUT
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nand2_2 DM_H[0] sky130_fd_io__hvsbt_xor_0/OUT sky130_fd_io__hvsbt_nand2_2/OUT
+ VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x2_3 VCC_IO VGND sky130_fd_io__hvsbt_inv_x2_3/IN sky130_fd_io__hvsbt_inv_x2_3/OUT
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_nand2_3 DM_H_N[0] sky130_fd_io__hvsbt_nand2_3/IN0 sky130_fd_io__hvsbt_nand2_3/OUT
+ VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_4 sky130_fd_io__hvsbt_nand2_4/IN1 PUEN_2OR1_H sky130_fd_io__hvsbt_nand2_4/OUT
+ VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_5 DM_H_N[1] DM_H_N[2] sky130_fd_io__hvsbt_nand2_6/IN1 VGND
+ VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_6 sky130_fd_io__hvsbt_nand2_6/IN1 DM_H_N[0] sky130_fd_io__hvsbt_nand2_6/OUT
+ VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_7 DM_H[0] DM_H[1] sky130_fd_io__hvsbt_nand2_7/OUT VGND
+ VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_xorv2_0 VCC_IO VGND DM_H[2] DM_H[0] sky130_fd_io__hvsbt_nor_2/IN0
+ VCC_IO sky130_fd_io__hvsbt_xorv2_0/a_566_375# VGND sky130_fd_io__hvsbt_xorv2_0/a_742_141#
+ sky130_fd_io__hvsbt_xorv2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x2_0/IN VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2_7/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x2_3/IN VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_inv_x1_3/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 sky130_fd_io__hvsbt_inv_x2_1/IN VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2_6/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_3 sky130_fd_io__hvsbt_inv_x1_3/OUT VCC_IO VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2_4/OUT VGND sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__gpio_dat_ls_1v2 IN OUT_H_N RST_H SET_H HLD_H_N OUT_H VPWR_KA
+ VGND VCC_IO
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X24 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X31 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X32 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X37 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X39 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X40 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__gpio_dat_lsv2 IN OUT_H_N RST_H SET_H HLD_H_N OUT_H VPWR_KA a_28_14#
+ VGND VCC_IO
X0 a_2251_36# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1 a_28_633# SET_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 a_1720_1202# HLD_H_N a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.5
X3 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X4 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X5 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X8 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X9 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X10 VPWR_KA a_2251_2228# a_2251_36# VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X12 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X13 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_28_633# a_28_14# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND IN a_2251_2228# VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 OUT_H a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X17 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X18 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X19 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X20 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X21 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X22 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X23 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X24 VGND a_28_633# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X25 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X26 a_2251_2228# IN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X28 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X29 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X30 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X31 a_2251_2228# IN VPWR_KA VPWR_KA sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X32 VGND a_28_633# a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X33 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X34 a_1484_128# VPWR_KA a_1251_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X35 VGND a_2251_36# a_1484_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X36 VGND a_2251_2228# a_2251_36# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X37 a_28_633# a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X38 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X39 a_28_14# a_28_633# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X40 a_1251_128# VPWR_KA a_1484_128# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X41 a_1251_128# HLD_H_N a_28_633# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X42 VCC_IO a_28_14# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_1484_128# a_2251_36# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X44 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X45 a_2080_128# VPWR_KA a_1720_1202# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X46 VGND RST_H a_28_14# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X47 OUT_H_N a_28_14# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X48 a_2080_128# a_2251_2228# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X49 VGND a_2251_2228# a_2080_128# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_io__com_cclat PU_DIS_H PD_DIS_H OE_H_N DRVLO_H_N DRVHI_H VGND VCC_IO
X0 a_947_1193# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X1 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X2 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X3 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 VGND DRVHI_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X6 VCC_IO PU_DIS_H a_638_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X10 a_2361_1095# DRVHI_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X11 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X15 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VGND PU_DIS_H a_638_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X17 a_4762_1193# DRVHI_H a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X18 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X19 VGND PD_DIS_H a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X20 a_505_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X21 VCC_IO a_638_279# a_947_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X22 a_3417_1193# DRVHI_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X23 a_2361_1095# PD_DIS_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X24 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X25 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X26 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X27 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X28 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X30 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 VCC_IO OE_H_N a_176_279# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X32 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X33 a_2361_1095# PD_DIS_H a_4762_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_987_279# DRVLO_H_N a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X35 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X36 DRVHI_H a_947_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X37 a_947_1193# a_176_279# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 VGND OE_H_N a_176_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X39 VCC_IO a_947_1193# DRVHI_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 VCC_IO a_2361_1095# DRVLO_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X41 DRVLO_H_N a_2361_1095# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X42 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X43 DRVHI_H a_947_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X44 VCC_IO a_505_1193# a_3417_1193# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X45 a_4762_1193# PD_DIS_H a_2361_1095# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X46 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X47 VGND a_947_1193# DRVHI_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X48 a_947_1193# a_638_279# a_1628_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X49 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X50 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X51 a_1628_279# DRVLO_H_N a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X52 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X53 a_505_1193# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X54 DRVLO_H_N a_2361_1095# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X55 VGND a_505_1193# a_2361_1095# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X56 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X57 VGND a_176_279# a_987_279# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X58 a_3417_1193# a_505_1193# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X59 VGND a_2361_1095# DRVLO_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X60 a_2361_1095# a_505_1193# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X61 a_987_279# a_176_279# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X62 a_1628_279# a_638_279# a_947_1193# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_opath_datoev2 DRVLO_H_N VCC_IO HLD_I_OVR_H OE_H a_5565_99#
+ OUT OE_N sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA DRVHI_H li_5565_99# sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ VGND OD_H
Xsky130_fd_io__gpio_dat_ls_1v2_0 OUT sky130_fd_io__com_cclat_0/PU_DIS_H VGND sky130_fd_io__gpio_dat_ls_1v2_0/SET_H
+ HLD_I_OVR_H sky130_fd_io__com_cclat_0/PD_DIS_H VPWR_KA VGND VCC_IO sky130_fd_io__gpio_dat_ls_1v2
Xsky130_fd_io__gpio_dat_lsv2_0 OE_N OE_H VGND OD_H HLD_I_OVR_H sky130_fd_io__com_cclat_0/OE_H_N
+ VPWR_KA a_28_1762# VGND VCC_IO sky130_fd_io__gpio_dat_lsv2
Xsky130_fd_io__com_cclat_0 sky130_fd_io__com_cclat_0/PU_DIS_H sky130_fd_io__com_cclat_0/PD_DIS_H
+ sky130_fd_io__com_cclat_0/OE_H_N DRVLO_H_N DRVHI_H VGND VCC_IO sky130_fd_io__com_cclat
.ends

.subckt sky130_fd_io__com_pdpredrvr_strong_slowv2 DRVLO_H_N PDEN_H_N VCC_IO VGND_IO
+ PD_H w_59_800#
X0 VCC_IO PDEN_H_N a_125_866# w_59_800# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 PD_H DRVLO_H_N VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 VGND_IO PDEN_H_N PD_H SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X3 a_125_866# DRVLO_H_N PD_H w_59_800# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X4 a_125_866# PDEN_H_N VCC_IO w_59_800# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X5 PD_H DRVLO_H_N a_125_866# w_59_800# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__com_pdpredrvr_weakv2 DRVLO_H_N PDEN_H_N PD_H VGND_IO VCC_IO
X0 PD_H DRVLO_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X1 a_73_866# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X2 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X3 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X4 VCC_IO PDEN_H_N a_73_866# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
.ends

.subckt sky130_fd_io__com_pdpredrvr_pbiasv2 EN_H VGND_IO PBIAS DRVLO_H_N EN_H_N PDEN_H_N
+ PD_H a_16899_3078# a_12434_3172# a_12120_4573# a_13911_2980# SUB a_18190_3078# VCC_IO
+ a_16799_2980#
X0 VGND_IO a_11581_4213# a_12120_4573# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
R0 m1_16797_3553# a_16899_3078# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X1 VCC_IO a_16799_2980# a_16899_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X2 VCC_IO a_13347_3873# a_16799_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X3 PBIAS PBIAS a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 VCC_IO a_16799_2980# a_16899_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 a_16899_3078# a_16799_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R1 m1_12556_4086# a_11581_4213# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X6 a_11781_4311# a_11581_4213# VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=1
X7 VCC_IO a_13911_2980# a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X8 a_11460_4784# a_11368_4652# a_11368_4652# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X9 a_11460_4784# DRVLO_H_N VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 PBIAS PBIAS a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X11 a_16899_3078# a_16799_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_18190_3078# a_12120_4573# a_12120_4573# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 a_16799_2980# a_18190_3078# a_18190_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 PBIAS PBIAS a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X15 a_13911_2980# PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R2 a_11368_4652# m1_13251_3471# sky130_fd_pr__res_generic_m1 w=0.64 l=10m
R3 m1_13288_3471# EN_H_N sky130_fd_pr__res_generic_m1 w=0.64 l=10m
R4 a_12578_4025# m1_12556_4086# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X16 a_13911_2980# a_13911_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X17 VGND_IO a_11460_4784# a_11581_4213# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X18 VGND_IO a_11581_4213# a_11781_4311# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X19 VCC_IO a_16799_2980# a_16899_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X20 a_16799_2980# a_18190_3078# a_18190_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R5 m1_11681_3387# PD_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R6 a_13911_2980# m1_15141_3027# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X21 a_13911_2980# a_13911_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X22 VCC_IO a_13911_2980# a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X23 a_13911_2980# PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X24 a_16899_3078# a_16799_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X25 VGND_IO PD_H a_12434_3172# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X26 a_18190_3078# a_18190_3078# a_16799_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
R7 PBIAS m1_12872_3935# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R8 m1_15178_3027# PBIAS sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X27 PBIAS a_11581_4213# VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X28 a_11581_4213# DRVLO_H_N VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X29 VCC_IO DRVLO_H_N a_13347_3873# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X30 a_12120_4573# a_12120_4573# a_18190_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X31 a_13219_3078# DRVLO_H_N a_11581_4213# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.795 ps=6.53 w=3 l=0.5
R9 a_11781_4311# m1_11840_4382# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 m1_12872_3935# a_12906_4025# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X32 VGND_IO PDEN_H_N a_11460_4784# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
R11 a_11368_4652# m1_11681_3387# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_12906_4025# a_11581_4213# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X34 VCC_IO EN_H_N a_13361_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.315 ps=3.21 w=3 l=0.5
X35 a_13911_2980# a_13911_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X36 PBIAS PBIAS a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X37 a_13911_2980# PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X38 a_16899_3078# a_16799_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X39 a_18190_3078# a_12120_4573# a_12120_4573# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 VGND_IO a_11581_4213# PBIAS SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=1
X41 VCC_IO a_13911_2980# a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X42 a_13347_3873# DRVLO_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X43 a_16799_2980# VGND_IO VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=8
R12 a_11460_4784# m1_11524_4738# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
X44 a_13347_3873# DRVLO_H_N VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X45 a_13361_3078# a_11368_4652# a_13219_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.315 pd=3.21 as=0.315 ps=3.21 w=3 l=0.5
X46 PBIAS a_13347_3873# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
R13 m1_11840_4382# PBIAS sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X47 VCC_IO EN_H PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X48 a_13911_2980# a_13911_2980# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X49 VCC_IO a_13911_2980# a_13911_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X50 a_12120_4573# a_12120_4573# a_18190_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X51 a_18190_3078# a_18190_3078# a_16799_2980# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X52 VGND_IO EN_H_N a_11581_4213# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X53 a_13911_2980# PBIAS PBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X54 VCC_IO a_16799_2980# a_16899_3078# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X55 a_12578_4025# PD_H a_12434_3172# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
R14 a_11368_4652# m1_11524_4701# sky130_fd_pr__res_generic_m1 w=2.5 l=10m
R15 a_13911_2980# m1_16797_3553# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
.ends

.subckt sky130_fd_io__gpiov2_octl_mux SEL_H_N A_H Y_H B_H SEL_H a_1266_1185# w_1191_2415#
X0 Y_H SEL_H A_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X1 A_H SEL_H_N Y_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X2 Y_H SEL_H B_H w_1191_2415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 B_H SEL_H_N Y_H a_1266_1185# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 DRVLO_H_N PD_I2C_H PDEN_H_N PD_H
+ VCC_IO I2C_MODE_H EN_FAST_N[0] EN_FAST_N[1] VGND_IO w_4658_n980#
X0 a_5469_n914# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X1 PD_H I2C_MODE_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 VCC_IO I2C_MODE_H a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X3 PD_I2C_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X4 a_4877_n914# I2C_MODE_H VCC_IO w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X5 PD_H DRVLO_H_N a_5781_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X6 PD_I2C_H DRVLO_H_N a_6596_n885# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X7 VCC_IO PDEN_H_N a_6596_n885# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X8 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X9 a_4877_n914# I2C_MODE_H VCC_IO w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X10 PD_I2C_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X11 a_5781_n914# EN_FAST_N[1] a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X12 a_7449_n1327# PDEN_H_N a_4877_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X13 a_4877_n914# EN_FAST_N[0] a_5469_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X14 a_7449_n1327# PDEN_H_N a_6596_n1327# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X15 a_6596_n1327# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X16 VGND_IO DRVLO_H_N PD_I2C_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X17 VCC_IO EN_FAST_N[1] a_7724_n1285# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=1
X18 VGND_IO PDEN_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X19 a_5781_n914# DRVLO_H_N PD_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X20 a_7724_n1285# DRVLO_H_N PD_I2C_H w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X21 PD_H DRVLO_H_N a_5469_n914# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X22 PD_I2C_H DRVLO_H_N a_7724_n1285# w_4658_n980# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X23 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 EN_FAST_N[0] EN_FAST_N[1] I2C_MODE_H
+ PDEN_H_N DRVLO_H_N PD_H VGND_IO VCC_IO
X0 a_1992_n250# PDEN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X1 VCC_IO EN_FAST_N[0] a_2168_n356# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X2 a_1139_172# I2C_MODE_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X3 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X4 a_2168_n356# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X5 a_1139_172# EN_FAST_N[1] a_1708_456# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X6 a_1992_n250# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=2
X7 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X8 VCC_IO I2C_MODE_H a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X9 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_1708_456# DRVLO_H_N PD_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.5
X11 PD_H DRVLO_H_N a_2477_n356# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X12 PD_H PDEN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X13 PD_H DRVLO_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X14 a_1708_456# EN_FAST_N[0] a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
X15 VGND_IO DRVLO_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X16 PD_H DRVLO_H_N a_1708_456# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
X17 PD_H DRVLO_H_N a_1592_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=2
X18 a_2477_n356# EN_FAST_N[1] VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X19 a_1592_172# PDEN_H_N a_1139_172# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=2
X20 VGND_IO PDEN_H_N PD_H VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_pdpredrvr_strong PD_H[3] PD_H[2] DRVLO_H_N PDEN_H_N I2C_MODE_H_N
+ PD_H[4] sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078# sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980# SLOW_H sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ m2_9346_3287# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172# sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ VCC_IO VGND
Xsky130_fd_io__com_pdpredrvr_pbiasv2_0 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H
+ VGND sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS DRVLO_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N
+ PDEN_H_N PD_H[4] sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573# sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ VGND sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078# VCC_IO sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__com_pdpredrvr_pbiasv2
Xsky130_fd_io__gpiov2_octl_mux_0 I2C_MODE_H_N sky130_fd_io__gpiov2_octl_mux_0/A_H
+ sky130_fd_io__gpiov2_octl_mux_0/Y_H DRVLO_H_N sky130_fd_io__hvsbt_nand2_1/IN0 VGND
+ VCC_IO sky130_fd_io__gpiov2_octl_mux
Xsky130_fd_io__hvsbt_nand2_0 SLOW_H I2C_MODE_H_N sky130_fd_io__hvsbt_nand2_0/OUT VGND
+ VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 SLOW_H sky130_fd_io__hvsbt_nand2_1/IN0 sky130_fd_io__hvsbt_nand2_1/OUT
+ VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_nr2_0 DRVLO_H_N PD_H[4] PDEN_H_N PD_H[2] VCC_IO
+ sky130_fd_io__hvsbt_inv_x1_1/OUT sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ VGND VCC_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VCC_IO VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2_0/OUT VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0]
+ sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] sky130_fd_io__hvsbt_inv_x1_1/OUT
+ PDEN_H_N sky130_fd_io__gpiov2_octl_mux_0/Y_H PD_H[3] VGND VCC_IO sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x1_1/OUT VCC_IO VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2_1/OUT VGND sky130_fd_io__hvsbt_inv_x1
R0 m1_9403_1623# m1_9430_1596# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0] m1_9575_2734# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R2 m1_9427_1780# sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
R3 m1_9575_2734# VCC_IO sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R4 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] m1_9830_1715# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[0] m1_9830_1752# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X1 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X2 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.21 ps=1.42 w=1 l=0.6
R6 sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS m1_9364_1624# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X3 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H PDEN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.335 ps=2.67 w=1 l=0.6
R7 m1_9364_1624# m1_9403_1623# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X4 VCC_IO sky130_fd_io__hvsbt_inv_x1_0/OUT a_8987_763# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.63 pd=3.42 as=0.42 ps=3.28 w=3 l=0.6
R8 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N m1_9562_1482# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X5 a_8987_763# PDEN_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=1 ps=6.67 w=3 l=0.6
R9 m1_9599_1482# sky130_fd_io__gpiov2_pdpredrvr_strong_nr3_0/EN_FAST_N[1] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X6 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.63 ps=3.42 w=3 l=0.6
X7 sky130_fd_io__hvsbt_nand2_1/IN0 I2C_MODE_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.6
X8 VGND PD_H[4] sky130_fd_io__gpiov2_octl_mux_0/A_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.5
R10 sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS m1_9427_1780# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X9 VGND sky130_fd_io__hvsbt_inv_x1_0/OUT sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.42 as=0.14 ps=1.28 w=1 l=0.6
R11 sky130_fd_io__com_pdpredrvr_pbiasv2_0/EN_H_N m1_9430_1559# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X10 VCC_IO PD_H[4] sky130_fd_io__gpiov2_octl_mux_0/A_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__com_pupredrvr_strong_slowv2 PUEN_H DRVHI_H PU_H_N VGND_IO a_93_102#
+ VCC_IO
X0 PU_H_N DRVHI_H a_93_102# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X1 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X2 a_93_102# PUEN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X3 VCC_IO PUEN_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X4 a_93_102# DRVHI_H PU_H_N VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X5 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X6 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X7 VGND_IO PUEN_H a_93_102# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
.ends

.subckt sky130_fd_io__feas_com_pupredrvr_weak DRVHI_H PUEN_H PU_H_N VGND_IO VCC_IO
+ w_21_799#
X0 VCC_IO DRVHI_H PU_H_N w_21_799# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X1 PU_H_N DRVHI_H VCC_IO w_21_799# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X2 a_280_102# PUEN_H VGND_IO SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X3 PU_H_N DRVHI_H a_280_102# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X4 VCC_IO PUEN_H PU_H_N w_21_799# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__feascom_pupredrvr_nbiasv2 EN_H_N EN_H NBIAS DRVHI_H PUEN_H PU_H_N
+ a_261_220# VGND_IO a_2821_220# a_2874_118# VCC_IO a_1772_220#
X0 VCC_IO DRVHI_H a_207_1014# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.192 pd=1.38 as=0.14 ps=1.28 w=1 l=0.5
X1 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X2 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X3 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X4 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X5 a_1672_194# a_207_1014# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X6 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.192 ps=1.38 w=1 l=0.8
X7 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X8 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R0 a_562_1898# m1_2838_1831# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 NBIAS m1_1014_127# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X9 VCC_IO a_250_1898# a_2874_118# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X10 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
R2 NBIAS m1_1014_800# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X11 VGND_IO a_1672_194# a_1772_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R3 EN_H m1_575_1252# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X12 VCC_IO DRVHI_H a_562_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.51 as=0.14 ps=1.28 w=1 l=0.5
X13 a_261_220# a_261_220# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R4 a_620_1263# m1_2838_1794# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 m1_612_1252# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X14 a_250_1898# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X15 VGND_IO DRVHI_H a_207_1014# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.324 pd=2.02 as=0.265 ps=2.53 w=1 l=0.6
X16 VGND_IO a_207_1014# NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X17 VGND_IO a_250_1898# a_1004_990# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=4
X18 NBIAS NBIAS a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R6 NBIAS m1_1409_1332# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X19 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X20 a_2874_118# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.04 ps=5.51 w=5 l=0.5
X21 a_583_914# EN_H VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.77 as=0.324 ps=2.02 w=1.5 l=0.5
X22 a_2821_220# a_2874_118# a_2874_118# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R7 m1_1608_646# a_1772_220# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X23 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X24 NBIAS a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X25 a_207_1014# DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X26 a_250_1898# a_562_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R8 a_2421_2014# m1_2596_1928# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X27 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X28 NBIAS EN_H_N VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X29 VCC_IO a_250_1898# a_1507_1397# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X30 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.04 pd=5.51 as=0.42 ps=3.28 w=3 l=0.5
X31 a_1772_220# a_1672_194# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X32 a_2821_220# a_2821_220# a_1672_194# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
R9 m1_2596_1928# a_250_1898# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 PU_H_N m1_702_1715# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R11 m1_1409_1332# a_1507_1397# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X33 a_1507_1397# a_250_1898# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
R12 m1_1046_126# a_261_220# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X34 VCC_IO EN_H a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X35 a_562_1898# PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X36 a_2421_2014# PU_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.185 ps=1.51 w=0.42 l=8
X37 a_737_914# a_620_1263# a_583_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.77 as=0.203 ps=1.77 w=1.5 l=0.5
R13 m1_702_1715# a_620_1263# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R14 m1_1014_800# a_1004_990# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X38 VCC_IO a_250_1898# NBIAS VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X39 a_261_220# NBIAS NBIAS VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X40 VGND_IO a_261_220# a_261_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
R15 a_261_220# m1_1608_646# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
X41 VCC_IO a_562_1898# a_250_1898# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X42 a_250_1898# DRVHI_H a_737_914# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.203 ps=1.77 w=1.5 l=0.5
X43 a_1672_194# a_2821_220# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X44 a_562_1898# a_620_1263# a_620_1263# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X45 a_1672_194# VCC_IO VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=8
X46 a_2874_118# a_2874_118# a_2821_220# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2 DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] PU_H_N VGND_IO a_158_632# VCC_IO
R0 m1_1184_866# PU_H_N sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X2 VGND_IO EN_FAST[3] a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
R1 a_158_632# m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X3 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X4 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X5 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
R2 PU_H_N a_1008_2434# sky130_fd_pr__res_generic_po w=0.33 l=4
X6 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
R3 a_158_632# a_1008_2434# sky130_fd_pr__res_generic_po w=0.33 l=11
X7 a_809_632# EN_FAST[2] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X8 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X9 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X10 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X11 PU_H_N DRVHI_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X12 VGND_IO PUEN_H a_158_109# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X13 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a DRVHI_H PUEN_H EN_FAST[0] EN_FAST[1]
+ EN_FAST[2] EN_FAST[3] PU_H_N VGND_IO a_353_606# a_609_606# VCC_IO
R0 m1_1184_866# PU_H_N sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X0 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.6
X1 a_311_632# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X2 VGND_IO a_353_606# a_311_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X3 VGND_IO PUEN_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
R1 a_158_632# m1_1184_866# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X4 PU_H_N DRVHI_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
X5 PU_H_N PUEN_H VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.6
X6 VCC_IO DRVHI_H PU_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.6
R2 PU_H_N a_1008_2434# sky130_fd_pr__res_generic_po w=0.33 l=4
X7 a_158_632# DRVHI_H a_809_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
R3 a_158_632# a_1008_2434# sky130_fd_pr__res_generic_po w=0.33 l=11
X8 a_809_632# a_609_606# VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
X9 a_158_632# DRVHI_H a_809_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.165 ps=1.72 w=1.5 l=0.5
X10 a_311_1060# DRVHI_H a_158_632# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.71 as=0.398 ps=3.53 w=1.5 l=0.5
X11 VGND_IO EN_FAST[0] a_311_1060# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.157 ps=1.71 w=1.5 l=1
X12 PU_H_N DRVHI_H a_158_199# VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=4
X13 a_809_1060# EN_FAST[1] VGND_IO VGND_IO sky130_fd_pr__nfet_g5v0d10v5 ad=0.165 pd=1.72 as=0.21 ps=1.78 w=1.5 l=1
.ends

.subckt sky130_fd_io__gpio_pupredrvr_strongv2 VCC_IO PU_H_N[3] PU_H_N[2] SLOW_H_N
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS SUB sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220# PUEN_H DRVHI_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
Xsky130_fd_io__feascom_pupredrvr_nbiasv2_0 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ DRVHI_H PUEN_H PU_H_N[2] sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220# SUB
+ sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220# sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ VCC_IO sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220# sky130_fd_io__feascom_pupredrvr_nbiasv2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] PU_H_N[3] SUB sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ VCC_IO sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xsky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0 DRVHI_H PUEN_H sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] PU_H_N[2] SUB sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3]
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] VCC_IO sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a
R0 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] m1_6556_1365# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R1 SUB m1_6555_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X0 VCC_IO PUEN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
R2 m1_6299_1273# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R3 SUB m1_6266_605# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R4 m1_5759_509# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X1 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SLOW_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
R5 m1_4777_1326# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R6 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS m1_5786_421# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 m1_4655_1468# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_a_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] m1_6266_568# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R9 m1_5786_421# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6300_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X2 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
R11 m1_6265_477# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[2] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R12 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H m1_5722_509# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R13 SUB m1_6299_1273# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R14 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[1] m1_6300_1365# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R15 m1_6555_1273# sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[0] sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6265_477# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X3 SUB PUEN_H a_483_1179# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 a_483_1179# SLOW_H_N sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H_N SUB SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
R17 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/EN_H m1_4740_1326# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R18 sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/EN_FAST[3] m1_6556_1402# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R19 sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS m1_4655_1468# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
.ends

.subckt sky130_fd_io__gpiov2_obpredrvr PD_H[3] PD_H[2] DRVLO_H_N PU_H_N[3] PU_H_N[2]
+ PU_H_N[1] PU_H_N[0] PD_H[0] PD_H[4] PUEN_H[1] PUEN_H[0] PDEN_H_N[0] SLOW_H_N I2C_MODE_H_N
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ SLOW_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ DRVHI_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102# sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ PD_H[1] SUB sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ PDEN_H_N[1] VCC_IO
Xsky130_fd_io__com_pdpredrvr_strong_slowv2_0 DRVLO_H_N PDEN_H_N[1] VCC_IO SUB PD_H[1]
+ VCC_IO sky130_fd_io__com_pdpredrvr_strong_slowv2
Xsky130_fd_io__com_pdpredrvr_weakv2_0 DRVLO_H_N PDEN_H_N[0] PD_H[0] SUB VCC_IO sky130_fd_io__com_pdpredrvr_weakv2
Xsky130_fd_io__gpiov2_pdpredrvr_strong_0 PD_H[3] PD_H[2] DRVLO_H_N PDEN_H_N[1] I2C_MODE_H_N
+ PD_H[4] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ SLOW_H sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ PUEN_H[1] sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H VCC_IO
+ SUB sky130_fd_io__gpiov2_pdpredrvr_strong
Xsky130_fd_io__com_pupredrvr_strong_slowv2_0 PUEN_H[1] DRVHI_H PU_H_N[1] SUB sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ VCC_IO sky130_fd_io__com_pupredrvr_strong_slowv2
Xsky130_fd_io__feas_com_pupredrvr_weak_0 DRVHI_H PUEN_H[0] PU_H_N[0] SUB VCC_IO VCC_IO
+ sky130_fd_io__feas_com_pupredrvr_weak
Xsky130_fd_io__gpio_pupredrvr_strongv2_0 VCC_IO PU_H_N[3] PU_H_N[2] SLOW_H_N sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ SUB sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ PUEN_H[1] DRVHI_H sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpio_pupredrvr_strongv2
.ends

.subckt sky130_fd_io__gpiov2_octl_dat VPWR_KA SLOW HLD_I_OVR_H OD_H SLOW_H_N DRVHI_H
+ PU_H_N[2] PU_H_N[1] PU_H_N[0] PD_H[1] PD_H[0] PD_H[4] DRVLO_H_N PD_H[3] PD_H[2]
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] DM_H[1] DM_H_N[0] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ DM_H_N[1] DM_H_N[2] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N sky130_fd_io__com_opath_datoev2_0/li_5565_99# sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N DM_H[2] sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ VPWR sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ PU_H_N[3] SUB
Xsky130_fd_io__gpiov2_octl_0 DM_H[0] DM_H[2] DM_H_N[0] DM_H_N[1] DM_H_N[2] sky130_fd_io__gpiov2_octl_0/PUEN_2OR1_H
+ DM_H[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0]
+ SLOW sky130_fd_io__gpiov2_octl_0/SLOW_H VCC_IO a_13335_4479# VCC_IO sky130_fd_io__gpiov2_obpredrvr_0/I2C_MODE_H_N
+ sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[1] VCC_IO SUB DM_H[0] VCC_IO VPWR DM_H[1]
+ DM_H[2] a_13335_4479# sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[0] VCC_IO SLOW_H_N
+ HLD_I_H_N SUB OD_H sky130_fd_io__gpiov2_octl
Xsky130_fd_io__com_opath_datoev2_0 DRVLO_H_N VCC_IO HLD_I_OVR_H sky130_fd_io__com_opath_datoev2_0/OE_H
+ SUB OUT OE_N sky130_fd_io__com_opath_datoev2_0/sky130_fd_io__com_cclat_0/PD_DIS_H
+ VPWR_KA DRVHI_H sky130_fd_io__com_opath_datoev2_0/li_5565_99# OD_H SUB OD_H sky130_fd_io__com_opath_datoev2
Xsky130_fd_io__gpiov2_obpredrvr_0 PD_H[3] PD_H[2] DRVLO_H_N PU_H_N[3] PU_H_N[2] PU_H_N[1]
+ PU_H_N[0] PD_H[0] PD_H[4] sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[1] sky130_fd_io__gpiov2_obpredrvr_0/PUEN_H[0]
+ sky130_fd_io__gpiov2_octl_0/PDEN_H_N[0] SLOW_H_N sky130_fd_io__gpiov2_obpredrvr_0/I2C_MODE_H_N
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_octl_0/SLOW_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ DRVHI_H sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ PD_H[1] SUB sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_octl_0/PDEN_H_N[1] VCC_IO sky130_fd_io__gpiov2_obpredrvr
.ends

.subckt sky130_fd_io__com_pudrvr_strong_slowv2 PU_H_N PAD w_122_n30# a_356_297#
X0 a_356_297# PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X1 PAD PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_122_n30# PU_H_N a_356_297# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X3 PAD PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_122_n30# PU_H_N a_356_297# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X5 w_122_n30# PU_H_N PAD w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X6 w_122_n30# PU_H_N PAD w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X7 a_356_297# PU_H_N w_122_n30# w_122_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
.ends

.subckt sky130_fd_io__com_res_weak_bentbigres a_419_6804# a_419_8054# a_n256_8772#
+ a_419_8146# a_n258_6046# a_419_9396# a_n2_6046#
R0 a_n258_6046# a_n256_8772# sky130_fd_pr__res_generic_po w=0.8 l=12
R1 a_419_8146# a_419_9396# sky130_fd_pr__res_generic_po w=0.8 l=6
R2 a_n258_6046# a_n2_6046# sky130_fd_pr__res_generic_po w=0.8 l=50
R3 a_419_6804# a_419_8054# sky130_fd_pr__res_generic_po w=0.8 l=6
.ends

.subckt sky130_fd_io__com_res_weak RB RA sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ li_n135_8054# a_n160_10423# li_n135_6820# a_n160_9488#
Xsky130_fd_io__com_res_weak_bentbigres_0 li_n135_6820# li_n135_8054# li_n135_6820#
+ li_n135_8054# sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046# a_n160_9488#
+ RA sky130_fd_io__com_res_weak_bentbigres
R0 a_n160_9838# a_n160_10423# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R1 a_n160_9488# a_n160_9838# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R2 m1_n147_10115# a_n160_10423# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 m1_n147_8777# a_n160_9488# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R4 m1_532_10115# a_n160_10423# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R5 m1_532_9534# a_517_9818# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R6 li_n135_8054# m1_n147_8777# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R7 a_n160_9838# m1_n147_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R8 a_517_9818# m1_532_10115# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R9 RB a_517_9818# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R10 RB m1_532_9534# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R11 m1_n147_9555# a_n160_9838# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R12 li_n135_8054# m1_n146_7735# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R13 a_517_9818# a_n160_10423# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R14 a_n160_9488# m1_n147_9555# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R15 li_n135_6820# m1_n146_7434# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270v2 w_415_600# a_2303_1380# a_13777_1380#
+ a_8817_1380# a_4287_1380# a_7263_1380# a_12223_1380# a_9247_1380# a_2865_1380# a_5841_1380#
+ a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380# a_12785_1380# a_7825_1380#
+ a_3295_1380# a_9809_1380# a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380#
+ a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_11793_1380# a_881_1380# a_6833_1380#
X0 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X1 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X3 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X4 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X7 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X8 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X10 a_1001_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X11 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X12 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X13 w_415_600# a_10239_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_1001_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 w_415_600# a_3295_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X16 w_415_600# a_2303_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_415_600# a_7263_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_1001_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X19 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X20 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X21 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X22 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X23 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_1001_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X26 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X27 a_1001_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X30 w_415_600# a_13215_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X31 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X32 w_415_600# a_6271_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X34 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X35 w_415_600# a_5279_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X36 a_1001_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X37 a_1001_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_415_600# a_9247_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X42 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X43 a_1001_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X44 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X45 a_1001_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X46 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 w_415_600# a_12223_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X48 a_1001_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X49 a_1001_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X50 a_1001_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X51 w_415_600# a_4287_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X52 w_415_600# a_14135_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X53 w_415_600# a_8255_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 a_1001_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X55 w_415_600# a_11231_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strongv2 PU_H_N[3] PU_H_N[2] VCC_IO TIE_HI_ESD m1_1330_n459#
+ m1_6027_281# m1_3418_50# VNB a_14575_n157# m1_6652_281# m1_3028_333# PAD m1_14880_n614#
+ li_9083_n155#
Xsky130_fd_io__pfet_con_diff_wo_abt_270v2_0 VCC_IO PU_H_N[2] m1_14229_1478# m1_8837_1478#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_8837_1478# PU_H_N[2] PU_H_N[3] PU_H_N[3] m1_10391_1478#
+ m1_14229_1478# PU_H_N[2] PU_H_N[2] PU_H_N[3] PU_H_N[2] m1_10391_1478# PAD PU_H_N[3]
+ PU_H_N[3] m1_11745_1478# m1_10391_1478# m1_8837_1478# PU_H_N[2] m1_13667_1478# PU_H_N[3]
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270v2
R0 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 PU_H_N[2] m2_12849_n185# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_10673_n208# m1_8837_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 PU_H_N[2] m2_11422_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 PU_H_N[2] m2_10673_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 TIE_HI_ESD m2_10197_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_11745_1478# m2_12608_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 TIE_HI_ESD m2_10945_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_11745_1478# m2_12849_116# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 PU_H_N[3] m2_12608_n185# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 PU_H_N[2] m2_14769_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 PU_H_N[3] m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 PU_H_N[3] m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 TIE_HI_ESD a_14575_n157# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R18 TIE_HI_ESD m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_8837_1478# m2_10197_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8837_1478# m2_10439_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 PU_H_N[3] m2_14532_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m2_11186_n208# m1_10391_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 TIE_HI_ESD m2_13593_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m2_13837_658# m1_13667_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 m2_12365_n184# m1_11745_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 PU_H_N[3] m2_10439_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 TIE_HI_ESD m2_12365_n184# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m2_14286_658# m1_14229_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 PU_H_N[2] m2_14075_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270v2 VCC_IO PAD a_10282_1285# a_5322_1285#
+ a_12266_1285# a_7306_1285# VSSIO a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285#
+ a_10844_1285# a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285#
+ a_4330_1285# a_3338_1285# a_11274_1285# a_6314_1285# a_8298_1285# a_13258_1285#
+ a_9290_1285# a_1916_1285# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285#
X0 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X1 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X3 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X4 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X7 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X8 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X10 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X11 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X12 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X13 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X16 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X19 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X20 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X21 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X22 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X23 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X26 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X27 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 VSSIO a_11274_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 VSSIO a_5322_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X30 PAD a_9852_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X31 PAD a_10844_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X32 VSSIO a_2346_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 PAD a_6876_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X34 VSSIO a_6314_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X35 PAD a_1916_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X36 VSSIO a_12266_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X37 PAD a_11836_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 PAD a_4892_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 VSSIO a_4330_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 VSSIO a_9290_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 PAD a_8860_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X42 VSSIO a_10282_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X43 PAD a_924_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X44 PAD a_3900_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X45 VSSIO a_3338_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X46 VSSIO a_8298_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 PAD a_2908_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X48 PAD a_7868_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X49 VSSIO a_13258_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X50 VSSIO a_7306_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X51 PAD a_13820_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X52 PAD a_12828_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X53 VSSIO a_1354_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 VSSIO a_14178_1285# PAD VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X55 PAD a_5884_1285# VSSIO VSSIO sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_pddrvr_strong VCC_IO PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO
+ VSSIO_AMX FORCE_LOVOL_H FORCE_LO_H PAD PD_H_I2C m2_8958_2367# m1_9569_2540# m1_225_1760#
+ w_n1000_1958# m1_4511_2373# m1_2390_2540# m1_320_1646#
Xsky130_fd_io__nfet_con_diff_wo_abt_270v2_0 VCC_IO PAD PD_H[3] m1_9769_3898# PD_H_I2C
+ m1_7657_3898# VGND_IO m1_11193_3898# m1_11193_3898# m1_8232_3898# m1_785_3898# PD_H[3]
+ m1_12747_3898# PD_H[2] m1_2135_3898# PD_H[2] m1_785_3898# m1_9769_3898# m1_11193_3898#
+ PD_H[3] m1_8232_3898# PD_H[2] m1_785_3898# PD_H[3] m1_12747_3898# m1_9769_3898#
+ m1_8232_3898# m1_12747_3898# PD_H[3] m1_12747_3898# PD_H[3] sky130_fd_io__nfet_con_diff_wo_abt_270v2
R0 m2_11758_1638# m1_11193_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 PD_H[3] m2_7233_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 PD_H[3] m2_13193_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 m2_8935_1638# m1_8232_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_9769_3898# m2_10846_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 m2_655_1638# m1_785_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_11193_3898# m2_11329_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m1_2135_3898# m2_1565_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_8232_3898# m2_8506_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m2_10415_1638# m1_9769_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 TIE_LO_ESD m2_1848_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_7657_3898# m2_7664_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 PD_H[2] m2_6804_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 PD_H[2] m2_12763_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 TIE_LO_ESD m2_13622_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 m2_7233_1638# m1_7657_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m1_12747_3898# m2_13193_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 PD_H[2] m2_1260_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 PD_H[2] m2_897_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_2135_3898# m2_1848_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 TIE_LO_ESD m2_12189_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R22 m1_7657_3898# m2_6804_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m1_12747_3898# m2_12763_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 PD_H[2] m2_9986_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 TIE_LO_ESD m2_414_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 TIE_LO_ESD m2_9366_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 m2_13622_1638# m1_12747_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_1260_1638# m1_2135_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m1_785_3898# m2_897_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 PD_H[3] m2_11758_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 PD_H[3] m2_8935_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 m1_11193_3898# m2_12189_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 TIE_LO_ESD m2_10846_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 PD_H[3] m2_655_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 m1_9769_3898# m2_9986_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 PD_H[2] m2_11329_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 m1_785_3898# m2_414_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m1_8232_3898# m2_9366_1938# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 PD_H[3] m2_1565_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 PD_H[2] m2_8506_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 PD_H[3] m2_10415_1638# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 TIE_LO_ESD m2_7664_1637# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__com_pudrvr_weakv2 PU_H_N PAD w_258_n30# a_756_297#
X0 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 PAD PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X3 w_258_n30# PU_H_N a_756_297# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X5 w_258_n30# PU_H_N PAD w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X6 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_756_297# PU_H_N w_258_n30# w_258_n30# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
.ends

.subckt sky130_fd_io__gpio_pddrvr_strong_slowv2 PD_H PAD dw_n122_n335# w_168_168#
X0 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X1 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X2 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X3 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__res250_sub_small a_10_2# a_2142_2#
R0 a_10_2# a_2142_2# sky130_fd_pr__res_generic_po w=2 l=10.1
.ends

.subckt sky130_fd_io__res250only_small PAD ROUT
Xsky130_fd_io__res250_sub_small_0 PAD ROUT sky130_fd_io__res250_sub_small
.ends

.subckt sky130_fd_io__gpio_pddrvr_weakv2 PD_H PAD dw_n122_84# w_168_168#
X0 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X1 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X2 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X3 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X4 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
X5 w_168_168# PD_H PAD w_168_168# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_odrvr_subv2 PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD
+ FORCE_HI_H_N FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX
+ TIE_HI_ESD m3_6107_13425# sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C w_n915_9930#
+ w_588_14893# li_5884_n9263# m2_8191_n10933# w_5497_14893# sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155# VGND_IO VGND PAD VCC_IO
Xsky130_fd_io__com_pudrvr_strong_slowv2_0 PU_H_N[1] sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD
+ VCC_IO sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD sky130_fd_io__com_pudrvr_strong_slowv2
Xsky130_fd_io__com_res_weak_0 sky130_fd_io__com_res_weak_0/RB sky130_fd_io__com_res_weak_0/RA
+ sky130_fd_io__com_res_weak_0/sky130_fd_io__com_res_weak_bentbigres_0/a_n258_6046#
+ sky130_fd_io__com_res_weak_0/li_n135_8054# sky130_fd_io__com_res_weak_0/a_n160_10423#
+ sky130_fd_io__com_res_weak_0/li_n135_6820# sky130_fd_io__com_res_weak_0/a_n160_9488#
+ sky130_fd_io__com_res_weak
Xsky130_fd_io__gpio_pudrvr_strongv2_0 PU_H_N[3] PU_H_N[2] VCC_IO TIE_HI_ESD VCC_IO
+ VCC_IO PU_H_N[0] VGND VCC_IO VCC_IO VCC_IO PAD sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155# sky130_fd_io__gpio_pudrvr_strongv2
Xsky130_fd_io__gpiov2_pddrvr_strong_0 VCC_IO PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO VCC_IO
+ VCC_IO VCC_IO PAD sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C w_5497_14893# PD_H[0]
+ sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD w_n915_9930# w_588_14893# PD_H[1] sky130_fd_io__com_res_weak_0/RA
+ sky130_fd_io__gpiov2_pddrvr_strong
Xsky130_fd_io__com_pudrvr_weakv2_0 PU_H_N[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ sky130_fd_io__com_res_weak_0/RA sky130_fd_io__com_pudrvr_weakv2
Xsky130_fd_io__gpio_pddrvr_strong_slowv2_0 PD_H[1] sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD
+ VCC_IO w_588_14893# sky130_fd_io__gpio_pddrvr_strong_slowv2
Xsky130_fd_io__res250only_small_0 PAD sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__gpio_pddrvr_weakv2_0 PD_H[0] sky130_fd_io__com_res_weak_0/RA VCC_IO
+ w_5497_14893# sky130_fd_io__gpio_pddrvr_weakv2
R0 a_10314_7886# sky130_fd_io__com_res_weak_0/RB sky130_fd_pr__res_generic_po w=2 l=2
R1 a_9612_7886# a_10314_7886# sky130_fd_pr__res_generic_po w=2 l=3
R2 m1_9882_7996# a_10314_7886# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R3 a_9612_7886# m1_9882_7996# sky130_fd_pr__res_generic_m1 w=1.32 l=10m
R4 sky130_fd_io__com_pudrvr_strong_slowv2_0/PAD a_9612_7886# sky130_fd_pr__res_generic_po w=2 l=5
.ends

.subckt sky130_fd_io__gpio_odrvrv2 PAD PD_H[0] PD_H[1] PD_H[2] PD_H[3] PU_H_N[0] PU_H_N[1]
+ PU_H_N[2] PU_H_N[3] TIE_HI_ESD FORCE_HI_H_N FORCE_LO_H VSSIO_AMX w_n915_9930# FORCE_LOVOL_H
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425# TIE_LO_ESD sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C
+ w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ w_5497_14893# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ SUB VCC_IO VGND_IO
Xsky130_fd_io__gpio_odrvr_subv2_0 PD_H[0] PD_H[2] PD_H[1] PD_H[3] TIE_LO_ESD FORCE_HI_H_N
+ FORCE_LO_H FORCE_LOVOL_H PU_H_N[0] PU_H_N[1] PU_H_N[2] PU_H_N[3] VSSIO_AMX TIE_HI_ESD
+ sky130_fd_io__gpio_odrvr_subv2_0/m3_6107_13425# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpiov2_pddrvr_strong_0/PD_H_I2C
+ w_n915_9930# w_588_14893# sky130_fd_io__gpio_odrvr_subv2_0/li_5884_n9263# sky130_fd_io__gpio_odrvr_subv2_0/m2_8191_n10933#
+ w_5497_14893# sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/m1_14880_n614#
+ sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ VGND_IO SUB PAD VCC_IO sky130_fd_io__gpio_odrvr_subv2
.ends

.subckt sky130_fd_io__gpio_opathv2 HLD_I_H_N OD_H SLOW VPWR TIE_HI_ESD HLD_I_OVR_H
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ DM_H[0] DM_H_N[0] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ DM_H_N[1] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ m1_4747_14860# sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ TIE_LO_ESD sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] m2_2157_n626# sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ m1_5007_14796# DM_H[1] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ PAD sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ DM_H_N[2] VSSIO_AMX sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ OE_N OUT VPWR_KA VCC_IO sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ SUB sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ DM_H[2]
Xsky130_fd_io__gpiov2_octl_dat_0 VPWR_KA SLOW HLD_I_OVR_H OD_H sky130_fd_io__gpiov2_octl_dat_0/SLOW_H_N
+ sky130_fd_io__gpiov2_octl_dat_0/DRVHI_H sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1] sky130_fd_io__gpio_odrvrv2_0/PD_H[0]
+ sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] sky130_fd_io__gpiov2_octl_dat_0/DRVLO_H_N
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__com_pupredrvr_strong_slowv2_0/a_93_102#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12120_4573#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_13911_2980#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_18190_3078#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_261_220#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2821_220#
+ DM_H[0] DM_H[1] DM_H_N[0] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16799_2980#
+ DM_H_N[1] DM_H_N[2] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_2874_118#
+ OE_N SUB sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__gpiov2_pupredrvr_strong_nd2_0/a_158_632#
+ HLD_I_H_N DM_H[2] sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_16899_3078#
+ VPWR sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/a_1772_220#
+ OUT sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ VCC_IO sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/a_12434_3172#
+ sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3] SUB sky130_fd_io__gpiov2_octl_dat
Xsky130_fd_io__gpio_odrvrv2_0 PAD sky130_fd_io__gpio_odrvrv2_0/PD_H[0] sky130_fd_io__gpio_odrvrv2_0/PD_H[1]
+ sky130_fd_io__gpio_odrvrv2_0/PD_H[2] sky130_fd_io__gpio_odrvrv2_0/PD_H[3] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[0]
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpio_odrvrv2_0/PU_H_N[3]
+ TIE_HI_ESD VSSIO_AMX VSSIO_AMX VSSIO_AMX w_n815_25161# VSSIO_AMX SUB TIE_LO_ESD
+ sky130_fd_io__gpiov2_octl_dat_0/PD_H[4] SUB SUB SUB SUB sky130_fd_io__gpio_odrvrv2_0/sky130_fd_io__gpio_odrvr_subv2_0/sky130_fd_io__gpio_pudrvr_strongv2_0/li_9083_n155#
+ sky130_fd_io__gpio_odrvrv2_0/PU_H_N[1] SUB VCC_IO SUB sky130_fd_io__gpio_odrvrv2
.ends

.subckt sky130_fd_io__amux_switch_1v2b AMUXBUS_HV PAD_HV_P0 PG_AMX_VDDA_H_N NG_AMX_VPMP_H
+ NG_PAD_VPMP_H PAD_HV_P1 PG_PAD_VDDIOQ_H_N PAD_HV_N0 PAD_HV_N1 VSSD PAD_HV_N2 PAD_HV_N3
+ VDDIO w_7010_315# w_3919_213# VDDA
X0 PAD_HV_N0 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X1 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X2 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X3 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X4 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X5 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X6 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X7 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.96 pd=14.6 as=1.23 ps=7.35 w=7 l=0.5
X8 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X9 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X10 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X11 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X12 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X13 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X14 w_3919_213# NG_PAD_VPMP_H PAD_HV_N1 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X15 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X16 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X17 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P0 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X18 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X19 AMUXBUS_HV PG_AMX_VDDA_H_N w_3919_213# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X20 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X21 AMUXBUS_HV NG_AMX_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X22 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X23 PAD_HV_P1 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X24 PAD_HV_N2 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=2.2 ps=14.6 w=7 l=0.5
X25 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X26 PAD_HV_N3 NG_PAD_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X27 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X28 PAD_HV_N1 NG_PAD_VPMP_H w_3919_213# w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X29 w_7010_315# NG_PAD_VPMP_H PAD_HV_N2 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X30 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X31 w_7010_315# NG_AMX_VPMP_H AMUXBUS_HV w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=1.23 pd=7.35 as=1.96 ps=14.6 w=7 l=0.5
X32 w_3919_213# PG_PAD_VDDIOQ_H_N PAD_HV_P1 VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X33 w_3919_213# PG_AMX_VDDA_H_N AMUXBUS_HV VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
X34 PAD_HV_P0 PG_PAD_VDDIOQ_H_N w_3919_213# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.23 pd=7.35 as=0.98 ps=7.28 w=7 l=0.5
X35 w_3919_213# NG_AMX_VPMP_H AMUXBUS_HV w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X36 w_3919_213# NG_PAD_VPMP_H PAD_HV_N0 w_3919_213# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X37 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X38 AMUXBUS_HV NG_AMX_VPMP_H w_7010_315# w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.23 ps=7.35 w=7 l=0.5
X39 w_7010_315# NG_PAD_VPMP_H PAD_HV_N3 w_7010_315# sky130_fd_pr__nfet_g5v0d10v5 ad=2.2 pd=14.6 as=0.98 ps=7.28 w=7 l=0.5
.ends

.subckt sky130_fd_io__res75only_small PAD ROUT
R0 PAD ROUT sky130_fd_pr__res_generic_po w=2 l=3.15
.ends

.subckt sky130_fd_io__gpiov2_amx_pucsd_inv VSSA VDA Y A SUB w_1_293#
X0 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 Y A VSSA SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.6
X2 Y A VSSA SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
X3 Y A VSSA SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X4 Y A VSSA SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X5 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 VSSA A Y SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X7 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X8 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X9 VDA A Y w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X11 Y A VDA w_1_293# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 VSSA A Y SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
X13 VSSA A Y SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_amx_inv4 A VDA VSSA Y w_0_284# SUB
X0 Y A VSSA SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.6
X1 VDA A Y w_0_284# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X2 Y A VDA w_0_284# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 VSSA A Y SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_lshv2hv VPWR_HV IN RST_H HLD_H_N IN_B OUT_H_N
+ a_n1424_3030# w_n1543_3062# a_n988_3146# VGND
X0 a_472_123# IN a_n988_3146# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 a_n988_3146# a_n1424_3030# VPWR_HV w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X2 a_n1424_3030# IN_B a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X3 VGND HLD_H_N a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X4 OUT_H_N a_n1424_3030# VPWR_HV w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X5 a_n988_3146# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X6 VPWR_HV a_n988_3146# a_n1424_3030# w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X7 a_n1424_3030# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X8 a_472_123# IN_B a_n1424_3030# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X9 VPWR_HV a_n1424_3030# OUT_H_N w_n1543_3062# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X10 a_472_123# IN_B a_n1424_3030# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X11 a_n988_3146# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X12 VGND a_n1424_3030# OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_lshv2hv2 IN RST_H HLD_H_N IN_B OUT_H_N VGND
+ a_319_123# VPWR_HV a_940_123#
X0 a_472_123# IN a_940_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 VPWR_HV a_319_123# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X2 a_319_123# IN_B a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X3 VGND HLD_H_N a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X4 OUT_H_N a_319_123# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X5 a_940_123# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X6 a_319_123# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X7 a_472_123# IN_B a_319_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X8 VPWR_HV a_319_123# a_940_123# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X9 a_319_123# a_940_123# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X10 a_472_123# IN_B a_319_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X11 a_940_123# IN a_472_123# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X12 VGND a_319_123# OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr_ls VPWR_LV RST_H OUT_H_N IN IN_B HLD_H_N OUT_H
+ a_398_158# VGND a_226_158# VPWR_HV
X0 a_226_158# VPWR_LV a_594_584# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X1 OUT_H OUT_H_N VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X2 OUT_H HLD_H_N a_594_584# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X3 a_226_158# IN_B VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X4 VGND RST_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X5 a_877_584# HLD_H_N OUT_H_N VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X6 a_594_584# VPWR_LV a_226_158# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 a_594_584# HLD_H_N OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X8 VGND IN_B a_226_158# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_877_584# VPWR_LV a_398_158# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X10 a_398_158# IN VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 OUT_H_N HLD_H_N a_877_584# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X12 a_398_158# VPWR_LV a_877_584# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X13 VPWR_HV OUT_H OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X14 VGND IN a_398_158# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X15 OUT_H RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
.ends

.subckt sky130_fd_io__amx_inv1 a_66_382# a_219_36# a_66_36# a_119_10# w_0_316#
X0 a_219_36# a_119_10# a_66_382# w_0_316# sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X1 a_219_36# a_119_10# a_66_36# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_drvr D_B NMIDA_VCCD_N NMIDA_VCCD NGA_PAD_VSWITCH_H_N
+ PD_CSD_VSWITCH_H_N NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H PD_CSD_VSWITCH_H NGB_AMX_VSWITCH_H
+ NGB_PAD_VSWITCH_H AMUX_EN_VDDA_H_N NMIDA_ON_N PU_ON_N PU_ON AMUXBUSA_ON_N AMUXBUSA_ON
+ AMUX_EN_VSWITCH_H_N PGB_AMX_VDDA_H_N NGA_AMX_VSWITCH_H VDDA AMUX_EN_VDDA_H AMUXBUSB_ON_N
+ PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N m1_19989_n11490# m1_17385_n10825# sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ m2_20051_n11486# m1_16633_n11615# m2_19532_n11610# m2_17426_n12074# m1_23401_n11569#
+ m1_18679_n11104# m1_17797_n11010# m1_18365_n10924# m2_16539_n11002# m1_17392_n6692#
+ PU_CSD_VDDIOQ_H_N m1_18084_n11662# sky130_fd_io__gpiov2_amx_pucsd_inv_0/A m1_16691_n12255#
+ m1_17928_n11059# sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158# m1_19746_n11489#
+ m2_19572_n11610# m2_17903_n11844# m1_18081_n11624# m2_16473_n11654# m1_18445_n10934#
+ m1_22876_n9465# m2_20912_n11926# m2_27137_n11400# m1_18222_n11662# sky130_fd_io__gpiov2_amx_inv4_5/A
+ m1_18834_n11164# m1_17472_n6718# m1_19518_n11662# AMUXBUSB_ON sky130_fd_io__hvsbt_inv_x2_1/IN
+ m1_17059_n11489# sky130_fd_io__gpiov2_amx_inv4_1/A m1_16789_n12170# m1_18772_n11178#
+ m1_19593_n11489# sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123# m1_17927_n11010#
+ AMUX_EN_VSWITCH_H m1_19972_n11538# sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ VCCD m2_16610_n11236# m1_17797_n11059# m1_18257_n10845# PGA_AMX_VDDA_H_N sky130_fd_io__gpiov2_amx_inv4_2/A
+ m2_16539_n11154# m2_16539_n11240# m1_16635_n11564# VSSA m1_17465_n10825# m1_23228_n10198#
+ m1_17925_n10825# sky130_fd_io__gpiov2_amx_inv4_4/A m2_17841_n11844# sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ m2_16539_n11563# PD_ON m1_16576_n12293# m2_19993_n11486# sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123# AMUX_EN_VDDIO_H PD_ON_N AMUX_EN_VDDIO_H_N
+ m2_16340_n11711# sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N VDDIO_Q m2_16478_n11164#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146# m1_17795_n11868# m2_16613_n11563#
+ sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158# m1_17457_n12126# m1_16696_n12226#
+ m1_18759_n11090# li_22905_n10879# VSWITCH m2_16276_n11768# m1_18389_n10980# m2_17340_n12074#
+ m1_23054_n9427# m2_16610_n11154# sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ VSSD sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N m1_18005_n10825#
Xsky130_fd_io__gpiov2_amx_pucsd_inv_0 VSSD VDDIO_Q PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amx_pucsd_inv_0/A
+ VSSD VDDIO_Q sky130_fd_io__gpiov2_amx_pucsd_inv
Xsky130_fd_io__gpiov2_amx_inv4_0 sky130_fd_io__gpiov2_amx_inv4_1/A VSWITCH VSSA NGB_PAD_VSWITCH_H
+ VSWITCH sky130_fd_io__gpiov2_amx_inv4_0/SUB sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_1 sky130_fd_io__gpiov2_amx_inv4_1/A VSWITCH VSSA NGB_AMX_VSWITCH_H
+ VSWITCH sky130_fd_io__gpiov2_amx_inv4_1/SUB sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_2 sky130_fd_io__gpiov2_amx_inv4_2/A VDDIO_Q VSSD PGB_PAD_VDDIOQ_H_N
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_3 sky130_fd_io__gpiov2_amx_inv4_5/A VSWITCH VSSA NGA_PAD_VSWITCH_H
+ VSWITCH sky130_fd_io__gpiov2_amx_inv4_3/SUB sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_4 sky130_fd_io__gpiov2_amx_inv4_4/A VDDIO_Q VSSD PGA_PAD_VDDIOQ_H_N
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amx_inv4_5 sky130_fd_io__gpiov2_amx_inv4_5/A VSWITCH VSSA NGA_AMX_VSWITCH_H
+ VSWITCH sky130_fd_io__gpiov2_amx_inv4_5/SUB sky130_fd_io__gpiov2_amx_inv4
Xsky130_fd_io__gpiov2_amux_drvr_lshv2hv_0 VDDA sky130_fd_io__gpiov2_amx_inv4_4/A AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N PGA_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146# VSSA sky130_fd_io__gpiov2_amux_drvr_lshv2hv
Xsky130_fd_io__hvsbt_inv_x2_0 VCCD VSSD NMIDA_ON_N NMIDA_VCCD VCCD VSSD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_inv_x2_1 VCCD VSSD sky130_fd_io__hvsbt_inv_x2_1/IN D_B VCCD VSSD
+ sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0 sky130_fd_io__gpiov2_amx_inv4_2/A AMUX_EN_VDDA_H_N
+ AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N PGB_AMX_VDDA_H_N VSSA
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123# VDDA sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123#
+ sky130_fd_io__gpiov2_amux_drvr_lshv2hv2
Xsky130_fd_io__gpiov2_amux_drvr_ls_0 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amx_inv4_1/A
+ AMUXBUSB_ON AMUXBUSB_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_0/OUT_H
+ sky130_fd_io__gpiov2_amux_drvr_ls_0/a_398_158# VSSA sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_1 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ AMUXBUSB_ON AMUXBUSB_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_inv4_2/A sky130_fd_io__gpiov2_amux_drvr_ls_1/a_398_158#
+ VSSD sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158# VDDIO_Q sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_2 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ PD_ON PD_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H sky130_fd_io__gpiov2_amux_drvr_ls_2/a_398_158#
+ VSSA sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158# VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_3 VCCD AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amx_inv4_5/A
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_3/OUT_H
+ sky130_fd_io__gpiov2_amux_drvr_ls_3/a_398_158# VSSA sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_5 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_5/OUT_H_N
+ PU_ON PU_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_pucsd_inv_0/A sky130_fd_io__gpiov2_amux_drvr_ls_5/a_398_158#
+ VSSD sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158# VDDIO_Q sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__gpiov2_amux_drvr_ls_4 VCCD AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ AMUXBUSA_ON AMUXBUSA_ON_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amx_inv4_4/A m1_16634_n13366#
+ VSSD m1_16775_n13156# VDDIO_Q sky130_fd_io__gpiov2_amux_drvr_ls
Xsky130_fd_io__amx_inv1_0 VSWITCH PD_CSD_VSWITCH_H_N VSSA PD_CSD_VSWITCH_H VSWITCH
+ sky130_fd_io__amx_inv1
Xsky130_fd_io__amx_inv1_1 VSWITCH NGB_PAD_VSWITCH_H_N VSSA NGB_PAD_VSWITCH_H VSWITCH
+ sky130_fd_io__amx_inv1
Xsky130_fd_io__amx_inv1_2 VSWITCH NGA_PAD_VSWITCH_H_N VSSA NGA_PAD_VSWITCH_H VSWITCH
+ sky130_fd_io__amx_inv1
Xsky130_fd_io__hvsbt_inv_x1_0 NMIDA_VCCD_N VCCD VSSD VCCD NMIDA_VCCD VSSD sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 D_B VCCD VSSD VCCD D_B VSSD sky130_fd_io__hvsbt_inv_x1
X0 VSSA AMUX_EN_VDDIO_H_N NGB_PAD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X1 VSWITCH sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N PD_CSD_VSWITCH_H VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=2
X2 VSSA VSSA PD_CSD_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X3 PD_CSD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X4 PD_CSD_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N VSWITCH VSWITCH sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=2
X5 NGB_AMX_VSWITCH_H AMUX_EN_VDDA_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X6 PD_CSD_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X7 VSSA AMUX_EN_VDDA_H_N NGA_AMX_VSWITCH_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X8 NGA_PAD_VSWITCH_H AMUX_EN_VDDIO_H_N VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_nand5 OUT IN1 IN0 IN3 IN2 IN4 VPWR VGND
X0 VPWR IN0 OUT VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 a_59_1018# OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X2 VPWR OUT a_59_1018# VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X3 VGND a_59_1018# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.52 pd=12.3 as=0.111 ps=1.37 w=0.42 l=0.5
X4 OUT IN1 a_854_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X5 a_542_228# IN4 a_386_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 a_854_228# IN2 a_698_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X7 a_386_228# IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.471 ps=3.65 w=5 l=0.5
X8 OUT a_59_1018# VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.155 ps=1.37 w=0.42 l=0.5
X9 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X10 VGND OUT a_59_1018# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.111 ps=1.37 w=0.42 l=0.5
X11 a_698_228# IN3 a_542_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
.ends

.subckt sky130_fd_io__inv_1 VPWR VGND Y A VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.83 as=0.386 ps=2.93 w=1.12 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.263 ps=2.19 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__xor2_1 VPWR VGND A B X VNB VPB
X0 VPWR B a_293_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.479 pd=3.44 as=0.176 ps=1.54 w=1.26 l=0.15
X1 a_297_69# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=1.08 as=0.118 ps=1.12 w=0.84 l=0.15
X2 a_125_367# B a_42_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.5 as=0.334 ps=3.05 w=1.26 l=0.15
X3 VGND a_42_367# X VNB sky130_fd_pr__nfet_01v8 ad=0.479 pd=2.82 as=0.244 ps=1.42 w=0.84 l=0.15
X4 a_42_367# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.223 ps=2.21 w=0.84 l=0.15
X5 X B a_297_69# VNB sky130_fd_pr__nfet_01v8 ad=0.244 pd=1.42 as=0.101 ps=1.08 w=0.84 l=0.15
X6 a_293_367# a_42_367# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.334 pd=3.05 as=0.359 ps=3.09 w=1.26 l=0.15
X7 a_293_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.176 pd=1.54 as=0.189 ps=1.56 w=1.26 l=0.15
X8 VPWR A a_125_367# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.189 pd=1.56 as=0.151 ps=1.5 w=1.26 l=0.15
X9 VGND A a_42_367# VNB sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.118 ps=1.12 w=0.84 l=0.15
.ends

.subckt sky130_fd_io__nor2_1 VPWR VGND B Y A VNB VPB
X0 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.151 pd=1.39 as=0.33 ps=2.83 w=1.12 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=1.02 as=0.211 ps=2.05 w=0.74 l=0.15
X2 Y B a_116_368# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.83 as=0.151 ps=1.39 w=1.12 l=0.15
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.104 ps=1.02 w=0.74 l=0.15
.ends

.subckt sky130_fd_io__gpiov2_amux_nand4 OUT IN1 IN0 IN3 IN2 VPWR VGND
X0 VGND a_59_1018# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.52 pd=12.3 as=0.111 ps=1.37 w=0.42 l=0.5
X1 OUT a_59_1018# VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.155 ps=1.37 w=0.42 l=0.5
X2 OUT IN0 VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X3 a_542_228# IN3 a_386_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X4 a_59_1018# OUT VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X5 VPWR IN0 OUT VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 OUT IN1 a_698_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X7 a_386_228# IN0 VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.471 ps=3.65 w=5 l=0.5
X8 VPWR OUT a_59_1018# VPWR sky130_fd_pr__pfet_g5v0d10v5 ad=0.155 pd=1.37 as=0.14 ps=1.28 w=1 l=0.6
X9 VGND OUT a_59_1018# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.471 pd=3.65 as=0.111 ps=1.37 w=0.42 l=0.5
X10 a_698_228# IN2 a_542_228# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
.ends

.subckt sky130_fd_io__nand2_1 VPWR VGND B Y A VNB VPB
X0 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0888 pd=0.98 as=0.211 ps=2.05 w=0.74 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.319 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.168 pd=1.42 as=0.319 ps=2.81 w=1.12 l=0.15
.ends

.subckt sky130_fd_io__gpiov2_amux_decoder NMIDA_ON_N D_B PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N
+ PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N PD_ON_N PU_ON PU_ON_N AMUXBUSB_ON AMUXBUSB_ON_N
+ OUT ANALOG_EN ANALOG_POL ANALOG_SEL AMUXBUSA_ON AMUXBUSA_ON_N NGB_PAD_VSWITCH_H
+ NGA_PAD_VSWITCH_H NGB_PAD_VSWITCH_H_N NMIDA_VCCD_N PU_VDDIOQ_H_N PD_VSWITCH_H_N
+ sky130_fd_io__inv_1_4/Y sky130_fd_io__gpiov2_amux_nand5_0/IN0 sky130_fd_io__xor2_1_0/X
+ NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_nand4_0/OUT sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_nand5_1/IN0 sky130_fd_io__nor2_1_2/Y PD_ON sky130_fd_io__hvsbt_nand2_2/OUT
+ sky130_fd_io__inv_1_7/A sky130_fd_io__nor2_1_1/Y sky130_fd_io__nor2_1_2/B sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__inv_1_3/Y sky130_fd_io__xor2_1_0/A sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_2/Y
+ VCCD SUB sky130_fd_io__hvsbt_nand2_3/OUT sky130_fd_io__inv_1_14/Y
Xsky130_fd_io__gpiov2_amux_nand5_0 sky130_fd_io__inv_1_7/A PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5_0/IN0
+ NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N NGB_PAD_VSWITCH_H_N VCCD SUB sky130_fd_io__gpiov2_amux_nand5
Xsky130_fd_io__gpiov2_amux_nand5_1 sky130_fd_io__inv_1_5/A PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_nand5_1/IN0
+ NGA_PAD_VSWITCH_H_N PGB_PAD_VDDIOQ_H_N NGB_PAD_VSWITCH_H_N VCCD SUB sky130_fd_io__gpiov2_amux_nand5
Xsky130_fd_io__inv_1_10 VCCD SUB sky130_fd_io__inv_1_11/A ANALOG_POL SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nor_0 NGA_PAD_VSWITCH_H sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nand2_3/OUT
+ VCCD SUB SUB VCCD sky130_fd_io__hvsbt_nor
Xsky130_fd_io__inv_1_11 VCCD SUB sky130_fd_io__xor2_1_0/A sky130_fd_io__inv_1_11/A
+ SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nor_1 NGB_PAD_VSWITCH_H sky130_fd_io__hvsbt_nand2_1/IN1 sky130_fd_io__hvsbt_nand2_2/OUT
+ VCCD SUB SUB VCCD sky130_fd_io__hvsbt_nor
Xsky130_fd_io__inv_1_12 VCCD SUB sky130_fd_io__inv_1_12/Y sky130_fd_io__inv_1_13/Y
+ SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_13 VCCD SUB sky130_fd_io__inv_1_13/Y ANALOG_SEL SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__xor2_1_0 VCCD SUB sky130_fd_io__xor2_1_0/A sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__xor2_1_0/X SUB VCCD sky130_fd_io__xor2_1
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__inv_1_14/Y
+ NMIDA_ON_N SUB VCCD VCCD SUB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_14 VCCD SUB sky130_fd_io__inv_1_14/Y sky130_fd_io__nor2_1_2/Y
+ SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_1/IN1 sky130_fd_io__inv_1_2/Y
+ D_B SUB VCCD VCCD SUB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_0 VCCD SUB PD_ON_N PD_ON SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_2 PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N sky130_fd_io__hvsbt_nand2_2/OUT
+ SUB VCCD VCCD SUB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_1 VCCD SUB PU_ON_N PU_ON SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_2 VCCD SUB sky130_fd_io__inv_1_2/Y sky130_fd_io__inv_1_2/A SUB
+ VCCD sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_nand2_3 PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__hvsbt_nand2_3/OUT
+ SUB VCCD VCCD SUB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_3 VCCD SUB sky130_fd_io__inv_1_3/Y sky130_fd_io__inv_1_4/Y SUB
+ VCCD sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_4 VCCD SUB sky130_fd_io__inv_1_4/Y OUT SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_5 VCCD SUB PU_ON sky130_fd_io__inv_1_5/A SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__inv_1_6 VCCD SUB sky130_fd_io__inv_1_6/Y ANALOG_EN SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_0 VCCD SUB sky130_fd_io__nor2_1_0/B sky130_fd_io__inv_1_2/A
+ sky130_fd_io__inv_1_6/Y SUB VCCD sky130_fd_io__nor2_1
Xsky130_fd_io__gpiov2_amux_nand4_0 sky130_fd_io__gpiov2_amux_nand4_0/OUT PU_VDDIOQ_H_N
+ sky130_fd_io__nor2_1_2/Y NMIDA_VCCD_N PD_VSWITCH_H_N VCCD SUB sky130_fd_io__gpiov2_amux_nand4
Xsky130_fd_io__inv_1_7 VCCD SUB PD_ON sky130_fd_io__inv_1_7/A SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_1 VCCD SUB sky130_fd_io__nor2_1_1/B sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__inv_1_6/Y SUB VCCD sky130_fd_io__nor2_1
Xsky130_fd_io__nor2_1_2 VCCD SUB sky130_fd_io__nor2_1_2/B sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__inv_1_6/Y SUB VCCD sky130_fd_io__nor2_1
Xsky130_fd_io__gpiov2_amux_nand4_1 AMUXBUSB_ON_N PU_VDDIOQ_H_N sky130_fd_io__inv_1_2/A
+ D_B PD_VSWITCH_H_N VCCD SUB sky130_fd_io__gpiov2_amux_nand4
Xsky130_fd_io__inv_1_8 VCCD SUB AMUXBUSA_ON AMUXBUSA_ON_N SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__nor2_1_3 VCCD SUB sky130_fd_io__nor2_1_3/B sky130_fd_io__nor2_1_3/Y
+ sky130_fd_io__inv_1_6/Y SUB VCCD sky130_fd_io__nor2_1
Xsky130_fd_io__inv_1_9 VCCD SUB AMUXBUSB_ON AMUXBUSB_ON_N SUB VCCD sky130_fd_io__inv_1
Xsky130_fd_io__nand2_1_0 VCCD SUB sky130_fd_io__inv_1_12/Y sky130_fd_io__nor2_1_0/B
+ sky130_fd_io__xor2_1_0/X SUB VCCD sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_1 VCCD SUB sky130_fd_io__xor2_1_0/X sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__inv_1_13/Y SUB VCCD sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_2 VCCD SUB sky130_fd_io__inv_1_4/Y sky130_fd_io__nor2_1_3/B
+ sky130_fd_io__inv_1_11/A SUB VCCD sky130_fd_io__nand2_1
Xsky130_fd_io__nand2_1_3 VCCD SUB sky130_fd_io__inv_1_3/Y sky130_fd_io__nor2_1_1/B
+ sky130_fd_io__xor2_1_0/A SUB VCCD sky130_fd_io__nand2_1
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_ls IN_B OUT_H_N OUT_H HLD_H_N RST_H IN VPWR_LV
+ VGND VPWR_HV
X0 a_209_617# IN a_292_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 OUT_H_N a_141_899# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X2 a_209_617# HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X3 OUT_H a_331_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X4 a_331_899# VPWR_LV a_292_617# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X5 a_292_617# IN a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X6 a_141_899# VPWR_LV a_636_617# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 a_209_617# IN_B a_636_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 a_292_617# VPWR_LV a_331_899# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X9 a_636_617# IN_B a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 VGND HLD_H_N a_209_617# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X11 VPWR_HV a_141_899# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X12 a_209_617# IN a_292_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_636_617# VPWR_LV a_141_899# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X14 a_636_617# IN_B a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 a_141_899# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X16 a_141_899# VPWR_LV a_636_617# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X17 a_141_899# a_331_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X18 a_292_617# IN a_209_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 a_331_899# VPWR_LV a_292_617# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X20 a_209_617# IN_B a_636_617# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X21 a_292_617# VPWR_LV a_331_899# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X22 VGND a_331_899# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X23 a_331_899# a_141_899# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_209_617# HLD_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X25 VGND HLD_H_N a_209_617# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X26 a_636_617# VPWR_LV a_141_899# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_inv_1 VPWR VGND OUT IN VNB VPB
X0 OUT IN VGND VNB sky130_fd_pr__nfet_01v8 ad=0.211 pd=2.05 as=0.263 ps=2.19 w=0.74 l=0.15
X1 OUT IN VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.295 pd=2.59 as=0.345 ps=2.69 w=1 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_lshv2hv IN_B IN RST_H OUT_H_N OUT_H HLD_H a_4133_651#
+ VGND a_3512_651# VPWR_HV
X0 a_4133_651# IN a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X1 VPWR_HV a_4133_651# OUT_H VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X2 a_3665_651# IN_B a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 OUT_H_N a_3512_651# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X4 VPWR_HV a_4133_651# a_3512_651# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X5 a_3665_651# IN a_4133_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X6 a_3665_651# IN_B a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X7 a_4133_651# a_3512_651# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X8 VGND RST_H a_3512_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X9 OUT_H_N a_3512_651# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X10 VGND HLD_H a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X11 a_4133_651# IN a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X12 OUT_H a_4133_651# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X13 a_3512_651# IN_B a_3665_651# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_lshv2hv2 IN_B IN RST_H OUT_H_N OUT_H HLD_H VGND
+ a_425_1501# a_291_2921# a_693_2921# a_467_555# a_391_3019# li_1122_1924# VPWR_HV
X0 a_425_665# IN a_578_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X1 a_578_665# IN_B a_693_2921# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X2 VGND HLD_H a_578_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X3 VGND a_693_2921# OUT_H_N a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X4 VPWR_HV a_693_2921# OUT_H_N VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X5 OUT_H a_425_665# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X6 a_693_2921# IN_B a_578_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X7 a_391_3019# a_291_2921# a_425_1501# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
X8 VPWR_HV a_291_2921# a_391_3019# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X9 a_578_665# IN a_425_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X10 a_693_2921# a_425_665# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=1
X11 a_578_665# IN a_425_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X12 a_693_2921# IN_B a_578_665# a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X13 a_391_3019# a_291_2921# VPWR_HV VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X14 OUT_H a_425_665# VGND a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.5
X15 VPWR_HV a_693_2921# a_425_665# VPWR_HV sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=1
X16 a_693_2921# RST_H VGND a_467_555# sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_amux_ls ANALOG_EN HLD_I_H HLD_I_H_N VSWITCH AMUX_EN_VDDA_H_N
+ AMUX_EN_VSWITCH_H_N ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H AMUX_EN_VDDA_H
+ VDDA w_1167_10569# sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_4133_651# VCCD sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/li_1122_1924# ENABLE_VDDA_H AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921# VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_3512_651#
Xsky130_fd_io__gpiov2_amux_ctl_ls_0 sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N
+ AMUX_EN_VDDIO_H HLD_I_H_N HLD_I_H sky130_fd_io__gpiov2_amux_ctl_ls_0/IN VCCD VSSD
+ VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_ls
Xsky130_fd_io__gpiov2_amux_ctl_inv_1_0 VCCD VSSD sky130_fd_io__gpiov2_amux_ctl_ls_0/IN
+ sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
Xsky130_fd_io__gpiov2_amux_ctl_inv_1_1 VCCD VSSD sky130_fd_io__gpiov2_amux_ctl_ls_0/IN_B
+ ANALOG_EN VSSD VCCD sky130_fd_io__gpiov2_amux_ctl_inv_1
Xsky130_fd_io__gpiov2_amux_ctl_lshv2hv_0 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ AMUX_EN_VSWITCH_H_N AMUX_EN_VSWITCH_H ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_4133_651#
+ VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/a_3512_651# VSWITCH sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xsky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0 AMUX_EN_VDDIO_H_N AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ AMUX_EN_VDDA_H_N AMUX_EN_VDDA_H ENABLE_VDDA_H VSSD VSSD ENABLE_VDDA_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ VSSD sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/li_1122_1924#
+ VDDA sky130_fd_io__gpiov2_amux_ctl_lshv2hv2
X0 sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H ENABLE_VSWITCH_H VSWITCH w_1167_10569# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X1 VSSD ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.185 ps=1.93 w=0.7 l=0.6
X2 VSWITCH ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H w_1167_10569# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_amux_ctl_logic NMIDA_VCCD PD_CSD_VSWITCH_H NGB_AMX_VSWITCH_H
+ NGA_AMX_VSWITCH_H NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H PGB_AMX_VDDA_H_N HLD_I_H_N
+ HLD_I_H AMUX_EN_VDDA_H_N VDDA sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ m1_31532_n4477# sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146#
+ ANALOG_POL sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/m2_27137_n11400# sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/PD_ON sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158#
+ ANALOG_SEL sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N
+ VDDIO_Q sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ ENABLE_VDDA_H m2_37354_n6053# sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT OUT sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ PGB_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N sky130_fd_io__gpiov2_amux_drvr_0/PGB_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123#
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A
+ VCCD m1_31532_n4418# sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A
+ PGA_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H ANALOG_EN sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N
+ PU_CSD_VDDIOQ_H_N D_B sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ SUB sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT
Xsky130_fd_io__gpiov2_amux_drvr_0 D_B sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ NMIDA_VCCD sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N NGA_PAD_VSWITCH_H PD_CSD_VSWITCH_H
+ NGB_AMX_VSWITCH_H NGB_PAD_VSWITCH_H AMUX_EN_VDDA_H_N sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N sky130_fd_io__gpiov2_amux_drvr_0/PU_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/PGB_AMX_VDDA_H_N
+ NGA_AMX_VSWITCH_H VDDA sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDA_H sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ PGB_PAD_VDDIOQ_H_N PGA_PAD_VDDIOQ_H_N AMUX_EN_VDDIO_H_N VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_3/a_226_158#
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11090#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934#
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H VSWITCH
+ PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_5/a_226_158#
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934#
+ NGA_PAD_VSWITCH_H sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/m2_27137_n11400#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H VSWITCH
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON
+ D_B AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_319_123#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n1424_3030#
+ VCCD sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ PGA_AMX_VDDA_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H SUB
+ VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N VSWITCH sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H sky130_fd_io__gpiov2_amux_drvr_0/PD_ON
+ sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_0/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv2_0/a_940_123#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N
+ AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ VDDIO_Q ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_lshv2hv_0/a_n988_3146#
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/a_226_158#
+ sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11090# D_B VSWITCH sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934# sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/a_226_158#
+ SUB sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ VSWITCH sky130_fd_io__gpiov2_amux_drvr
Xsky130_fd_io__gpiov2_amux_decoder_0 sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N D_B
+ PGB_AMX_VDDA_H_N PGB_PAD_VDDIOQ_H_N PGA_AMX_VDDA_H_N PGA_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/PU_ON sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ OUT ANALOG_EN ANALOG_POL ANALOG_SEL sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N NGB_PAD_VSWITCH_H NGA_PAD_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ PU_CSD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X
+ sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y sky130_fd_io__gpiov2_amux_drvr_0/PD_ON
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/B
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_3/Y sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y VCCD SUB sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT
+ sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y sky130_fd_io__gpiov2_amux_decoder
Xsky130_fd_io__gpiov2_amux_ls_0 ANALOG_EN HLD_I_H HLD_I_H_N VSWITCH AMUX_EN_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N ENABLE_VSWITCH_H AMUX_EN_VDDIO_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDA_H
+ VDDA VSWITCH sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_ls_0/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H sky130_fd_io__gpiov2_amux_drvr_0/m1_18445_n10934#
+ VCCD sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv_0/RST_H
+ SUB VSWITCH ENABLE_VDDA_H sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/a_693_2921#
+ VDDIO_Q sky130_fd_io__gpiov2_amux_drvr_0/m1_18759_n11090# sky130_fd_io__gpiov2_amux_ls
.ends

.subckt sky130_fd_io__gpiov2_amux AMUXBUS_B AMUXBUS_A VDDA OUT HLD_I_H_N HLD_I_H ANALOG_SEL
+ ANALOG_POL sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N ENABLE_VSWITCH_H w_11765_4495#
+ ANALOG_EN w_11765_6609# a_14152_3009# VCCD PAD VSSIO_Q ENABLE_VDDA_H VSWITCH w_8674_6609#
+ a_5735_n215# w_8674_4393# VSSD VDDIO_Q
Xsky130_fd_io__amux_switch_1v2b_0 AMUXBUS_A sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small_3/ROUT VSSD sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__res75only_small_10/ROUT VDDIO_Q w_11765_6609# w_8674_6609# VDDA sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__amux_switch_1v2b_1 AMUXBUS_B sky130_fd_io__res75only_small_13/ROUT
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H sky130_fd_io__res75only_small_0/ROUT
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small_3/ROUT VSSD sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__res75only_small_10/ROUT VDDIO_Q w_11765_4495# w_8674_4393# VDDA sky130_fd_io__amux_switch_1v2b
Xsky130_fd_io__res75only_small_10 sky130_fd_io__res75only_small_10/PAD sky130_fd_io__res75only_small_10/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_11 PAD sky130_fd_io__res75only_small_10/PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_12 PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_13 PAD sky130_fd_io__res75only_small_13/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_0 PAD sky130_fd_io__res75only_small_0/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 PAD sky130_fd_io__res75only_small_3/PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD sky130_fd_io__res75only_small_3/ROUT
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_4 PAD sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_amux_ctl_logic_0 sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__amux_switch_1v2b_1/NG_AMX_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/NG_AMX_VPMP_H sky130_fd_io__amux_switch_1v2b_1/NG_PAD_VPMP_H
+ sky130_fd_io__amux_switch_1v2b_0/NG_PAD_VPMP_H sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ HLD_I_H_N HLD_I_H sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDA_H_N VDDA m1_n215_3811#
+ m1_n9_5040# sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N m1_8063_323# m2_405_5685#
+ ANALOG_POL m1_2332_3811# VSSD m1_n215_2973# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PD_ON
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_4/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_4/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_VCCD_N
+ m1_10523_323# ANALOG_SEL m1_497_8129# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PU_ON
+ ENABLE_VSWITCH_H sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_0/IN1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NGB_PAD_VSWITCH_H_N
+ VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_3/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_1/A
+ ENABLE_VDDA_H VCCD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_7/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_2/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_2/OUT
+ OUT sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NMIDA_ON_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON
+ sky130_fd_io__amux_switch_1v2b_1/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/PD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_12/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSA_ON_N
+ sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N m1_408_8055# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__xor2_1_0/X
+ VSWITCH sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_5/A
+ VCCD sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_inv4_4/A
+ sky130_fd_io__amux_switch_1v2b_0/PG_PAD_VDDIOQ_H_N sky130_fd_io__amux_switch_1v2b_0/PG_AMX_VDDA_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/NGA_PAD_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amx_pucsd_inv_0/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/Y
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/AMUX_EN_VDDIO_H_N sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_14/Y
+ m1_1492_5537# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VDDIO_H
+ ANALOG_EN sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PU_ON_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/AMUX_EN_VSWITCH_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/PD_ON_N sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/AMUXBUSB_ON
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__nor2_1_1/Y
+ VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__inv_1_2/A
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_drvr_0/sky130_fd_io__gpiov2_amux_drvr_ls_1/OUT_H_N
+ sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_decoder_0/sky130_fd_io__hvsbt_nand2_3/OUT
+ sky130_fd_io__gpiov2_amux_ctl_logic
Xsky130_fd_io__res75only_small_5 PAD sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_6 VSSD sky130_fd_io__res75only_small_6/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_7 VSSD sky130_fd_io__res75only_small_7/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_8 VSSD sky130_fd_io__res75only_small_8/ROUT sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_9 VSSD sky130_fd_io__res75only_small_9/ROUT sky130_fd_io__res75only_small
X0 VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H w_11765_6609# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X1 VSSD sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H w_8674_4393# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X2 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X3 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X4 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=4.2 ps=30.6 w=15 l=0.5
X6 VSSD a_14152_3009# w_8674_6609# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X7 w_8674_6609# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X8 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X10 VSSD a_14152_3009# w_11765_4495# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X11 w_11765_4495# sky130_fd_io__gpiov2_amux_ctl_logic_0/sky130_fd_io__gpiov2_amux_ls_0/sky130_fd_io__gpiov2_amux_ctl_lshv2hv2_0/RST_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X12 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X13 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=4.2 pd=30.6 as=2.1 ps=15.3 w=15 l=0.5
X14 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_4/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X15 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X16 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X17 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X18 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X19 w_11765_6609# sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD sky130_fd_io__res75only_small_9/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X20 VDDIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N sky130_fd_io__res75only_small_5/ROUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X21 w_11765_4495# sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__res75only_small_7/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X22 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X23 w_8674_4393# sky130_fd_io__gpiov2_amux_ctl_logic_0/D_B sky130_fd_io__res75only_small_6/ROUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X24 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X25 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X26 sky130_fd_io__res75only_small_8/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/NMIDA_VCCD w_8674_6609# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X27 w_11765_6609# a_14152_3009# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
X28 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_5/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 sky130_fd_io__res75only_small_5/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H VSSIO_Q VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X30 VSSIO_Q sky130_fd_io__gpiov2_amux_ctl_logic_0/PD_CSD_VSWITCH_H sky130_fd_io__res75only_small_4/ROUT VSSIO_Q sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X31 sky130_fd_io__res75only_small_4/ROUT sky130_fd_io__gpiov2_amux_ctl_logic_0/PU_CSD_VDDIOQ_H_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=2.1 pd=15.3 as=2.1 ps=15.3 w=15 l=0.5
X32 w_8674_4393# a_14152_3009# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_ipath_hvls OUT OUT_B MODE_NORMAL_N IN_VCCHIB INB_VCCHIB
+ IN_VDDIO MODE_VCCHIB_N MODE_NORMAL MODE_VCCHIB VSSD VDDIO_Q
X0 a_1290_2876# MODE_VCCHIB_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X1 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X2 a_1752_1955# a_1175_2172# OUT_B VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X3 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X4 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X5 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_621_2778# MODE_VCCHIB_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X8 a_2024_2876# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X9 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X10 VDDIO_Q MODE_VCCHIB_N a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X11 a_1930_201# IN_VCCHIB a_602_2876# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X12 a_621_2778# INB_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X13 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X15 VSSD MODE_VCCHIB a_1752_1955# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X16 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X17 VSSD MODE_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X18 a_621_2778# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X19 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X20 a_1290_2876# a_1175_2172# OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X21 VDDIO_Q MODE_NORMAL_N a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X22 a_1752_2267# MODE_NORMAL VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X23 a_881_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X24 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X25 a_1175_2172# a_602_2876# VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X26 VDDIO_Q MODE_NORMAL a_2911_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X27 VDDIO_Q OUT_B OUT VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X28 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X29 VDDIO_Q a_621_2778# a_602_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X30 a_2024_2876# IN_VDDIO OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X31 OUT_B a_1175_2172# a_1290_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X32 OUT_B IN_VDDIO a_1752_2267# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X33 VSSD MODE_VCCHIB a_881_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X34 a_881_201# INB_VCCHIB a_621_2778# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X35 a_602_2876# IN_VCCHIB a_1930_201# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X36 a_2911_2876# MODE_VCCHIB OUT_B VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X37 OUT OUT_B VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X38 a_1930_201# MODE_VCCHIB VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X39 OUT_B IN_VDDIO a_2024_2876# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X40 a_1175_2172# a_602_2876# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_vcchib_in_buf IN_H MODE_VCCHIB_LV_N OUT OUT_N VSSD VCCHIB
X0 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X1 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=4.58 pd=36.7 as=0.265 ps=2.53 w=1 l=0.8
X2 a_612_2476# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X3 VCCHIB MODE_VCCHIB_LV_N a_612_2476# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.25
X4 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X5 a_538_595# a_591_563# a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X6 a_446_3055# MODE_VCCHIB_LV_N VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X7 VCCHIB a_446_3055# OUT_N VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X8 VSSD a_446_3055# OUT_N VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X9 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X10 a_751_595# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X11 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X12 VCCHIB MODE_VCCHIB_LV_N a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X13 VSSD MODE_VCCHIB_LV_N a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X14 a_446_3055# a_591_563# a_612_3332# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X15 a_612_3332# a_591_563# a_446_3055# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X16 a_446_3055# a_591_563# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X17 a_751_595# a_591_563# a_538_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X18 VSSD OUT_N OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X19 VSSD IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X20 a_751_595# IN_H a_591_563# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X21 a_591_563# IN_H a_612_2476# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X22 a_591_563# IN_H a_751_595# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X23 a_538_595# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
X24 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0 ps=0 w=5 l=0.8
X25 a_612_2476# IN_H a_591_563# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X26 VSSD a_591_563# a_446_3055# VSSD sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X27 OUT OUT_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_in_buf OUT OUT_N MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H
+ VTRIP_SEL_H_N VDDIO_Q VSSD m1_n467_n748#
Xsky130_fd_io__hvsbt_nor_0 VTRIP_SEL_H li_3458_2405# MODE_NORMAL_N VDDIO_Q VSSD VSSD
+ VDDIO_Q sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VSSD VDDIO_Q
+ li_3458_2405# VSSD sky130_fd_io__hvsbt_inv_x1
X0 a_1761_1865# sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X1 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X2 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X3 VSSD a_36_n802# a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.5
X4 VDDIO_Q VDDIO_Q VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=11.5 pd=89.5 as=1.33 ps=10.5 w=5 l=0.8
X5 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X6 VDDIO_Q MODE_NORMAL_N a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X7 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X8 a_219_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X9 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X10 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=118 as=1.33 ps=10.5 w=5 l=0.8
X11 a_2385_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X12 a_36_n802# IN_H a_219_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X13 VDDIO_Q MODE_NORMAL_N a_2073_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X14 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.8
X15 a_917_1865# sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X16 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X17 VDDIO_Q a_2651_1865# OUT_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X18 OUT OUT_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X19 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X20 a_2651_1865# a_36_n802# a_2385_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.5
X21 VDDIO_Q sky130_fd_io__hvsbt_inv_x1_0/OUT a_1761_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X22 a_2073_1865# MODE_NORMAL_N VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X23 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X24 a_2651_1865# MODE_NORMAL_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X25 a_249_n802# IN_H a_36_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.8
X26 a_36_n802# IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X27 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X28 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.8
X29 a_2073_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.8
X30 a_249_n802# a_36_n802# a_2073_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.8
X31 a_249_n802# IN_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X32 VSSD IN_VT a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X33 VSSD IN_H a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=1.33 ps=10.5 w=5 l=0.8
X34 VSSD VTRIP_SEL_H_N IN_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=1
X35 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.33 ps=10.5 w=5 l=0.8
X36 VDDIO_Q sky130_fd_io__hvsbt_inv_x1_0/OUT a_917_1865# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X37 a_249_n802# a_36_n802# a_1761_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X38 a_917_1865# IN_H a_36_n802# VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X39 a_1761_1865# a_36_n802# a_249_n802# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X40 VSSD MODE_NORMAL_N a_2651_1865# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X41 a_2651_1865# a_36_n802# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X42 VSSD a_2651_1865# OUT_N VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X43 OUT OUT_N VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
.ends

.subckt sky130_fd_io__gpiov2_ipath_lvls IN_VCCHIB IN_VDDIO MODE_NORMAL_LV MODE_NORMAL_LV_N
+ MODE_VCCHIB_LV MODE_VCCHIB_LV_N OUT OUT_B VSSD a_323_2354# VCCHIB
X0 VSSD OUT_B OUT VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X1 VCCHIB MODE_NORMAL_LV_N a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X2 VCCHIB MODE_VCCHIB_LV_N a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X3 a_823_n317# MODE_NORMAL_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X4 a_1679_n317# IN_VCCHIB OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X5 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X6 a_114_2354# IN_VDDIO VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X7 a_1504_2754# IN_VCCHIB OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X8 a_323_2354# a_114_2354# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X9 a_436_2754# MODE_NORMAL_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X10 OUT_B a_323_2354# a_436_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X11 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X12 VCCHIB MODE_NORMAL_LV a_114_2354# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.25
X13 VCCHIB OUT_B OUT VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X14 a_823_n317# a_323_2354# OUT_B VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X15 a_1679_n317# MODE_VCCHIB_LV VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X16 a_2141_2754# MODE_NORMAL_LV OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X17 a_1504_2754# MODE_VCCHIB_LV_N VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X18 VSSD MODE_NORMAL_LV a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X19 VSSD MODE_VCCHIB_LV a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X20 a_316_n17# IN_VDDIO a_114_2354# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.398 ps=3.53 w=1.5 l=0.5
X21 VCCHIB MODE_VCCHIB_LV a_2141_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.25
X22 VCCHIB IN_VDDIO a_114_2354# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X23 OUT_B IN_VCCHIB a_1504_2754# VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X24 VSSD MODE_NORMAL_LV a_316_n17# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X25 OUT OUT_B VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X26 a_436_2754# a_323_2354# OUT_B VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X27 a_323_2354# a_114_2354# VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.25
X28 OUT OUT_B VCCHIB VCCHIB sky130_fd_pr__pfet_01v8 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.25
X29 OUT_B a_323_2354# a_823_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
X30 OUT_B IN_VCCHIB a_1679_n317# VSSD sky130_fd_pr__nfet_01v8 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_inbuf_lvinv_x1 IN OUT VPWR VGND
X0 VPWR IN OUT VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.25
X1 VGND IN OUT VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.25
.ends

.subckt sky130_fd_io__gpiov2_ibuf_se VTRIP_SEL_H_N VCCHIB ENABLE_VDDIO_LV MODE_NORMAL_N
+ IBUFMUX_OUT IN_VT IN_H VTRIP_SEL_H MODE_VCCHIB_N IBUFMUX_OUT_H sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ VDDIO_Q VSSD sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354#
Xsky130_fd_io__gpiov2_ipath_hvls_0 IBUFMUX_OUT_H sky130_fd_io__gpiov2_ipath_hvls_0/OUT_B
+ MODE_NORMAL_N sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N
+ sky130_fd_io__gpiov2_in_buf_0/OUT MODE_VCCHIB_N sky130_fd_io__hvsbt_nand2_1/IN1
+ sky130_fd_io__hvsbt_nand2_0/IN1 VSSD VDDIO_Q sky130_fd_io__gpiov2_ipath_hvls
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 ENABLE_VDDIO_LV sky130_fd_io__hvsbt_nand2_0/OUT
+ VSSD VCCHIB VCCHIB VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__gpiov2_vcchib_in_buf_0 IN_H sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT
+ sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT_N VSSD VCCHIB sky130_fd_io__gpiov2_vcchib_in_buf
Xsky130_fd_io__hvsbt_nand2_1 sky130_fd_io__hvsbt_nand2_1/IN1 ENABLE_VDDIO_LV sky130_fd_io__hvsbt_nand2_1/OUT
+ VSSD VCCHIB VCCHIB VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__gpiov2_in_buf_0 sky130_fd_io__gpiov2_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT_N
+ MODE_NORMAL_N IN_H IN_VT VTRIP_SEL_H VTRIP_SEL_H_N VDDIO_Q VSSD sky130_fd_io__gpiov2_in_buf_0/m1_n467_n748#
+ sky130_fd_io__gpiov2_in_buf
Xsky130_fd_io__gpiov2_ipath_lvls_0 sky130_fd_io__gpiov2_vcchib_in_buf_0/OUT sky130_fd_io__gpiov2_in_buf_0/OUT
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT sky130_fd_io__hvsbt_nand2_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT
+ sky130_fd_io__hvsbt_nand2_0/OUT IBUFMUX_OUT sky130_fd_io__gpiov2_ipath_lvls_0/OUT_B
+ VSSD sky130_fd_io__gpiov2_ipath_lvls_0/a_323_2354# VCCHIB sky130_fd_io__gpiov2_ipath_lvls
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_0 sky130_fd_io__hvsbt_nand2_1/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_0/OUT
+ VCCHIB VSSD sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__gpiov2_inbuf_lvinv_x1_1 sky130_fd_io__hvsbt_nand2_0/OUT sky130_fd_io__gpiov2_inbuf_lvinv_x1_1/OUT
+ VCCHIB VSSD sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_nand2_0/IN1 VDDIO_Q VSSD VDDIO_Q
+ MODE_VCCHIB_N VSSD sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_nand2_1/IN1 VDDIO_Q VSSD VDDIO_Q
+ MODE_NORMAL_N VSSD sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__hvsbt_nand2v2 IN1 IN0 OUT VGND VPWR SUB w_n34_415#
X0 VPWR IN1 OUT w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X1 OUT IN0 VPWR w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X2 OUT IN1 a_239_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X3 a_239_144# IN0 VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X4 VPWR IN1 OUT w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 OUT IN0 VPWR w_n34_415# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__gpiov2_ictl_logic INP_DIS_I_H_N INP_DIS_I_H INP_DIS_H_N DM_H_N[2]
+ DM_H_N[1] DM_H_N[0] IB_MODE_SEL_H_N VTRIP_SEL_H_N MODE_NORMAL_N MODE_VCCHIB_N TRIPSEL_I_H
+ TRIPSEL_I_H_N IB_MODE_SEL_H VSSD VDDIO_Q
Xsky130_fd_io__hvsbt_nand2v2_0 DM_H_N[0] DM_H_N[1] sky130_fd_io__hvsbt_nand2v2_0/OUT
+ VSSD VDDIO_Q VSSD VDDIO_Q sky130_fd_io__hvsbt_nand2v2
Xsky130_fd_io__hvsbt_nor_0 VTRIP_SEL_H_N TRIPSEL_I_H MODE_NORMAL_N VDDIO_Q VSSD VSSD
+ VDDIO_Q sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 IB_MODE_SEL_H INP_DIS_I_H_N MODE_VCCHIB_N VSSD VDDIO_Q
+ VDDIO_Q VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_1 IB_MODE_SEL_H_N INP_DIS_I_H_N MODE_NORMAL_N VSSD VDDIO_Q
+ VDDIO_Q VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_2 INP_DIS_H_N sky130_fd_io__hvsbt_nand2_3/OUT INP_DIS_I_H
+ VSSD VDDIO_Q VDDIO_Q VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_nand2_3 sky130_fd_io__hvsbt_nand2_3/IN1 DM_H_N[2] sky130_fd_io__hvsbt_nand2_3/OUT
+ VSSD VDDIO_Q VDDIO_Q VSSD sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x1_0 INP_DIS_I_H_N VDDIO_Q VSSD VDDIO_Q INP_DIS_I_H VSSD
+ sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_nand2_3/IN1 VDDIO_Q VSSD VDDIO_Q
+ sky130_fd_io__hvsbt_nand2v2_0/OUT VSSD sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 TRIPSEL_I_H_N VDDIO_Q VSSD VDDIO_Q TRIPSEL_I_H VSSD
+ sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__signal_5_sym_hv_local_5term GATE NWELLRING VGND IN m1_204_67#
+ NBODY
X0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 ad=3.73 pd=11.4 as=3.73 ps=11.4 w=5.75 l=0.6
R0 NBODY m1_534_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
R1 NWELLRING m1_204_67# sky130_fd_pr__res_generic_m1 w=0.02 l=5m
.ends

.subckt sky130_fd_io__gpiov2_buf_localesd VTRIP_SEL_H OUT_VT VDDIO_Q VSSD OUT_H IN_H
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VSSD VDDIO_Q VSSD OUT_H VDDIO_Q VSSD
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VSSD VDDIO_Q OUT_H VDDIO_Q VDDIO_Q VSSD
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 IN_H OUT_H sky130_fd_io__res250only_small
X0 OUT_H VTRIP_SEL_H OUT_VT VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__gpiov2_ipath ENABLE_VDDIO_LV OUT_H MODE_VCCHIB_N VCCHIB DM_H_N[1]
+ DM_H_N[0] DM_H_N[2] IB_MODE_SEL_H_N VTRIP_SEL_H_N PAD OUT m1_2058_35701# INP_DIS_H_N
+ VDDIO_Q IB_MODE_SEL_H SUB
Xsky130_fd_io__gpiov2_ibuf_se_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N VCCHIB
+ ENABLE_VDDIO_LV sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N OUT sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ sky130_fd_io__gpiov2_ibuf_se_0/IN_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H MODE_VCCHIB_N
+ OUT_H PAD VDDIO_Q SUB m2_15184_37210# sky130_fd_io__gpiov2_ibuf_se
Xsky130_fd_io__gpiov2_ictl_logic_0 sky130_fd_io__gpiov2_ictl_logic_0/INP_DIS_I_H_N
+ sky130_fd_io__gpiov2_ictl_logic_0/INP_DIS_I_H INP_DIS_H_N DM_H_N[2] DM_H_N[1] DM_H_N[0]
+ IB_MODE_SEL_H_N VTRIP_SEL_H_N sky130_fd_io__gpiov2_ibuf_se_0/MODE_NORMAL_N MODE_VCCHIB_N
+ sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H_N
+ IB_MODE_SEL_H SUB VDDIO_Q sky130_fd_io__gpiov2_ictl_logic
Xsky130_fd_io__gpiov2_buf_localesd_0 sky130_fd_io__gpiov2_ibuf_se_0/VTRIP_SEL_H sky130_fd_io__gpiov2_ibuf_se_0/IN_VT
+ VDDIO_Q SUB sky130_fd_io__gpiov2_ibuf_se_0/IN_H PAD sky130_fd_io__gpiov2_buf_localesd
.ends

.subckt sky130_fd_io__com_ctl_ls_en_1_v2 DM[1] VPB OUT_H_N OUT_H RST_H SET_H VPWR
+ HLD_H_N a_1150_n777# w_1114_n948# VCC_IO a_1762_n1276# a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X7 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X8 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X9 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X10 a_1150_n777# DM[1] a_992_934# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 a_634_829# a_992_934# a_1150_n777# w_1114_n948# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X22 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X23 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X24 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X25 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X26 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X27 a_1762_n1276# DM[1] a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X28 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X29 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X30 a_634_829# a_992_934# a_1762_n1276# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__com_ctl_ls_v2 OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N VPB
+ VCC_IO a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__com_ctl_lsv2 SET_H HLD_H_N OUT_H OUT_H_N RST_H IN VPWR m1_5675_1428#
+ w_5775_333# w_4727_n1281# VGND m1_5585_1428# VCC_IO
X0 a_4739_1530# HLD_H_N a_4700_968# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X1 OUT_H a_4739_1530# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X2 OUT_H_N a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X3 a_4700_638# VPWR a_4933_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X4 VGND SET_H a_4739_1530# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X5 VGND a_4739_1530# OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X6 VCC_IO a_4793_n866# a_4739_1530# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X7 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X8 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 a_4793_n866# RST_H VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X10 VGND IN a_4944_2496# VGND sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X11 a_4933_968# a_4944_2840# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X13 a_4933_638# HLD_H_N a_4793_n866# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X14 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X15 a_4700_968# VPWR a_4933_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X16 VCC_IO a_4793_n866# OUT_H_N VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X17 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_4944_2496# a_4700_638# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X20 a_4944_2840# a_4944_2496# VPWR w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X21 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.9
X22 VCC_IO a_4739_1530# a_4793_n866# w_4727_n1281# sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X23 a_4739_1530# a_4793_n866# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=1
X24 a_4933_638# VPWR a_4700_638# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_4944_2840# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X26 VGND a_4944_2840# a_4933_968# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X27 a_4793_n866# a_4739_1530# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=1
X28 a_4933_968# VPWR a_4700_968# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.9
X29 VPWR IN a_4944_2496# w_5775_333# sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X30 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 a_4700_638# a_4944_2496# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
.ends

.subckt sky130_fd_io__com_ctl_ls_1v2 OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N VPB
+ VCC_IO a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__gpiov2_ctl_lsbank VTRIP_SEL_H VTRIP_SEL INP_DIS INP_DIS_H DM[0]
+ DM_H[0] DM[2] DM_H[2] DM_H_N[2] VCC_IO STARTUP_ST_H STARTUP_RST_H OD_I_H IB_MODE_SEL_H_N
+ IB_MODE_SEL sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276# sky130_fd_io__com_ctl_lsv2_0/VCC_IO
+ DM_H[1] INP_DIS_H_N w_15552_2653# m1_2266_545# DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ HLD_I_H_N VGND IB_MODE_SEL_H VPWR
Xsky130_fd_io__com_ctl_ls_en_1_v2_0 DM[1] VPWR DM_H_N[1] DM_H[1] sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H VPWR HLD_I_H_N VPWR VPWR VCC_IO sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VGND sky130_fd_io__com_ctl_ls_en_1_v2
Xsky130_fd_io__com_ctl_ls_v2_0 DM_H_N[2] DM_H[2] DM[2] sky130_fd_io__com_ctl_ls_v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_v2_0/SET_H VPWR HLD_I_H_N VPWR VCC_IO VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_1 INP_DIS_H_N INP_DIS_H INP_DIS sky130_fd_io__com_ctl_ls_v2_1/RST_H
+ sky130_fd_io__com_ctl_ls_v2_1/SET_H VPWR HLD_I_H_N VPWR VCC_IO VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_ls_v2_2 DM_H_N[0] DM_H[0] DM[0] sky130_fd_io__com_ctl_ls_v2_2/RST_H
+ sky130_fd_io__com_ctl_ls_v2_2/SET_H VPWR HLD_I_H_N VPWR VCC_IO VGND sky130_fd_io__com_ctl_ls_v2
Xsky130_fd_io__com_ctl_lsv2_0 sky130_fd_io__com_ctl_lsv2_0/SET_H HLD_I_H_N IB_MODE_SEL_H
+ IB_MODE_SEL_H_N sky130_fd_io__com_ctl_lsv2_0/RST_H IB_MODE_SEL VPWR VGND VPWR w_15552_2653#
+ VGND VGND sky130_fd_io__com_ctl_lsv2_0/VCC_IO sky130_fd_io__com_ctl_lsv2
Xsky130_fd_io__com_ctl_ls_1v2_0 VTRIP_SEL_H_N VTRIP_SEL_H VTRIP_SEL sky130_fd_io__com_ctl_ls_1v2_0/RST_H
+ sky130_fd_io__com_ctl_ls_1v2_0/SET_H VPWR HLD_I_H_N VPWR VCC_IO VGND sky130_fd_io__com_ctl_ls_1v2
R0 m1_2266_320# sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 m1_14183_362# sky130_fd_io__com_ctl_ls_1v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R2 STARTUP_ST_H m1_6620_334# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R3 sky130_fd_io__com_ctl_lsv2_0/SET_H m2_15089_329# sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R4 m1_6420_507# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R5 STARTUP_RST_H m1_5875_412# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R6 STARTUP_ST_H m1_6148_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R7 sky130_fd_io__com_ctl_ls_v2_0/SET_H m1_10303_506# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 m1_6620_334# sky130_fd_io__com_ctl_ls_v2_1/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R9 OD_I_H m1_14183_362# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R10 m1_6148_320# sky130_fd_io__com_ctl_ls_v2_2/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R11 OD_I_H m1_10303_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R12 OD_I_H m1_10029_412# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R13 m2_15027_104# sky130_fd_io__com_ctl_lsv2_0/SET_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R14 sky130_fd_io__com_ctl_ls_v2_1/RST_H m1_6707_412# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R15 STARTUP_ST_H m1_6421_319# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R16 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14456_624# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R17 STARTUP_ST_H m1_5955_333# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R18 OD_I_H m1_14457_430# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R19 OD_I_H m2_14799_410# sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R20 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6421_356# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R21 m2_14799_410# sky130_fd_io__com_ctl_lsv2_0/RST_H sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R22 m2_15089_329# VGND sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R23 m1_14456_624# VGND sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R24 sky130_fd_io__com_ctl_ls_v2_2/RST_H m1_5955_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R25 sky130_fd_io__com_ctl_ls_1v2_0/SET_H m1_14457_467# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R26 VGND m1_10109_333# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R27 VGND m1_10302_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R28 m1_2553_412# m1_2266_545# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R29 sky130_fd_io__com_ctl_ls_v2_0/RST_H m1_10109_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R30 m1_10302_320# sky130_fd_io__com_ctl_ls_v2_0/SET_H sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R31 sky130_fd_io__com_ctl_ls_en_1_v2_0/SET_H m1_2267_506# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R32 sky130_fd_io__com_ctl_ls_1v2_0/RST_H m1_14263_617# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R33 VGND m1_2467_333# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R34 m1_2266_545# m1_2267_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R35 VGND m1_14263_654# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R36 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2467_370# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R37 sky130_fd_io__com_ctl_ls_v2_2/SET_H m1_6149_506# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R38 sky130_fd_io__com_ctl_lsv2_0/RST_H m1_14911_509# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R39 m1_10029_412# sky130_fd_io__com_ctl_ls_v2_0/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R40 OD_I_H m2_14990_104# sky130_fd_pr__res_generic_m2 w=0.26 l=10m
R41 STARTUP_RST_H m1_6149_543# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R42 sky130_fd_io__com_ctl_ls_en_1_v2_0/RST_H m1_2553_412# sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R43 VGND m1_14911_546# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R44 VGND m1_2266_320# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R45 m1_6744_412# STARTUP_RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R46 m1_5875_412# sky130_fd_io__com_ctl_ls_v2_2/RST_H sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R47 sky130_fd_io__com_ctl_ls_v2_1/SET_H m1_6420_507# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
.ends

.subckt sky130_fd_io__hvsbt_inv_x8 IN VPWR VGND OUT w_n42_416# SUB
X0 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X2 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X3 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X6 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X8 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X9 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X13 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X14 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X15 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X16 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X18 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X19 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X21 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X22 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X23 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__hvsbt_inv_x4 IN OUT w_n42_416# SUB a_66_144# a_66_482#
X0 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 a_66_144# IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X2 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X3 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X4 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X5 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X6 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X7 a_66_144# IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X8 OUT IN a_66_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X9 a_66_482# IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 OUT IN a_66_144# SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X11 OUT IN a_66_482# w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_ls OUT_H_N OUT_H IN RST_H SET_H VPWR HLD_H_N VPB VCC_IO
+ a_n17_1379#
X0 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X1 VCC_IO a_130_181# OUT_H VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X2 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X3 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X5 a_361_1391# HLD_H_N a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=0.6
X6 a_634_829# a_992_934# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X7 a_361_1391# VPWR a_128_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X8 a_n17_1379# a_634_829# a_128_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X9 OUT_H_N a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X10 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X11 a_128_1391# a_634_829# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X13 a_65_861# HLD_H_N a_957_1391# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.6
X14 OUT_H a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.6
X15 a_n17_1379# a_992_934# a_724_1391# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X16 a_65_861# a_130_181# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X17 a_724_1391# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8_lvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X18 a_n17_1379# a_65_861# a_130_181# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=1
X19 VPWR IN a_992_934# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X20 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X21 a_n17_1379# IN a_992_934# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.25
X22 a_n17_1379# a_65_861# OUT_H_N a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.6
X23 a_130_181# a_65_861# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X24 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X25 a_957_1391# VPWR a_724_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.9
X26 a_65_861# a_130_181# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=1
X27 a_634_829# a_992_934# a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_01v8 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.25
X28 a_130_181# SET_H a_n17_1379# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.42 ps=3.28 w=3 l=0.6
X29 a_724_1391# VPWR a_957_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
X30 a_n17_1379# RST_H a_65_861# a_n17_1379# sky130_fd_pr__nfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.6
X31 a_128_1391# VPWR a_361_1391# a_n17_1379# sky130_fd_pr__nfet_05v0_nvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.9
.ends

.subckt sky130_fd_io__hvsbt_inv_x8v2 IN VPWR VGND OUT w_n42_416# SUB
X0 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X1 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X2 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X3 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X4 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X5 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
X6 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X7 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X8 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X9 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X10 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X11 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X12 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X13 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X14 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X15 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.185 ps=1.93 w=0.7 l=0.6
X16 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X17 VGND IN OUT SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.185 pd=1.93 as=0.098 ps=0.98 w=0.7 l=0.6
X18 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X19 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X20 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.6
X21 OUT IN VGND SUB sky130_fd_pr__nfet_g5v0d10v5 ad=0.098 pd=0.98 as=0.098 ps=0.98 w=0.7 l=0.6
X22 OUT IN VPWR w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.6
X23 VPWR IN OUT w_n42_416# sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.6
.ends

.subckt sky130_fd_io__com_ctl_hldv2 HLD_OVR VGND HLD_I_H_N OD_I_H HLD_I_H li_8226_3758#
+ VPWR sky130_fd_io__hvsbt_nand2_0/IN1 m2_3556_4143# m1_3684_4201# sky130_fd_io__hvsbt_nand2_0/IN0
+ VCC_IO m2_3665_4182#
Xsky130_fd_io__hvsbt_inv_x8_0 sky130_fd_io__hvsbt_inv_x8_0/IN VCC_IO VGND sky130_fd_io__hvsbt_inv_x8_0/OUT
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x8
Xsky130_fd_io__hvsbt_inv_x4_0 sky130_fd_io__hvsbt_inv_x4_0/IN OD_I_H VCC_IO VGND VGND
+ VCC_IO sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__hvsbt_inv_x4_1 sky130_fd_io__hvsbt_nor_0/IN0 sky130_fd_io__hvsbt_inv_x8_0/IN
+ VCC_IO VGND VGND VCC_IO sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__hvsbt_nor_0 sky130_fd_io__hvsbt_nor_0/IN0 li_8312_3766# sky130_fd_io__com_ctl_ls_0/OUT_H
+ VCC_IO VGND VGND VCC_IO sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nor_1 OD_I_H li_8226_3758# li_8312_3766# VCC_IO VGND VGND VCC_IO
+ sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 sky130_fd_io__hvsbt_nand2_0/IN1 sky130_fd_io__hvsbt_nand2_0/IN0
+ sky130_fd_io__hvsbt_nand2_0/OUT VGND VCC_IO VCC_IO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__com_ctl_ls_0 sky130_fd_io__com_ctl_ls_0/OUT_H_N sky130_fd_io__com_ctl_ls_0/OUT_H
+ HLD_OVR sky130_fd_io__hvsbt_inv_x1_0/OUT VGND VPWR sky130_fd_io__hvsbt_nor_0/IN0
+ VPWR VCC_IO VGND sky130_fd_io__com_ctl_ls
Xsky130_fd_io__hvsbt_inv_x8v2_0 sky130_fd_io__hvsbt_inv_x8_0/IN VCC_IO VGND sky130_fd_io__hvsbt_inv_x8v2_0/OUT
+ VCC_IO VGND sky130_fd_io__hvsbt_inv_x8v2
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VCC_IO VGND VCC_IO
+ sky130_fd_io__hvsbt_nand2_0/IN0 VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_1 sky130_fd_io__hvsbt_inv_x4_0/IN VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_inv_x1_0/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__hvsbt_inv_x1_2 sky130_fd_io__hvsbt_nor_0/IN0 VCC_IO VGND VCC_IO sky130_fd_io__hvsbt_nand2_0/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
R0 HLD_I_H sky130_fd_io__hvsbt_inv_x8_0/IN sky130_fd_pr__res_generic_m1 w=0.23 l=10m
R1 sky130_fd_io__hvsbt_inv_x8v2_0/OUT HLD_I_H_N sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
R2 HLD_I_H_N sky130_fd_io__hvsbt_inv_x8_0/OUT sky130_fd_pr__res_generic_m1 w=0.23 l=0.025
.ends

.subckt sky130_fd_io__gpiov2_ctl VTRIP_SEL_H_N DM[0] DM[2] DM_H[0] HLD_OVR DM_H[2]
+ DM_H_N[1] INP_DIS INP_DIS_H_N VTRIP_SEL_H VTRIP_SEL HLD_H_N INP_STARTUP_EN_H IB_MODE_SEL_H_N
+ IB_MODE_SEL ENABLE_INP_H HLD_I_OVR_H ENABLE_H DM[1] li_11745_4176# li_18199_5031#
+ DM_H_N[0] OD_I_H IB_MODE_SEL_H sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ DM_H_N[2] DM_H[1] SUB HLD_I_H_N VPWR sky130_fd_io__com_ctl_hldv2_0/HLD_I_H VCC_IO
Xsky130_fd_io__gpiov2_ctl_lsbank_0 VTRIP_SEL_H VTRIP_SEL INP_DIS sky130_fd_io__gpiov2_ctl_lsbank_0/INP_DIS_H
+ DM[0] DM_H[0] DM[2] DM_H[2] DM_H_N[2] VCC_IO INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ OD_I_H IB_MODE_SEL_H_N IB_MODE_SEL sky130_fd_io__gpiov2_ctl_lsbank_0/sky130_fd_io__com_ctl_ls_en_1_v2_0/a_1762_n1276#
+ VCC_IO DM_H[1] INP_DIS_H_N VCC_IO OD_I_H DM_H_N[1] DM[1] DM_H_N[0] VTRIP_SEL_H_N
+ HLD_I_H_N SUB IB_MODE_SEL_H VPWR sky130_fd_io__gpiov2_ctl_lsbank
Xsky130_fd_io__com_ctl_hldv2_0 HLD_OVR SUB HLD_I_H_N OD_I_H sky130_fd_io__com_ctl_hldv2_0/HLD_I_H
+ HLD_I_OVR_H VPWR HLD_H_N OD_I_H OD_I_H ENABLE_H VCC_IO OD_I_H sky130_fd_io__com_ctl_hldv2
Xsky130_fd_io__hvsbt_nor_0 ENABLE_INP_H sky130_fd_io__gpiov2_ctl_lsbank_0/STARTUP_RST_H
+ li_11745_4176# VCC_IO SUB SUB VCC_IO sky130_fd_io__hvsbt_nor
Xsky130_fd_io__hvsbt_nand2_0 ENABLE_INP_H OD_I_H sky130_fd_io__hvsbt_nand2_0/OUT SUB
+ VCC_IO VCC_IO SUB sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__hvsbt_inv_x1_0 INP_STARTUP_EN_H VCC_IO SUB VCC_IO sky130_fd_io__hvsbt_nand2_0/OUT
+ SUB sky130_fd_io__hvsbt_inv_x1
.ends

.subckt sky130_fd_io__top_gpiov2 VSSIO_Q ANALOG_POL ENABLE_VDDIO IN_H IN ANALOG_EN
+ OUT TIE_HI_ESD PAD_A_ESD_1_H DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL
+ OE_N SLOW TIE_LO_ESD PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16869# sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16869# w_12765_14755# w_9674_14653# HLD_H_N PAD VSWITCH a_12875_50# VCCHIB
+ VDDIO VDDIO_Q VDDA AMUXBUS_B AMUXBUS_A VCCD VSSD
Xsky130_fd_io__gpio_opathv2_0 sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N sky130_fd_io__gpiov2_ctl_0/OD_I_H
+ SLOW VCCD TIE_HI_ESD sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H li_9062_7268# li_7854_5377#
+ sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__gpiov2_octl_mux_0/Y_H
+ sky130_fd_io__gpiov2_ctl_0/DM_H[0] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] li_10974_4971#
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] li_3302_6400# VSSD PAD li_7636_6398# li_3442_6400#
+ TIE_LO_ESD sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpio_odrvrv2_0/PU_H_N[2] sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N
+ li_5278_5352# VSSD sky130_fd_io__gpiov2_ctl_0/DM_H[1] li_2678_6400# PAD li_5245_3919#
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] VDDA sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpiov2_pdpredrvr_strong_0/sky130_fd_io__com_pdpredrvr_pbiasv2_0/PBIAS
+ li_4745_6400# OE_N OUT VCCHIB VDDIO sky130_fd_io__gpio_opathv2_0/sky130_fd_io__gpiov2_octl_dat_0/sky130_fd_io__gpiov2_obpredrvr_0/sky130_fd_io__gpio_pupredrvr_strongv2_0/sky130_fd_io__feascom_pupredrvr_nbiasv2_0/NBIAS
+ VSSD li_3958_5352# li_3334_5352# sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpio_opathv2
Xsky130_fd_io__gpiov2_amux_0 AMUXBUS_B AMUXBUS_A VDDA OUT sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N
+ sky130_fd_io__gpiov2_amux_0/HLD_I_H ANALOG_SEL ANALOG_POL sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ ENABLE_VSWITCH_H w_12765_14755# ANALOG_EN w_12765_16869# sky130_fd_io__gpiov2_amux_0/HLD_I_H
+ VCCD PAD VSSIO_Q ENABLE_VDDA_H VSWITCH w_9674_16869# VSSD w_9674_14653# VSSD VDDIO_Q
+ sky130_fd_io__gpiov2_amux
Xsky130_fd_io__res75only_small_0 PAD_A_ESD_1_H sky130_fd_io__res75only_small_1/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_1 sky130_fd_io__res75only_small_1/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_2 PAD_A_ESD_0_H sky130_fd_io__res75only_small_3/PAD
+ sky130_fd_io__res75only_small
Xsky130_fd_io__res75only_small_3 sky130_fd_io__res75only_small_3/PAD PAD sky130_fd_io__res75only_small
Xsky130_fd_io__gpiov2_ipath_0 ENABLE_VDDIO IN_H sky130_fd_io__gpiov2_ipath_0/MODE_VCCHIB_N
+ VCCHIB sky130_fd_io__gpiov2_ctl_0/DM_H_N[1] sky130_fd_io__gpiov2_ctl_0/DM_H_N[0]
+ sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N PAD IN VDDIO sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N
+ VDDIO_Q sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H VSSD sky130_fd_io__gpiov2_ipath
Xsky130_fd_io__gpiov2_ctl_0 sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H_N DM[0] DM[2] sky130_fd_io__gpiov2_ctl_0/DM_H[0]
+ HLD_OVR sky130_fd_io__gpiov2_ctl_0/DM_H[2] sky130_fd_io__gpiov2_ctl_0/DM_H_N[1]
+ INP_DIS sky130_fd_io__gpiov2_ctl_0/INP_DIS_H_N sky130_fd_io__gpiov2_ctl_0/VTRIP_SEL_H
+ VTRIP_SEL HLD_H_N sky130_fd_io__gpiov2_ctl_0/INP_STARTUP_EN_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H_N
+ IB_MODE_SEL ENABLE_INP_H sky130_fd_io__gpiov2_ctl_0/HLD_I_OVR_H ENABLE_H DM[1] ENABLE_H
+ PAD sky130_fd_io__gpiov2_ctl_0/DM_H_N[0] sky130_fd_io__gpiov2_ctl_0/OD_I_H sky130_fd_io__gpiov2_ctl_0/IB_MODE_SEL_H
+ VSSD sky130_fd_io__gpiov2_ctl_0/DM_H_N[2] sky130_fd_io__gpiov2_ctl_0/DM_H[1] VSSD
+ sky130_fd_io__gpiov2_ctl_0/HLD_I_H_N VCCD sky130_fd_io__gpiov2_amux_0/HLD_I_H VDDIO_Q
+ sky130_fd_io__gpiov2_ctl
R0 PAD PAD sky130_fd_pr__res_generic_m3 w=1.07 l=0.035
R1 PAD PAD sky130_fd_pr__res_generic_m3 w=12.4 l=0.035
.ends

.subckt sky130_ef_io__gpiov2_pad DM[0] IB_MODE_SEL ENABLE_H ENABLE_INP_H SLOW VTRIP_SEL
+ ENABLE_VDDIO ENABLE_VDDA_H ANALOG_POL HLD_H_N w_9674_16462# DM[1] w_12765_14348#
+ DM[2] w_9674_14246# PAD_A_ESD_1_H ENABLE_VSWITCH_H TIE_HI_ESD TIE_LO_ESD OE_N w_12765_16462#
+ VSWITCH ANALOG_SEL IN_H VDDIO INP_DIS OUT HLD_OVR VCCD PAD VCCHIB PAD_A_ESD_0_H
+ ANALOG_EN AMUXBUS_B AMUXBUS_A VDDA VDDIO_Q VSSIO_Q IN SUB
Xsky130_fd_io__top_gpiov2_0 VSSIO_Q ANALOG_POL ENABLE_VDDIO IN_H IN ANALOG_EN OUT
+ TIE_HI_ESD PAD_A_ESD_1_H DM[0] DM[1] DM[2] HLD_OVR INP_DIS ENABLE_VDDA_H VTRIP_SEL
+ OE_N SLOW TIE_LO_ESD PAD_A_ESD_0_H ANALOG_SEL ENABLE_INP_H ENABLE_H IB_MODE_SEL
+ ENABLE_VSWITCH_H sky130_fd_io__top_gpiov2_0/sky130_fd_io__overlay_gpiov2_m4_0/sky130_fd_io__top_gpio_pad_0/b_1500_19531#
+ w_9674_16462# sky130_fd_io__top_gpiov2_0/sky130_fd_io__gpiov2_amux_0/sky130_fd_io__amux_switch_1v2b_1/PG_AMX_VDDA_H_N
+ w_12765_16462# w_12765_14348# w_9674_14246# HLD_H_N PAD VSWITCH SUB VCCHIB VDDIO
+ VDDIO_Q VDDA AMUXBUS_B AMUXBUS_A VCCD SUB sky130_fd_io__top_gpiov2
.ends

.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_ESD_0_H PAD_A_ESD_1_H DM[2] DM[1]
+ DM[0] IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H OE_N TIE_HI_ESD
+ TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO ENABLE_VSWITCH_H
+ ANALOG_POL OUT VDDIO_Q w_9674_19062# HLD_H_N VSSIO_Q w_12765_19062# VCCD AMUXBUS_B
+ AMUXBUS_A VSWITCH VDDA w_12765_16948# VDDIO SUB w_9674_16846# PAD VCCHIB
Xgpio DM[0] IB_MODE_SEL ENABLE_H ENABLE_INP_H SLOW VTRIP_SEL ENABLE_VDDIO ENABLE_VDDA_H
+ ANALOG_POL HLD_H_N w_9674_19062# DM[1] w_12765_16948# DM[2] w_9674_16846# PAD_A_ESD_1_H
+ ENABLE_VSWITCH_H TIE_HI_ESD TIE_LO_ESD OE_N w_12765_19062# VSWITCH ANALOG_SEL IN_H
+ VDDIO INP_DIS OUT HLD_OVR VCCD PAD VCCHIB PAD_A_ESD_0_H ANALOG_EN AMUXBUS_B AMUXBUS_A
+ VDDA VDDIO_Q VSSIO_Q IN SUB sky130_ef_io__gpiov2_pad
.ends

.subckt sky130_fd_io__pad_esd m4_960_20017# m5_1354_20500#
R0 m4_960_20017# m5_1354_20500# sky130_fd_pr__res_generic_m5 w=253 l=0.1
.ends

.subckt sky130_fd_io__com_busses_esd sky130_fd_io__com_bus_hookup_0/VCCHIB sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_bus_hookup_0/VSSD sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_bus_hookup_0/AMUXBUS_B sky130_fd_io__com_bus_hookup_0/VDDIO
+ sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_bus_hookup_0/VSSIO_Q sky130_fd_io__com_bus_hookup_0/VDDIO_Q
Xsky130_fd_io__pad_esd_0 sky130_fd_io__pad_esd_0/m4_960_20017# sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__pad_esd
.ends

.subckt sky130_fd_io__gnd2gnd_sub_dnwl sky130_fd_io__gnd2gnd_tap_0[4]/sky130_fd_io__gnd2gnd_strap_0/li_0_0#
+ sky130_fd_io__gnd2gnd_tap_0[3]/sky130_fd_io__gnd2gnd_strap_0/li_0_0# sky130_fd_io__gnd2gnd_tap_0[2]/sky130_fd_io__gnd2gnd_strap_0/li_0_0#
+ sky130_fd_io__gnd2gnd_tap_0[1]/sky130_fd_io__gnd2gnd_strap_0/li_0_0# sky130_fd_io__gnd2gnd_tap_0[0]/sky130_fd_io__gnd2gnd_strap_0/li_0_0#
+ sky130_fd_io__gnd2gnd_tap_0[4]/SUB
.ends

.subckt sky130_fd_io__gnd2gnd_120x2_lv_isosub SUB
Xsky130_fd_io__gnd2gnd_sub_dnwl_0 SUB SUB SUB SUB SUB SUB sky130_fd_io__gnd2gnd_sub_dnwl
Xsky130_fd_io__gnd2gnd_sub_dnwl_1 SUB SUB SUB SUB SUB SUB sky130_fd_io__gnd2gnd_sub_dnwl
.ends

.subckt sky130_fd_io__top_power_lvc_wpad VSSIO_Q VCCHIB VDDA VDDIO_Q P_PAD P_CORE
+ OGC_LVC AMUXBUS_B DRN_LVC2 DRN_LVC1 SRC_BDY_LVC2 VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A
+ VSSA
Xsky130_fd_io__com_busses_esd_0 VCCHIB P_PAD VSSD P_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__gnd2gnd_120x2_lv_isosub_0 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=687 pd=3.1k as=0.7 ps=5.28 w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=25u pd=5m as=0.98 ps=7.28 w=7 l=8
X12 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X15 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X22 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R0 DRN_LVC1 a_414_306# sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X23 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X26 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X27 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X30 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
R1 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X41 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X42 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X45 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X47 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X48 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X49 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X50 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X51 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X52 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X53 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R2 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X54 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X55 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X56 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X57 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X58 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X59 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X61 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X62 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X63 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X64 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X65 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X66 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X67 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X68 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X69 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X70 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X71 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X72 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X73 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X74 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X75 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X76 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X77 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X78 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X79 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X82 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X83 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X84 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X85 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X86 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X87 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X88 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X89 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X90 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X91 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X92 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X93 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X95 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X96 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X97 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X98 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X99 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X100 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X102 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X103 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X104 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X105 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X107 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X108 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X109 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X110 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X112 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X113 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X114 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X115 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X116 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X117 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X118 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X119 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X120 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X121 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X122 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X125 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X126 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X127 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X128 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X129 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X130 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X131 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X132 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X133 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X134 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X135 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X136 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X137 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X138 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X139 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X140 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X141 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X143 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X144 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X145 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X146 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X147 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X148 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X149 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X150 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X151 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X152 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X153 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X154 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X155 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X156 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X157 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X158 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X159 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X160 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X161 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X162 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X163 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X164 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X165 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X166 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X167 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X169 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X170 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X171 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X172 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X173 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X174 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X175 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X176 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X177 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X178 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X180 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X181 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X182 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X183 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X184 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X185 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X186 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X187 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X188 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X189 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X190 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X191 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X192 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X194 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X195 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X196 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X197 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X198 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X199 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X200 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X201 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X203 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X204 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X205 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X206 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X207 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X208 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X209 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X210 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R3 a_13955_3836# DRN_LVC2 sky130_fd_pr__res_generic_po w=0.33 l=900
X212 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X213 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X214 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R4 a_2183_16816# a_1871_4484# sky130_fd_pr__res_generic_po w=0.33 l=720
X215 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X216 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X217 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X218 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X219 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X221 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X222 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X223 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X224 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X226 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X227 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X228 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X229 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X230 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X233 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X235 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X236 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X237 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X238 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X239 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X240 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X241 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X242 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X243 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X244 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X245 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X246 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X247 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X248 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X250 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X251 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X252 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X253 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X254 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X255 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X256 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X257 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X258 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X259 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X260 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X261 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X262 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X263 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X264 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X265 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X266 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X267 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X269 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X270 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X271 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X272 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X273 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X274 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X275 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X276 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X277 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X278 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X279 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X280 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X281 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X282 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X283 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X284 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X285 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X286 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X287 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X288 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X290 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X291 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X292 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X293 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X295 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X296 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X297 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X298 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X299 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X300 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X301 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X302 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X303 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X304 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X305 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X306 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X307 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X308 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X309 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X311 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X312 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X313 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X314 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X315 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X317 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X318 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X319 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X320 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X321 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X322 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X323 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X324 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X325 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X326 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X328 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X329 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X330 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X331 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X332 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X333 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X334 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X335 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X336 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X340 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X341 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X342 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X343 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X344 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X345 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X346 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X347 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X349 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X350 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X351 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X352 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X353 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X354 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X355 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X356 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X357 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X358 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X361 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X362 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X363 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X364 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X365 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X366 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X367 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X368 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X369 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X371 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X372 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X373 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X374 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X375 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X377 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X378 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X379 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X380 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X381 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X382 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X383 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X384 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X385 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X386 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X389 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X390 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X391 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X392 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X393 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X394 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X395 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X396 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X397 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X398 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X399 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X400 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X401 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X402 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X403 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X404 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X405 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X406 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X408 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X409 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X410 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X411 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X412 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X413 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X414 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X415 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X416 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X417 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X418 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X420 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X421 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X422 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X423 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X424 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X425 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X426 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X427 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X428 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X430 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.33 ps=10.5 w=5 l=4
X432 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X433 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X434 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X435 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X437 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X438 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X440 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X441 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X442 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X445 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X447 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X448 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X449 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X450 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X451 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X452 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
.ends

.subckt sky130_ef_io__vccd_lvc_clamped_pad VDDA VCCHIB AMUXBUS_B AMUXBUS_A VCCD_PAD
+ VCCD VDDIO VSWITCH VDDIO_Q SUB VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VCCD SUB
+ AMUXBUS_B VCCD VCCD SUB SUB VDDIO SUB VSWITCH VCCD AMUXBUS_A SUB sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_sc_hd__buf_16 A VGND VPWR X VNB VPB
X0 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X11 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X13 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X17 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X19 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 VGND A a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X25 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X32 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X34 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X35 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X36 VPWR A a_109_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 X a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 X a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X40 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 VPWR a_109_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X42 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND a_109_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=0.48 l=0.045
R1 VGND LO sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt constant_block zero vccd one SUB
Xconst_zero_buf const_source/LO SUB vccd zero SUB vccd sky130_fd_sc_hd__buf_16
Xconst_source SUB SUB vccd vccd const_source/HI const_source/LO sky130_fd_sc_hd__conb_1
Xconst_one_buf const_source/HI SUB vccd one SUB vccd sky130_fd_sc_hd__buf_16
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_W5U4AW c2_n3079_n3000# m4_n3179_n3100#
X0 c2_n3079_n3000# m4_n3179_n3100# sky130_fd_pr__cap_mim_m3_2 l=30 w=30
.ends

.subckt sky130_fd_sc_hvl__buf_8 A VGND VPWR X VNB VPB
X0 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X1 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X2 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 a_45_443# A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.203 ps=1.29 w=0.75 l=0.5
X4 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X5 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.203 pd=1.29 as=0.214 ps=2.07 w=0.75 l=0.5
X7 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X8 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 VPWR A a_45_443# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=2.06 as=0.428 ps=3.57 w=1.5 l=0.5
X10 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X11 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X12 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X13 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X15 VGND A a_45_443# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X16 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X17 X a_45_443# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X18 VGND a_45_443# X VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X19 X a_45_443# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X20 VPWR a_45_443# X VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X21 a_45_443# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.42 ps=2.06 w=1.5 l=0.5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ a_n683_n200# a_n189_n297# a_29_n297# a_189_n200#
+ a_n901_n200# a_247_n297# a_n407_n297# a_465_n297# a_407_n200# a_n625_n297# a_683_n297#
+ a_625_n200# a_n843_n297# w_n1101_n497# a_843_n200# a_n29_n200# a_n247_n200# a_n465_n200#
X0 a_n247_n200# a_n407_n297# a_n465_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_843_n200# a_683_n297# a_625_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X2 a_407_n200# a_247_n297# a_189_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X3 a_189_n200# a_29_n297# a_n29_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n465_n200# a_n625_n297# a_n683_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_625_n200# a_465_n297# a_407_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_n29_n200# a_n189_n297# a_n247_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X7 a_n683_n200# a_n843_n297# a_n901_n200# w_n1101_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_TGFUGS a_n792_n200# a_298_n200# a_516_n200# a_734_n200#
+ a_n926_n422# a_138_n288# a_n298_n288# a_80_n200# a_356_n288# a_n516_n288# a_574_n288#
+ a_n734_n288# a_n138_n200# a_n356_n200# a_n574_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n288# a_n792_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n288# a_516_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n288# a_80_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n288# a_n356_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n288# a_n574_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n288# a_298_n200# a_n926_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p69_S5N9F3 a_n1806_2500# a_n4122_n2932# a_n5280_2500#
+ a_2054_n2932# a_896_n2932# a_4756_2500# a_3598_n2932# a_3212_2500# a_n3736_n2932#
+ a_1668_n2932# a_n1806_n2932# a_5142_n2932# a_896_2500# a_510_n2932# a_n3350_2500#
+ a_n4508_2500# a_3212_n2932# a_n4894_2500# a_n5410_n3062# a_1282_2500# a_4756_n2932#
+ a_2826_2500# a_2826_n2932# a_n2192_n2932# a_n1034_2500# a_n2578_2500# a_n1420_2500#
+ a_n2964_2500# a_n648_n2932# a_n648_2500# a_n5280_n2932# a_n3350_n2932# a_4370_2500#
+ a_1282_n2932# a_124_n2932# a_n1420_n2932# a_n4894_n2932# a_124_2500# a_n2964_n2932#
+ a_n4122_2500# a_2054_2500# a_510_2500# a_n4508_n2932# a_4370_n2932# a_3598_2500#
+ a_3984_2500# a_2440_n2932# a_2440_2500# a_3984_n2932# a_n2192_2500# a_n3736_2500#
+ a_1668_2500# a_n262_n2932# a_n262_2500# a_n1034_n2932# a_5142_2500# a_n2578_n2932#
X0 a_n2578_n2932# a_n2578_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X1 a_n1420_n2932# a_n1420_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X2 a_n1806_n2932# a_n1806_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X3 a_3212_n2932# a_3212_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X4 a_3598_n2932# a_3598_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X5 a_n2964_n2932# a_n2964_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X6 a_2826_n2932# a_2826_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X7 a_4370_n2932# a_4370_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X8 a_3984_n2932# a_3984_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X9 a_n262_n2932# a_n262_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X10 a_n3350_n2932# a_n3350_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X11 a_n4122_n2932# a_n4122_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X12 a_n3736_n2932# a_n3736_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X13 a_5142_n2932# a_5142_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X14 a_n4894_n2932# a_n4894_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X15 a_1282_n2932# a_1282_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X16 a_4756_n2932# a_4756_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X17 a_124_n2932# a_124_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X18 a_510_n2932# a_510_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X19 a_896_n2932# a_896_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X20 a_n648_n2932# a_n648_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X21 a_n5280_n2932# a_n5280_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X22 a_n4508_n2932# a_n4508_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X23 a_n1034_n2932# a_n1034_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X24 a_n2192_n2932# a_n2192_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X25 a_2054_n2932# a_2054_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X26 a_1668_n2932# a_1668_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
X27 a_2440_n2932# a_2440_2500# a_n5410_n3062# sky130_fd_pr__res_xhigh_po_0p69 l=25
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_3YBPVB a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__schmittbuf_1 A VGND VPWR X VNB VPB
X0 X a_117_181# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.316 ps=1.45 w=0.75 l=0.5
X1 a_217_207# a_117_181# a_64_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.111 ps=1.37 w=0.42 l=0.5
X2 VPWR A a_231_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.341 pd=1.73 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND A a_217_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.316 pd=1.45 as=0.0588 ps=0.7 w=0.42 l=0.5
X4 a_78_463# VGND VNB sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.36
X5 a_64_207# VPWR VPB sky130_fd_pr__res_generic_pd__hv w=0.29 l=3.11
X6 X a_117_181# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.341 ps=1.73 w=1.5 l=0.5
X7 a_231_463# A a_117_181# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=0.5
X8 a_231_463# a_117_181# a_78_463# VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X9 a_217_207# A a_117_181# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.111 ps=1.37 w=0.42 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_PKVMTM a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPXE a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC a_80_n200# a_n272_n422# a_n138_n200# a_n80_n288#
X0 a_80_n200# a_n80_n288# a_n138_n200# a_n272_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_WRT4AW c1_n3036_n3000# m3_n3136_n3100#
X0 c1_n3036_n3000# m3_n3136_n3100# sky130_fd_pr__cap_mim_m3_1 l=30 w=30
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YEUEBV a_n792_n200# a_138_n297# a_n298_n297#
+ a_298_n200# a_356_n297# a_n516_n297# a_574_n297# a_516_n200# a_n734_n297# a_734_n200#
+ a_n80_n297# a_80_n200# a_n138_n200# a_n356_n200# a_n574_n200# w_n992_n497#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X1 a_n574_n200# a_n734_n297# a_n792_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.8
X2 a_734_n200# a_574_n297# a_516_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.8
X3 a_298_n200# a_138_n297# a_80_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X4 a_n138_n200# a_n298_n297# a_n356_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X5 a_n356_n200# a_n516_n297# a_n574_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
X6 a_516_n200# a_356_n297# a_298_n200# w_n992_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.29 ps=2.29 w=2 l=0.8
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YUHPBG a_n80_n297# a_80_n200# w_n338_n497# a_n138_n200#
X0 a_80_n200# a_n80_n297# a_n138_n200# w_n338_n497# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.8
.ends

.subckt sky130_fd_sc_hvl__inv_8 A VGND VPWR Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X1 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X2 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.157 pd=1.17 as=0.105 ps=1.03 w=0.75 l=0.5
X3 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X4 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.206 pd=2.05 as=0.105 ps=1.03 w=0.75 l=0.5
X5 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X6 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X7 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X8 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X9 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.157 ps=1.17 w=0.75 l=0.5
X10 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X11 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X12 VPWR A Y VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X13 Y A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X14 VGND A Y VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X15 Y A VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.199 ps=2.03 w=0.75 l=0.5
.ends

.subckt simple_por vdd3v3 vdd1v8 porb_h por_l porb_l vss1v8 vss3v3
Xsky130_fd_pr__cap_mim_m3_2_W5U4AW_0 vss3v3 sky130_fd_sc_hvl__schmittbuf_1_0/A sky130_fd_pr__cap_mim_m3_2_W5U4AW
Xsky130_fd_sc_hvl__buf_8_1 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vdd1v8 porb_l vss1v8
+ vdd1v8 sky130_fd_sc_hvl__buf_8
Xsky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ_0 m1_502_7653# m1_502_7653# m1_502_7653# m1_502_7653#
+ vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653# vdd3v3 m1_502_7653# m1_502_7653# m1_502_7653#
+ m1_502_7653# vdd3v3 vdd3v3 vdd3v3 m1_502_7653# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_ZEUEFZ
Xsky130_fd_pr__nfet_g5v0d10v5_TGFUGS_0 m1_721_6815# vss3v3 m1_721_6815# vss3v3 vss3v3
+ m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815# m1_721_6815#
+ vss3v3 m1_721_6815# vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_TGFUGS
Xsky130_fd_pr__res_xhigh_po_0p69_S5N9F3_0 li_3322_5813# li_1391_165# vss3v3 li_7567_165#
+ li_6023_165# vdd3v3 li_9111_165# li_8726_5813# li_1391_165# li_6795_165# li_3707_165#
+ vss3v3 li_6410_5813# li_6023_165# li_1778_5813# li_1006_5813# li_8339_165# vss3v3
+ vss3v3 li_6410_5813# li_9883_165# li_7954_5813# li_8339_165# li_2935_165# li_4094_5813#
+ li_2550_5813# li_4094_5813# li_2550_5813# li_4479_165# li_4866_5813# vss3v3 li_2163_165#
+ li_9498_5813# li_6795_165# li_5251_165# li_3707_165# li_619_165# li_5638_5813# li_2163_165#
+ li_1006_5813# li_7182_5813# li_5638_5813# li_619_165# li_9883_165# li_8726_5813#
+ li_9498_5813# li_7567_165# li_7954_5813# li_9111_165# li_3322_5813# li_1778_5813#
+ li_7182_5813# li_5251_165# li_4866_5813# li_4479_165# vss3v3 li_2935_165# sky130_fd_pr__res_xhigh_po_0p69_S5N9F3
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_0 m1_185_6573# m1_721_6815# vdd3v3 m1_2993_7658#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_1 m1_2756_6573# m1_4283_8081# vdd3v3 m1_2756_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_sc_hvl__schmittbuf_1_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 vdd3v3
+ sky130_fd_sc_hvl__inv_8_0/A vss3v3 vdd3v3 sky130_fd_sc_hvl__schmittbuf_1
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_2 m1_2756_6573# sky130_fd_sc_hvl__schmittbuf_1_0/A
+ vdd3v3 m1_6249_7690# sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__pfet_g5v0d10v5_3YBPVB_3 m1_185_6573# m1_502_7653# vdd3v3 m1_185_6573#
+ sky130_fd_pr__pfet_g5v0d10v5_3YBPVB
Xsky130_fd_pr__nfet_g5v0d10v5_PKVMTM_0 m1_2756_6573# vss3v3 vss3v3 m1_721_6815# sky130_fd_pr__nfet_g5v0d10v5_PKVMTM
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPXE_0 m1_4283_8081# m1_6249_7690# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPXE
Xsky130_fd_pr__nfet_g5v0d10v5_ZK8HQC_1 m1_185_6573# vss3v3 vss3v3 li_2550_5813# sky130_fd_pr__nfet_g5v0d10v5_ZK8HQC
Xsky130_fd_pr__cap_mim_m3_1_WRT4AW_0 sky130_fd_sc_hvl__schmittbuf_1_0/A vss3v3 sky130_fd_pr__cap_mim_m3_1_WRT4AW
Xsky130_fd_pr__pfet_g5v0d10v5_YEUEBV_0 vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ m1_4283_8081# m1_4283_8081# m1_4283_8081# vdd3v3 m1_4283_8081# m1_4283_8081# m1_4283_8081#
+ vdd3v3 m1_4283_8081# vdd3v3 m1_4283_8081# vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YEUEBV
Xsky130_fd_pr__pfet_g5v0d10v5_YUHPBG_0 m1_502_7653# m1_2993_7658# vdd3v3 vdd3v3 sky130_fd_pr__pfet_g5v0d10v5_YUHPBG
Xsky130_fd_sc_hvl__buf_8_0 sky130_fd_sc_hvl__inv_8_0/A vss3v3 vdd3v3 porb_h vss3v3
+ vdd3v3 sky130_fd_sc_hvl__buf_8
Xsky130_fd_sc_hvl__inv_8_0 sky130_fd_sc_hvl__inv_8_0/A vss1v8 vdd1v8 por_l vss1v8
+ vdd1v8 sky130_fd_sc_hvl__inv_8
.ends

.subckt sky130_fd_io__sio_clamp_pcap_4x5 a_36_36# a_229_118#
X0 a_36_36# a_229_118# a_36_36# a_36_36# sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=2.65 ps=21.1 w=5 l=4
.ends

.subckt sky130_fd_io__esd_rcclamp_nfetcap a_179_100# a_n14_18#
X0 a_n14_18# a_179_100# a_n14_18# a_n14_18# sky130_fd_pr__nfet_g5v0d10v5 ad=2.65 pd=21.1 as=1.33 ps=10.5 w=5 l=8
.ends

.subckt sky130_fd_io__hvc_clampv2 m2_5179_0# w_1040_5785# sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q w_2676_441#
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
Xsky130_fd_io__sio_clamp_pcap_4x5_0[0] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[1] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_0[2] w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCHIB
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__pad_esd_0/m5_1354_20500# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSD
+ m3_99_0# sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_A
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VCCD sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/AMUXBUS_B
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSWITCH sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSA
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDA sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VSSIO_Q
+ sky130_fd_io__com_busses_esd_0/sky130_fd_io__com_bus_hookup_0/VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1 w_2676_441# a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# w_2676_441# sky130_fd_io__esd_rcclamp_nfetcap
X0 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X1 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X3 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X5 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X6 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X7 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X8 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X9 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X10 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X11 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X12 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X13 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X14 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X15 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X16 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X18 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X21 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X22 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X23 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X24 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X25 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X26 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X27 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X28 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X29 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X30 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X31 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X32 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X33 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X37 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X38 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X39 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X40 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X41 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X42 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X44 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X45 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X46 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X47 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X48 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X50 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X51 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X52 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X53 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X54 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X55 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X57 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X58 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X59 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X60 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X61 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X62 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X63 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X64 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X65 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X66 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X67 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X68 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X69 w_2676_441# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=74.2 pd=498 as=1.33 ps=10.5 w=5 l=4
X70 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X71 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X72 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X73 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X74 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X75 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X76 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X77 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X78 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X79 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X80 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X81 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
R0 a_1672_8570# a_1268_5934# sky130_fd_pr__res_generic_po w=0.33 l=470
X82 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X83 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X84 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X85 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X86 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X87 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X88 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X89 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X90 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X91 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X92 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X93 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X94 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X95 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X96 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X97 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X98 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X99 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X100 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X101 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X102 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X103 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X104 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X105 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X106 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X107 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X108 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X109 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X110 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X112 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X113 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X114 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X115 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X116 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X117 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X118 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X119 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X120 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X121 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X122 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X123 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X124 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X125 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X126 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X127 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X128 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X129 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X130 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X131 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R1 a_214_8570# w_1040_5785# sky130_fd_pr__res_generic_po w=0.33 l=700
X133 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X134 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X136 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X137 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X138 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X139 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X140 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X141 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X142 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X143 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X144 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X145 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X146 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X147 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X148 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X149 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X150 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X151 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
R2 a_214_8570# a_1672_8570# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X152 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X153 w_2676_441# a_1268_5934# a_1368_5960# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X154 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X155 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X156 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X157 a_1368_5960# a_1268_5934# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X158 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X159 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X160 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X161 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X162 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X163 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X164 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X165 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X166 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X167 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X168 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X169 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X170 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X171 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X172 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X173 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X174 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X175 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X176 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X177 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X178 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X179 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X180 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X181 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X182 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X183 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X184 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X185 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X186 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X187 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X188 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X189 w_1040_5785# a_1268_5934# a_1368_5960# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X190 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X191 a_1368_5960# a_1268_5934# w_1040_5785# w_1040_5785# sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X192 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X193 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X194 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X195 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X196 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X197 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X198 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X199 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X200 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X201 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X202 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X203 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X204 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X205 w_1040_5785# a_1368_5960# w_2676_441# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X206 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X207 w_2676_441# a_1368_5960# w_1040_5785# w_2676_441# sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
.ends

.subckt sky130_fd_io__top_power_hvc_wpadv2 SRC_BDY_HVC OGC_HVC AMUXBUS_B VSSIO_Q P_PAD
+ VDDIO_Q P_CORE DRN_HVC VCCHIB VDDIO VDDA VCCD VSWITCH VSSA AMUXBUS_A SUB VSSIO
Xsky130_fd_io__hvc_clampv2_0 OGC_HVC DRN_HVC P_PAD VDDIO_Q AMUXBUS_B VSSIO_Q SRC_BDY_HVC
+ VDDIO VCCHIB VSSIO VDDA SUB P_CORE VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__hvc_clampv2
.ends

.subckt sky130_ef_io__vddio_hvc_clamped_pad VSSA VDDA SUB VSSIO_Q VDDIO_PAD AMUXBUS_B
+ VSWITCH AMUXBUS_A VCCD VCCHIB VDDIO VSSIO
Xsky130_fd_io__top_power_hvc_wpadv2_0 VSSIO VDDIO AMUXBUS_B VSSIO_Q VDDIO_PAD VDDIO
+ VDDIO VDDIO VCCHIB VDDIO VDDA VCCD VSWITCH VSSA AMUXBUS_A SUB VSSIO sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__top_ground_hvc_wpad G_PAD VCCHIB VDDA VDDIO_Q VSSIO_Q OGC_HVC
+ G_CORE DRN_HVC AMUXBUS_B VDDIO VSSIO VSSD VSWITCH VCCD AMUXBUS_A VSSA SRC_BDY_HVC
Xsky130_fd_io__sio_clamp_pcap_4x5_0 SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__sio_clamp_pcap_4x5_1[0] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[1] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__sio_clamp_pcap_4x5_1[2] SRC_BDY_HVC a_1268_5934# sky130_fd_io__sio_clamp_pcap_4x5
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|0] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|1] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|2] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|3] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[0|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[1|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
Xsky130_fd_io__esd_rcclamp_nfetcap_0[2|4] a_1268_5934# SRC_BDY_HVC sky130_fd_io__esd_rcclamp_nfetcap
X0 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
X1 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X2 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X3 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X4 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X5 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X6 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X7 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X8 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X9 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X10 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X11 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X12 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X13 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X14 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X15 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X16 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X17 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X18 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X19 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X20 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X21 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X22 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X23 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X24 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X25 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X26 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X27 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X28 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X29 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X30 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X31 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X32 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X33 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X34 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X35 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X36 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X37 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X38 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X39 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X40 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X41 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X42 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X43 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X44 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X45 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X46 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X47 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X48 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X49 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X50 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X51 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X52 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X53 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X54 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X55 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X56 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X57 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X58 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X59 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X60 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X61 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X62 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X63 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X64 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X65 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X66 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X67 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X68 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X69 SRC_BDY_HVC a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=685 pd=2.25k as=1.33 ps=10.5 w=5 l=4
X70 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X71 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X72 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X73 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X74 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X75 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X76 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X77 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X78 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X79 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X80 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X81 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X82 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X83 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X84 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X85 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X86 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X87 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X88 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X89 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X90 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X91 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X92 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X93 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X94 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X95 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X96 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X97 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X98 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X99 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X100 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X101 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X102 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X103 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X104 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X105 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X106 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X107 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X108 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X109 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X110 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X111 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X112 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X113 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X114 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X115 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X116 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X117 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X118 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X119 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X120 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X121 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X122 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X123 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X124 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X125 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X126 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X127 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X128 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X129 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X130 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X131 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X132 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
R0 a_214_8638# DRN_HVC sky130_fd_pr__res_generic_po w=0.33 l=700
X133 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X134 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X135 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X136 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X137 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X138 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X139 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X140 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X141 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X142 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X143 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X144 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X145 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X146 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X147 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X148 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X149 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X150 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X151 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=1.86 pd=14.5 as=0.98 ps=7.28 w=7 l=0.5
R1 a_214_8638# a_1672_8638# sky130_fd_pr__res_generic_po w=0.33 l=1.55k
X152 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X153 SRC_BDY_HVC a_1268_5934# a_1368_5960# SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X154 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X155 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=1.86 ps=14.5 w=7 l=0.5
X156 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X157 a_1368_5960# a_1268_5934# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X158 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
R2 a_1672_8638# a_1268_5934# sky130_fd_pr__res_generic_po w=0.33 l=470
X159 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X160 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X161 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X162 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X163 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X164 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X165 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X166 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X167 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X168 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X169 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X170 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X171 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X172 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X173 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X174 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X175 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X176 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X177 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X178 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X179 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X180 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X181 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X182 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X183 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X184 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X185 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X186 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X187 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X188 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X189 DRN_HVC a_1268_5934# a_1368_5960# DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X190 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X191 a_1368_5960# a_1268_5934# DRN_HVC DRN_HVC sky130_fd_pr__pfet_g5v0d10v5 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.5
X192 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X193 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X194 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X195 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X196 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=6.95 pd=21.4 as=7.55 ps=11.5 w=10 l=0.5
X197 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X198 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X199 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X200 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=15.1 pd=21.5 as=13.9 ps=41.4 w=20 l=0.5
X201 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X202 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X203 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X204 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X205 DRN_HVC a_1368_5960# SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=7.55 pd=11.5 as=6.95 ps=21.4 w=10 l=0.5
X206 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
X207 SRC_BDY_HVC a_1368_5960# DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 ad=13.9 pd=41.4 as=15.1 ps=21.5 w=20 l=0.5
.ends

.subckt sky130_ef_io__vssio_hvc_clamped_pad VDDA SUB VSSA AMUXBUS_B AMUXBUS_A VSSIO_PAD
+ VDDIO VDDIO_Q VSSIO VSWITCH VCCHIB VCCD
Xsky130_fd_io__top_ground_hvc_wpad_0 VSSIO_PAD VCCHIB VDDA VDDIO_Q VSSIO VDDIO VSSIO
+ VDDIO AMUXBUS_B VDDIO VSSIO SUB VSWITCH VCCD AMUXBUS_A VSSA VSSIO sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt sky130_ef_io__vdda_hvc_clamped_pad VSSIO_Q VDDA_PAD VSSIO VCCHIB VSWITCH AMUXBUS_B
+ AMUXBUS_A VDDIO_Q VCCD VDDA SUB VSSA VDDIO
Xsky130_fd_io__top_power_hvc_wpadv2_0 VSSA VDDIO AMUXBUS_B VSSIO_Q VDDA_PAD VDDIO_Q
+ VDDA VDDA VCCHIB VDDIO VDDA VCCD VSWITCH VSSA AMUXBUS_A SUB VSSIO sky130_fd_io__top_power_hvc_wpadv2
.ends

.subckt sky130_fd_io__top_ground_lvc_wpad VSSIO_Q VCCHIB VDDA VDDIO_Q G_PAD G_CORE
+ OGC_LVC AMUXBUS_B DRN_LVC2 DRN_LVC1 SRC_BDY_LVC2 VSSIO VDDIO VSSD VSWITCH VCCD AMUXBUS_A
+ VSSA
Xsky130_fd_io__com_busses_esd_0 VCCHIB G_PAD VSSD G_CORE AMUXBUS_A VCCD AMUXBUS_B
+ VDDIO VSSIO VSWITCH VSSA VDDA VSSIO_Q VDDIO_Q sky130_fd_io__com_busses_esd
Xsky130_fd_io__gnd2gnd_120x2_lv_isosub_0 VSSD sky130_fd_io__gnd2gnd_120x2_lv_isosub
X0 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X1 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X2 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X3 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=687 pd=3.1k as=0.7 ps=5.28 w=5 l=8
X4 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X5 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X6 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X7 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X8 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X9 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X10 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X11 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=25u pd=5m as=0.98 ps=7.28 w=7 l=8
X12 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X13 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X14 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X15 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X16 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X17 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X18 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X19 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X20 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X21 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X22 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R0 DRN_LVC1 a_414_306# sky130_fd_pr__res_generic_po w=0.33 l=1.95k
X23 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X24 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X25 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X26 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X27 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X28 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X29 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X30 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X31 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X32 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X33 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X34 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X35 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X36 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X37 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X38 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X39 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X40 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
R1 a_2183_16816# a_2595_15129# sky130_fd_pr__res_generic_po w=0.33 l=200
X41 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X42 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X43 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X44 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X45 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X46 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X47 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X48 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X49 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X50 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X51 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X52 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X53 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
R2 a_1871_4484# a_13955_3836# sky130_fd_pr__res_generic_po w=0.33 l=300
X54 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X55 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X56 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X57 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X58 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X59 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X60 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X61 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X62 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X63 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X64 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X65 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X66 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X67 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X68 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X69 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X70 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X71 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X72 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X73 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X74 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X75 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X76 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X77 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X78 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X79 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X80 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X81 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X82 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X83 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X84 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X85 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X86 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X87 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X88 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X89 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X90 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X91 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X92 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X93 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X94 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X95 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X96 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X97 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X98 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X99 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X100 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X101 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X102 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X103 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X104 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X105 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X106 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X107 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X108 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X109 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X110 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X111 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X112 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X113 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X114 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X115 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X116 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X117 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X118 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X119 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X120 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X121 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X122 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X123 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X124 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X125 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X126 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X127 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X128 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X129 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X130 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X131 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X132 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X133 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X134 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X135 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X136 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X137 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X138 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X139 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X140 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X141 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X142 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X143 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X144 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X145 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X146 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X147 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X148 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X149 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X150 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X151 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X152 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X153 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X154 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X155 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X156 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X157 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X158 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X159 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X160 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X161 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X162 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X163 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X164 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X165 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X166 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X167 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X168 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X169 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X170 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X171 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X172 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X173 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X174 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X175 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X176 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X177 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X178 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X179 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X180 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X181 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X182 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X183 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X184 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X185 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X186 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X187 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X188 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X189 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X190 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X191 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X192 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X193 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X194 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X195 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X196 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X197 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X198 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X199 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X200 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X201 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X202 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X203 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X204 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.7 pd=5.28 as=0 ps=0 w=5 l=8
X205 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X206 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X207 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X208 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X209 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X210 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X211 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R3 a_13955_3836# DRN_LVC2 sky130_fd_pr__res_generic_po w=0.33 l=900
X212 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X213 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X214 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
R4 a_2183_16816# a_1871_4484# sky130_fd_pr__res_generic_po w=0.33 l=720
X215 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X216 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X217 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X218 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X219 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X220 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X221 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X222 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X223 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X224 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X225 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X226 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X227 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X228 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X229 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X230 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X231 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X232 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X233 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X234 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X235 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X236 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X237 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X238 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X239 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X240 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X241 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X242 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X243 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X244 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X245 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X246 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X247 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X248 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X249 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X250 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X251 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X252 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X253 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X254 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X255 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X256 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X257 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X258 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X259 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X260 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X261 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X262 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X263 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X264 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X265 SRC_BDY_LVC2 a_2595_15129# a_2872_5340# SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X266 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X267 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X268 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X269 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X270 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X271 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X272 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X273 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X274 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X275 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X276 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X277 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X278 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X279 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X280 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X281 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X282 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X283 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X284 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X285 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X286 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X287 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X288 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X289 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X290 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X291 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X292 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X293 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X294 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X295 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X296 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X297 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X298 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X299 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X300 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X301 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X302 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X303 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X304 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X305 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X306 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X307 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X308 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X309 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X310 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X311 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X312 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X313 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X314 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X315 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X316 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X317 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X318 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X319 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X320 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=1.96 pd=14.6 as=0.98 ps=7.28 w=7 l=0.18
X321 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X322 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X323 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X324 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X325 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X326 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X327 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X328 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X329 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X330 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X331 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X332 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X333 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X334 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X335 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X336 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X337 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X338 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X339 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X340 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X341 VSSD a_414_306# a_450_404# VSSD sky130_fd_pr__nfet_01v8 ad=2.4 pd=7.68 as=4.76 ps=15.4 w=7 l=0.18
X342 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=2.4 ps=7.68 w=7 l=8
X343 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X344 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X345 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X346 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X347 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X348 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X349 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X350 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X351 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X352 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X353 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X354 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X355 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X356 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X357 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X358 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X359 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X360 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X361 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=1.96 ps=14.6 w=7 l=0.18
X362 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X363 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X364 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X365 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X366 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X367 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X368 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X369 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X370 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X371 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X372 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X373 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X374 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X375 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X376 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X377 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X378 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X379 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X380 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X381 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X382 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X383 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X384 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0.98 pd=7.28 as=0 ps=0 w=7 l=8
X385 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X386 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X387 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X388 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X389 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X390 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X391 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X392 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X393 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X394 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X395 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=5.62 pd=12.2 as=2.92 ps=6.17 w=5 l=0.18
X396 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X397 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X398 a_450_404# a_414_306# DRN_LVC1 DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X399 a_2872_5340# a_2595_15129# DRN_LVC2 DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X400 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X401 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X402 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X403 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X404 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X405 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X406 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X407 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X408 VSSD a_414_306# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=8
X409 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X410 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X411 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X412 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X413 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.7 ps=5.28 w=5 l=8
X414 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X415 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X416 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X417 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X418 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X419 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X420 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X421 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X422 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X423 DRN_LVC1 a_414_306# a_450_404# DRN_LVC1 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X424 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X425 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X426 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X427 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X428 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X429 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X430 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X431 SRC_BDY_LVC2 a_2595_15129# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=1.33 ps=10.5 w=5 l=4
X432 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X433 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X434 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X435 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X436 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X437 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
X438 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X439 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X440 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X441 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X442 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=2.92 pd=6.17 as=5.62 ps=12.2 w=5 l=0.18
X443 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X444 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X445 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=3.54 pd=8.01 as=3.5 ps=15 w=7 l=0.18
X446 SRC_BDY_LVC2 a_2872_5340# DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.5 pd=11 as=2.53 ps=6.01 w=5 l=0.18
X447 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X448 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=7.88 pd=16.2 as=4.09 ps=8.17 w=7 l=0.18
X449 DRN_LVC2 a_2595_15129# a_2872_5340# DRN_LVC2 sky130_fd_pr__pfet_01v8 ad=0.98 pd=7.28 as=0.98 ps=7.28 w=7 l=0.18
X450 DRN_LVC2 a_2872_5340# SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 ad=2.53 pd=6.01 as=2.5 ps=11 w=5 l=0.18
X451 VSSD a_450_404# DRN_LVC1 VSSD sky130_fd_pr__nfet_01v8 ad=3.5 pd=15 as=3.54 ps=8.01 w=7 l=0.18
X452 DRN_LVC1 a_450_404# VSSD VSSD sky130_fd_pr__nfet_01v8 ad=4.09 pd=8.17 as=7.88 ps=16.2 w=7 l=0.18
.ends

.subckt sky130_ef_io__vssd_lvc_clamped3_pad VSSA VDDA VSWITCH VSSD_PAD VCCD1 VSSIO_Q
+ VDDIO VCCHIB VCCD AMUXBUS_B VDDIO_Q AMUXBUS_A SUB
Xsky130_fd_io__top_ground_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD SUB SUB
+ AMUXBUS_B VCCD1 VCCD1 SUB SUB VDDIO SUB VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_ground_lvc_wpad
.ends

.subckt sky130_ef_io__vssd_lvc_clamped_pad VDDA VSWITCH VSSD_PAD VDDIO VCCD AMUXBUS_B
+ AMUXBUS_A VDDIO_Q VCCHIB VSSIO_Q SUB
Xsky130_fd_io__top_ground_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VSSD_PAD SUB SUB
+ AMUXBUS_B VCCD VCCD SUB SUB VDDIO SUB VSWITCH VCCD AMUXBUS_A SUB sky130_fd_io__top_ground_lvc_wpad
.ends

.subckt sky130_ef_io__vccd_lvc_clamped3_pad VDDA VCCHIB VDDIO VSWITCH AMUXBUS_B AMUXBUS_A
+ VCCD VCCD_PAD VCCD1 SUB VSSA VDDIO_Q VSSIO_Q
Xsky130_fd_io__top_power_lvc_wpad_0 VSSIO_Q VCCHIB VDDA VDDIO_Q VCCD_PAD VCCD1 SUB
+ AMUXBUS_B VCCD1 VCCD1 SUB SUB VDDIO SUB VSWITCH VCCD AMUXBUS_A VSSA sky130_fd_io__top_power_lvc_wpad
.ends

.subckt sky130_fd_sc_hvl__decap_4 VGND VPWR VNB VPB
X0 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.412 pd=4.1 as=0.199 ps=2.03 w=0.75 l=1
X1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.55 pd=5.1 as=0.265 ps=2.53 w=1 l=1
.ends

.subckt sky130_fd_sc_hvl__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=7.68 as=0.275 ps=2.55 w=1 l=1
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.623 pd=6.16 as=0.199 ps=2.03 w=0.75 l=1
X2 VPWR VGND VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.14 ps=1.28 w=1 l=1
X3 VGND VPWR VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0 ps=0 w=0.75 l=1
.ends

.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VPB VPWR VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_11v0 pj=3.16 area=0.607
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A VGND VPWR X VNB VPB LVPWR
X0 a_30_1337# A VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X1 VGND a_30_1337# a_30_207# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X2 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X3 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X4 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X5 VGND a_30_207# a_389_141# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X6 VGND A a_30_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X7 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X8 a_389_141# a_30_207# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X9 VGND a_30_1337# a_389_1337# VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X10 LVPWR a_389_141# X LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.4 as=0.297 ps=2.77 w=1.12 l=0.15
X11 VGND a_389_141# X VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=2.01 as=0.196 ps=2.01 w=0.74 l=0.15
X12 a_389_1337# a_30_1337# VGND VNB sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X13 LVPWR a_389_1337# a_389_141# LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.297 ps=2.77 w=1.12 l=0.15
X14 a_30_207# a_30_1337# VPWR VPB sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X15 a_389_1337# a_389_141# LVPWR LVPWR sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.157 ps=1.4 w=1.12 l=0.15
.ends

.subckt xres_buf A X LVPWR LVGND VPWR VGND
XFILLER_0_24 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_16 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_4
XANTENNA_lvlshiftdown_A A VGND VPWR VPWR VGND sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_0 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_8 VGND VPWR VGND VPWR sky130_fd_sc_hvl__decap_8
Xlvlshiftdown A VGND VPWR X VGND VPWR LVPWR sky130_fd_sc_hvl__lsbufhv2lv_1
.ends

.subckt sky130_ef_io__vssa_hvc_clamped_pad SUB VDDIO VSSA_PAD VSSA VCCHIB VSWITCH
+ VSSIO VDDIO_Q VDDA VCCD VSSIO_Q AMUXBUS_A AMUXBUS_B
Xsky130_fd_io__top_ground_hvc_wpad_0 VSSA_PAD VCCHIB VDDA VDDIO_Q VSSIO_Q VDDIO VSSA
+ VDDA AMUXBUS_B VDDIO VSSIO SUB VSWITCH VCCD AMUXBUS_A VSSA VSSA sky130_fd_io__top_ground_hvc_wpad
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.452 pd=4.52 as=0.226 ps=2.26 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.286 pd=3.24 as=0.143 ps=1.62 w=0.55 l=1.97
.ends

.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[14]
+ mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20]
+ mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27]
+ mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5]
+ mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[28] mask_rev[13] SUB VPWR
Xmask_rev_value\[1\] SUB SUB VPWR VPWR mask_rev_value\[1\]/HI mask_rev[1] sky130_fd_sc_hd__conb_1
XFILLER_6_12 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[30\] SUB SUB VPWR VPWR mask_rev_value\[30\]/HI mask_rev[30] sky130_fd_sc_hd__conb_1
XFILLER_0_47 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[23\] SUB SUB VPWR VPWR mask_rev_value\[23\]/HI mask_rev[23] sky130_fd_sc_hd__conb_1
XFILLER_0_15 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[16\] SUB SUB VPWR VPWR mask_rev_value\[16\]/HI mask_rev[16] sky130_fd_sc_hd__conb_1
XFILLER_0_39 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[21\] SUB SUB VPWR VPWR mask_rev_value\[21\]/HI mask_rev[21] sky130_fd_sc_hd__conb_1
XFILLER_3_6 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_28 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XPHY_0 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_18 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[14\] SUB SUB VPWR VPWR mask_rev_value\[14\]/HI mask_rev[14] sky130_fd_sc_hd__conb_1
XPHY_1 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[8\] SUB SUB VPWR VPWR mask_rev_value\[8\]/HI mask_rev[8] sky130_fd_sc_hd__conb_1
XPHY_2 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_6 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XPHY_3 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[12\] SUB SUB VPWR VPWR mask_rev_value\[12\]/HI mask_rev[12] sky130_fd_sc_hd__conb_1
XPHY_4 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_10 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[6\] SUB SUB VPWR VPWR mask_rev_value\[6\]/HI mask_rev[6] sky130_fd_sc_hd__conb_1
XFILLER_1_33 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XPHY_5 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XPHY_6 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[28\] SUB SUB VPWR VPWR mask_rev_value\[28\]/HI mask_rev[28] sky130_fd_sc_hd__conb_1
XFILLER_8_3 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[10\] SUB SUB VPWR VPWR mask_rev_value\[10\]/HI mask_rev[10] sky130_fd_sc_hd__conb_1
XFILLER_1_24 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XPHY_7 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_46 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[4\] SUB SUB VPWR VPWR mask_rev_value\[4\]/HI mask_rev[4] sky130_fd_sc_hd__conb_1
XFILLER_7_46 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
XPHY_8 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XPHY_9 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_26 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[26\] SUB SUB VPWR VPWR mask_rev_value\[26\]/HI mask_rev[26] sky130_fd_sc_hd__conb_1
XFILLER_6_3 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_15 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[19\] SUB SUB VPWR VPWR mask_rev_value\[19\]/HI mask_rev[19] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[2\] SUB SUB VPWR VPWR mask_rev_value\[2\]/HI mask_rev[2] sky130_fd_sc_hd__conb_1
XFILLER_7_27 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[31\] SUB SUB VPWR VPWR mask_rev_value\[31\]/HI mask_rev[31] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[24\] SUB SUB VPWR VPWR mask_rev_value\[24\]/HI mask_rev[24] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[17\] SUB SUB VPWR VPWR mask_rev_value\[17\]/HI mask_rev[17] sky130_fd_sc_hd__conb_1
XFILLER_5_40 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
Xmask_rev_value\[0\] SUB SUB VPWR VPWR mask_rev_value\[0\]/HI mask_rev[11] sky130_fd_sc_hd__conb_1
XFILLER_5_31 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[22\] SUB SUB VPWR VPWR mask_rev_value\[22\]/HI mask_rev[22] sky130_fd_sc_hd__conb_1
XFILLER_2_32 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[15\] SUB SUB VPWR VPWR mask_rev_value\[15\]/HI mask_rev[15] sky130_fd_sc_hd__conb_1
XFILLER_2_44 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_32 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_11 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[9\] SUB SUB VPWR VPWR mask_rev_value\[9\]/HI mask_rev[9] sky130_fd_sc_hd__conb_1
XFILLER_8_44 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_23 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
Xmask_rev_value\[20\] SUB SUB VPWR VPWR mask_rev_value\[20\]/HI mask_rev[20] sky130_fd_sc_hd__conb_1
XPHY_10 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[13\] SUB SUB VPWR VPWR mask_rev_value\[13\]/HI mask_rev[13] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[7\] SUB SUB VPWR VPWR mask_rev_value\[7\]/HI mask_rev[7] sky130_fd_sc_hd__conb_1
XPHY_11 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XPHY_12 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
Xmask_rev_value\[29\] SUB SUB VPWR VPWR mask_rev_value\[29\]/HI mask_rev[29] sky130_fd_sc_hd__conb_1
XPHY_13 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[11\] SUB SUB VPWR VPWR mask_rev_value\[11\]/HI mask_rev[0] sky130_fd_sc_hd__conb_1
XPHY_14 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[5\] SUB SUB VPWR VPWR mask_rev_value\[5\]/HI mask_rev[5] sky130_fd_sc_hd__conb_1
XPHY_15 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
Xmask_rev_value\[27\] SUB SUB VPWR VPWR mask_rev_value\[27\]/HI mask_rev[27] sky130_fd_sc_hd__conb_1
XFILLER_6_40 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
XPHY_16 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_12
XPHY_17 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_42 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[3\] SUB SUB VPWR VPWR mask_rev_value\[3\]/HI mask_rev[3] sky130_fd_sc_hd__conb_1
XFILLER_6_32 SUB VPWR SUB VPWR sky130_fd_sc_hd__decap_4
Xmask_rev_value\[25\] SUB SUB VPWR VPWR mask_rev_value\[25\]/HI mask_rev[25] sky130_fd_sc_hd__conb_1
Xmask_rev_value\[18\] SUB SUB VPWR VPWR mask_rev_value\[18\]/HI mask_rev[18] sky130_fd_sc_hd__conb_1
.ends

.subckt sky130_fd_io__com_res_weak_v2 a_n281_1306# a_534_6146#
R0 a_n13_3671# m1_3_3617# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R1 a_n283_2797# a_n283_3382# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R2 a_n283_2797# m1_n268_3094# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R3 a_n281_1306# m1_n268_1364# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R4 a_n13_2329# m1_3_3580# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 a_n13_2329# a_n13_3671# sky130_fd_pr__res_generic_po w=0.8 l=6
R6 a_n283_2447# a_n283_2797# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R7 m1_n268_1924# a_n283_2447# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R8 m1_n268_2513# a_n283_2797# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R9 a_n283_3382# a_n13_2329# sky130_fd_pr__res_generic_po w=0.8 l=6
R10 m1_2_2233# a_n13_2329# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R11 a_n281_1656# m1_n268_1924# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R12 a_n13_6243# a_534_6146# sky130_fd_pr__res_generic_po w=0.8 l=50
R13 a_n13_3671# a_n13_6243# sky130_fd_pr__res_generic_po w=0.8 l=12
R14 a_n283_2447# m1_n268_2513# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R15 a_n283_3382# m1_2_2233# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R16 a_n281_1656# a_n283_2447# sky130_fd_pr__res_generic_po w=0.8 l=1.5
R17 m1_n268_3094# a_n283_3382# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R18 m1_n268_1364# a_n281_1656# sky130_fd_pr__res_generic_m1 w=0.66 l=10m
R19 a_n281_1306# a_n281_1656# sky130_fd_pr__res_generic_po w=0.8 l=1.5
.ends

.subckt sky130_fd_io__xres4v2_in_buf IN_H VNORMAL VNORMAL_B PAD ENABLE_HV IN_H_N ENABLE_VDDIO_LV
+ VDDIO a_n445_2580# m2_288_2575# w_4058_2188# a_n32352_n9635# VCCHIB VGND
Xsky130_fd_io__hvsbt_nand2_0 ENABLE_HV VNORMAL_B sky130_fd_io__hvsbt_nand2_0/OUT VGND
+ VDDIO VDDIO VGND sky130_fd_io__hvsbt_nand2
Xsky130_fd_io__inv_1_0 VCCHIB VGND sky130_fd_io__inv_1_0/Y ENABLE_VDDIO_LV VGND VCCHIB
+ sky130_fd_io__inv_1
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO VGND VDDIO sky130_fd_io__hvsbt_nand2_0/OUT
+ VGND sky130_fd_io__hvsbt_inv_x1
X0 a_n445_2580# sky130_fd_io__inv_1_0/Y VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X1 VDDIO VNORMAL a_157_2580# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X2 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X3 a_n29280_n8739# VNORMAL_B a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
X4 a_n11573_n8777# sky130_fd_io__hvsbt_inv_x1_0/OUT VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X5 VGND a_n176_869# a_2300_3398# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 a_1560_2580# ENABLE_HV VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X7 VGND IN_H_N IN_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.5
X8 VGND PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X9 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.8
X10 a_2165_2545# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X11 VGND a_2165_2545# a_2356_3115# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X12 VDDIO a_2356_3115# a_2300_3398# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.0588 pd=0.7 as=0.118 ps=1.4 w=0.42 l=0.5
X13 IN_H_N a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X14 a_n176_869# PAD w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.8
X15 a_n16_901# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.8
X16 a_1560_2580# ENABLE_HV VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.33 ps=10.5 w=5 l=0.5
X17 a_n232_901# PAD VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X18 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=0.5
X19 IN_H_N a_2300_3398# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.795 ps=6.53 w=3 l=0.5
X20 a_2356_3115# a_2165_2545# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X21 VDDIO sky130_fd_io__hvsbt_inv_x1_0/OUT a_n29280_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X22 a_n176_869# PAD a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.8
X23 a_n9813_4210# VNORMAL_B a_n11573_n8777# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X24 a_2300_3398# a_n176_869# VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X25 w_4058_2188# sky130_fd_io__hvsbt_inv_x1_0/OUT a_n445_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X26 VGND VGND VGND VGND sky130_fd_pr__nfet_05v0_nvt ad=8.81 pd=68.6 as=2.65 ps=20.5 w=10 l=0.9
X27 a_2165_2545# a_n176_869# w_4058_2188# w_4058_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.5
X28 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=0.5
X29 IN_H IN_H_N VGND VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.5
X30 a_469_2037# a_n176_869# a_n232_901# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X31 a_n31524_n8739# a_n29280_n8739# VGND sky130_fd_pr__res_generic_nd__hv w=0.29 l=1.08k
X32 VDDIO IN_H_N IN_H VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.42 ps=3.28 w=3 l=0.5
X33 a_n232_901# PAD a_n176_869# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X34 a_n757_2580# sky130_fd_io__hvsbt_inv_x1_0/OUT w_5030_2188# VGND sky130_fd_pr__nfet_05v0_nvt ad=2.8 pd=20.6 as=2.8 ps=20.6 w=10 l=0.9
X35 a_n16_901# VNORMAL_B VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X36 VCCHIB sky130_fd_io__inv_1_0/Y a_n757_2580# VCCHIB sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.4 ps=10.6 w=5 l=0.5
R0 a_n11573_n8777# a_n9813_4210# sky130_fd_pr__res_generic_po w=0.4 l=714
X37 w_5030_2188# w_5030_2188# w_5030_2188# w_5030_2188# sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=7.68 as=0.28 ps=2.56 w=1 l=0.8
X38 a_n232_901# a_n176_869# a_469_2037# VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.8
X39 a_n176_869# PAD a_n31524_n8739# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=1.4 ps=10.6 w=5 l=0.5
X40 a_2165_2545# a_n176_869# a_n9813_4210# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.4 pd=10.6 as=0.7 ps=5.28 w=5 l=0.5
X41 a_469_2037# PAD a_157_2580# VGND sky130_fd_pr__nfet_05v0_nvt ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.9
X42 IN_H IN_H_N VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.795 ps=6.53 w=3 l=0.5
X43 a_2356_3115# a_2300_3398# VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.0588 ps=0.7 w=0.42 l=0.5
.ends

.subckt sky130_fd_io__xres_inv_hysv2 OUT_H VSSD a_122_112# a_322_144# a_322_604# VCC_IO
X0 a_578_144# a_122_112# a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.42 ps=3.28 w=3 l=1
X1 a_322_144# OUT_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=1
X2 a_322_144# a_122_112# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=1
X3 a_578_144# a_122_112# a_322_144# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.14 ps=1.28 w=1 l=1
X4 OUT_H a_578_144# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X5 VCC_IO OUT_H a_322_604# VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.118 pd=1.4 as=0.118 ps=1.4 w=0.42 l=1
X6 OUT_H a_578_144# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.28 pd=2.56 as=0.28 ps=2.56 w=1 l=0.5
X7 a_322_604# a_122_112# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0.42 pd=3.28 as=0.84 ps=6.56 w=3 l=1
.ends

.subckt sky130_fd_io__gpio_buf_localesdv2 VTRIP_SEL_H OUT_H OUT_VT sky130_fd_io__res250only_small_0/PAD
+ VGND VCC_IO
Xsky130_fd_io__signal_5_sym_hv_local_5term_0 VGND VCC_IO OUT_VT VCC_IO VCC_IO VGND
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_1 VGND VCC_IO VGND OUT_VT VCC_IO VGND sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_2 VGND VCC_IO OUT_H VCC_IO VCC_IO VGND
+ sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__signal_5_sym_hv_local_5term_3 VGND VCC_IO VGND OUT_H VCC_IO VGND sky130_fd_io__signal_5_sym_hv_local_5term
Xsky130_fd_io__res250only_small_0 sky130_fd_io__res250only_small_0/PAD OUT_H sky130_fd_io__res250only_small
X0 OUT_VT VTRIP_SEL_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 ad=0.795 pd=6.53 as=0.795 ps=6.53 w=3 l=1
.ends

.subckt sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 VCC_IO a_10282_1285# a_5322_1285#
+ a_8980_1457# a_7988_1457# a_2036_1457# a_13940_1457# a_12948_1457# a_12266_1285#
+ a_7306_1285# a_5012_1457# a_3900_1285# a_2908_1285# a_5884_1285# a_14178_1285# a_10844_1285#
+ a_1354_1285# a_7868_1285# a_12828_1285# a_8860_1285# a_13820_1285# a_4330_1285#
+ a_3338_1285# a_6996_1457# a_11956_1457# a_1044_1457# a_11274_1285# a_6314_1285#
+ w_469_785# a_9972_1457# a_4020_1457# a_3028_1457# a_8298_1285# a_13258_1285# a_9290_1285#
+ a_1916_1285# a_6004_1457# a_4892_1285# a_6876_1285# a_924_1285# a_11836_1285# a_2346_1285#
+ a_9852_1285# a_10964_1457#
X0 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X1 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X3 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X4 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X7 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X8 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X10 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X11 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X12 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X13 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X16 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X19 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X20 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X21 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X22 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X23 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X26 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X27 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_469_785# a_11274_1285# a_10964_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 w_469_785# a_5322_1285# a_5012_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X30 a_9972_1457# a_9852_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X31 a_10964_1457# a_10844_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X32 w_469_785# a_2346_1285# a_2036_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_6996_1457# a_6876_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X34 w_469_785# a_6314_1285# a_6004_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X35 a_2036_1457# a_1916_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X36 w_469_785# a_12266_1285# a_11956_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X37 a_11956_1457# a_11836_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_5012_1457# a_4892_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_469_785# a_4330_1285# a_4020_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_469_785# a_9290_1285# a_8980_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_8980_1457# a_8860_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X42 w_469_785# a_10282_1285# a_9972_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X43 a_1044_1457# a_924_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.42 ps=11.4 w=5 l=0.6
X44 a_4020_1457# a_3900_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X45 w_469_785# a_3338_1285# a_3028_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X46 w_469_785# a_8298_1285# a_7988_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 a_3028_1457# a_2908_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X48 a_7988_1457# a_7868_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X49 w_469_785# a_13258_1285# a_12948_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X50 w_469_785# a_7306_1285# a_6996_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X51 a_13940_1457# a_13820_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X52 a_12948_1457# a_12828_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X53 w_469_785# a_1354_1285# a_1044_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 w_469_785# a_14178_1285# a_13940_1457# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.42 pd=11.4 as=2.97 ps=6.19 w=5 l=0.6
X55 a_6004_1457# a_5884_1285# w_469_785# w_469_785# sky130_fd_pr__nfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pddrvr_strong_xres4v2 PD_H[2] PD_H[3] TIE_LO_ESD VGND_IO
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457# m1_785_3898# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ VCC_IO
Xsky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0 VCC_IO PD_H[3] m1_9769_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_8980_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_7988_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_2036_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_13940_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_12948_1457#
+ m1_2697_3903# m1_7657_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_5012_1457#
+ m1_11193_3903# m1_11193_3903# m1_8232_3903# m1_785_3898# PD_H[3] m1_12747_3903#
+ PD_H[2] m1_2135_3903# PD_H[2] m1_785_3898# m1_9769_3903# m1_11193_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6996_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_11956_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_1044_1457#
+ PD_H[3] m1_8232_3903# w_335_3259# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_9972_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_4020_1457# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_3028_1457#
+ PD_H[2] m1_785_3898# PD_H[3] m1_12747_3903# sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_6004_1457#
+ m1_9769_3903# m1_8232_3903# m1_12747_3903# PD_H[3] m1_12747_3903# PD_H[3] sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2_0/a_10964_1457#
+ sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2
R0 PD_H[2] m2_6804_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 PD_H[2] m2_12763_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 m1_2135_3903# m2_1848_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R3 TIE_LO_ESD m2_13622_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_12747_3903# m2_12763_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 PD_H[2] m2_1260_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_7657_3903# m2_6804_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 PD_H[2] m2_897_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m2_13622_1100# m1_12747_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m2_1260_1100# m1_2135_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 m1_785_3898# m2_897_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 TIE_LO_ESD m2_12189_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 PD_H[2] m2_9986_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 TIE_LO_ESD m2_413_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 PD_H[3] m2_3095_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 TIE_LO_ESD m2_9366_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 m1_11193_3903# m2_12189_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 m1_9769_3903# m2_9986_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 m2_413_1100# m1_785_3898# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 m1_2697_3903# m2_3095_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m1_8232_3903# m2_9366_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 PD_H[3] m2_11758_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 m2_11758_1100# m1_11193_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 PD_H[3] m2_8935_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 TIE_LO_ESD m2_10846_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 PD_H[3] m2_656_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 PD_H[2] m2_11329_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 PD_H[3] m2_1565_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 TIE_LO_ESD m2_3378_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m2_8935_1100# m1_8232_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 m1_9769_3903# m2_10846_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R31 m1_11193_3903# m2_11329_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R32 PD_H[2] m2_8506_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R33 PD_H[3] m2_10415_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R34 m1_785_3898# m2_656_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R35 TIE_LO_ESD m2_7664_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R36 m1_2135_3903# m2_1565_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R37 m1_2697_3903# m2_3378_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R38 m1_8232_3903# m2_8506_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R39 m2_10415_1100# m1_9769_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R40 m1_7657_3903# m2_7664_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R41 PD_H[3] m2_7233_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R42 PD_H[3] m2_13193_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R43 PD_H[2] m2_2790_1100# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R44 m2_7233_1100# m1_7657_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R45 m1_12747_3903# m2_13193_1400# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R46 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po w=0.5 l=10.2
R47 TIE_LO_ESD m2_1848_1099# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R48 m2_2790_1100# m1_2697_3903# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__tk_tie_r_out_esd A B
R0 A B sky130_fd_pr__res_generic_po w=0.5 l=10.2
.ends

.subckt sky130_fd_io__xres2v2_rcfilter_lpfv2 IN a_9105_2295# a_1381_4189# a_7373_4189#
+ a_3949_4189# a_2237_4189# a_525_4189# a_472_471# a_7393_2295# a_472_1087# a_8249_2295#
+ a_5661_4189# a_472_779# a_336_26# a_472_317# a_472_1549# a_6517_4189# a_6537_2295#
+ a_9941_4189# a_472_163# a_3093_4189# a_472_1395# a_4805_4189# a_9961_2295# a_9085_4189#
+ VCC_IO a_472_1857#
X0 a_472_317# a_472_1087# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=25.3 pd=189 as=0.98 ps=7.28 w=7 l=4
X1 a_9941_4189# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R0 a_11618_2147# m1_14480_2172# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R1 a_11618_3071# m1_14484_3300# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R2 a_7373_4189# m1_14480_4922# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R3 IN m1_14484_4202# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R4 a_7373_4189# m1_11613_5471# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R5 m1_14328_5846# a_5661_4189# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X2 a_3382_6882# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X3 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R6 a_472_6420# m1_3338_6444# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R7 a_5661_4189# m1_14480_5846# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R8 m1_3363_1728# a_3382_1703# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R9 a_11618_3071# m1_14480_3096# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R10 a_7373_4189# m1_14484_5126# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R11 a_472_317# m1_3338_341# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R12 a_472_7344# m1_3338_7368# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R13 a_472_1395# m1_467_1384# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R14 a_472_779# m1_467_769# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X4 VCC_IO a_2237_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=25.3 pd=189 as=0.653 ps=4.85 w=6.12 l=4
X5 a_11618_3379# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R15 a_472_1087# m1_3334_1112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R16 a_472_1857# m1_5939_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R17 m1_3363_496# a_3382_471# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X6 a_472_7036# a_3382_7190# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X7 a_472_317# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R18 a_11618_2455# m1_14484_2684# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X8 a_9085_4189# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R19 a_472_1395# m1_10927_1419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X9 a_6517_4189# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R20 a_472_6728# m1_3338_6752# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X10 a_472_6728# a_472_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R21 a_7373_4189# m1_14484_5434# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R22 a_472_317# m1_5624_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X11 a_472_317# a_7393_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R23 a_472_7652# m1_3338_7676# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X12 a_11618_3687# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R24 a_472_317# m1_6480_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R25 m1_3363_1112# a_3382_1087# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X13 a_3382_7190# a_9085_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X14 a_472_317# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R26 a_11618_2763# m1_14484_2992# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R27 a_472_1395# m1_14299_5846# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R28 a_472_317# m1_467_432# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R29 a_472_317# m1_4825_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X15 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
R30 a_472_317# m1_6537_426# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R31 a_472_317# m1_4768_1042# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X16 a_472_6728# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X17 a_472_1549# a_3382_1703# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R32 a_6517_4189# m1_14484_5742# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X18 a_472_6112# a_472_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X19 a_7373_4189# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X20 a_472_317# a_8249_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R33 a_472_7036# m1_3338_7060# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X21 a_472_7036# a_472_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R34 a_472_471# m1_467_461# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R35 a_472_7344# m1_3338_7419# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X22 a_472_1087# a_3382_1087# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R36 a_472_1549# m1_2201_1652# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
R37 a_472_317# m1_3338_700# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X23 VCC_IO a_7373_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=6.12 l=4
X24 a_3382_1703# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R38 a_472_779# m1_10929_804# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X25 a_472_6420# a_472_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X26 a_472_6112# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X27 a_472_779# a_3382_779# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R39 a_7373_4189# m1_11741_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R40 a_472_6728# m1_3338_6803# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X28 a_472_7344# a_472_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X29 a_472_7036# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R41 a_472_7652# m1_3338_7727# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X30 a_472_1395# a_3382_1395# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R42 a_472_317# m1_2201_1681# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X31 a_472_317# a_472_779# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
X32 a_3382_1087# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R43 a_472_163# m1_10929_188# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X33 a_11618_2147# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R44 a_472_1549# m1_466_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X34 a_472_317# a_472_1857# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
X35 a_472_317# a_472_471# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R45 a_472_6112# m1_3338_6187# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R46 a_472_6728# m1_3334_6907# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X36 a_472_6420# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X37 a_472_7652# a_472_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X38 a_472_7344# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X39 a_472_163# a_3382_163# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X40 VCC_IO a_3949_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
X41 VCC_IO a_5661_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
X42 a_3382_1395# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R47 a_472_471# m1_10929_496# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X43 a_11618_2455# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R48 a_472_7036# m1_3338_7111# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X44 a_11618_3379# a_12884_625# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R49 a_472_6420# m1_3338_6495# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R50 a_472_317# m1_3338_392# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X45 a_7373_4189# a_12884_6728# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X46 a_472_317# a_6537_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R51 m1_3363_6907# a_3382_6882# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X47 a_472_7652# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X48 a_9085_4189# a_12884_7344# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R52 a_11618_2147# m1_14484_2325# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X49 a_472_471# a_3382_471# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R53 m1_10958_804# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R54 a_11618_3071# m1_14484_3249# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R55 a_472_7036# m1_3334_7215# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R56 a_472_317# m1_3338_1265# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X50 a_11618_2763# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R57 a_472_1395# m1_10927_1470# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X51 VCC_IO a_6517_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
R58 a_472_6420# m1_3334_6599# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X52 a_11618_3687# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R59 a_472_317# m1_3113_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R60 a_9941_4189# m1_14484_4459# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X53 a_3382_779# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X54 a_6517_4189# a_12884_6420# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R61 a_472_317# m1_3056_1350# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R62 m1_10958_188# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X55 a_7373_4189# a_12884_7036# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X56 a_472_317# a_9105_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R63 a_11618_2455# m1_14484_2633# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X57 a_472_317# a_472_1549# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.86 ps=14.5 w=7 l=4
R64 a_11618_3379# m1_14484_3557# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X58 a_472_317# a_472_1395# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R65 a_472_1549# m1_3338_1573# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X59 a_472_1549# a_472_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R66 a_472_7344# m1_3334_7523# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R67 a_5661_4189# m1_11613_5808# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R68 m1_3363_7215# a_3382_7190# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R69 m1_14509_2480# a_12884_1549# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R70 m1_3363_6599# a_3382_6574# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R71 a_472_1549# m1_10929_1728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R72 a_9085_4189# m1_14484_4767# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X60 VCC_IO a_3093_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
R73 m1_14509_4306# a_12884_7652# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R74 a_472_779# m1_3334_804# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R75 a_472_317# m1_3338_1008# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X61 VCC_IO a_525_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.928 ps=7.26 w=6.12 l=4
X62 a_5661_4189# a_12884_6112# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X63 a_11618_3071# a_12884_933# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R76 m1_10958_496# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R77 a_11618_2763# m1_14484_2941# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R78 a_9941_4189# m1_11613_4547# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R79 m1_14509_5230# a_12884_6728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X64 a_472_7652# a_3382_7806# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R80 a_472_1857# m1_1345_1960# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
X65 a_3382_163# a_11618_3687# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X66 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R81 a_472_1857# m1_3338_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R82 a_11618_3687# m1_14484_3865# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X67 a_472_1857# a_472_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X68 a_472_1549# a_12884_1549# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R83 a_472_7652# m1_3334_7831# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R84 m1_14509_3404# a_12884_625# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X69 a_9941_4189# a_12884_7652# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X70 a_11618_2455# a_11618_2455# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R85 m1_3363_7523# a_3382_7498# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R86 a_472_163# m1_3334_188# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R87 m1_14509_2788# a_12884_1241# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X71 a_472_6112# a_3382_6266# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R88 a_472_1549# m1_595_1664# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
X72 a_472_317# a_472_163# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
R89 m1_14509_4614# a_12884_7344# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R90 a_472_6112# m1_3334_6291# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R91 a_472_317# m1_3338_1316# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R92 m1_10958_1728# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R93 a_9085_4189# m1_11613_4576# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R94 a_472_317# m1_1345_1989# sky130_fd_pr__res_generic_m1 w=0.29 l=10m
R95 a_472_1087# m1_10929_1112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R96 IN m1_14484_4151# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R97 a_9085_4189# m1_11613_4855# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R98 m1_14509_5538# a_12884_6420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X73 a_3382_7806# IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X74 a_3382_471# a_11618_3379# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R99 a_11618_2455# m1_14480_2480# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R100 a_9941_4189# m1_14484_4510# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R101 a_7373_4189# m1_14484_5075# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R102 a_6517_4189# m1_11613_5779# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X75 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X76 a_472_1857# a_12884_1857# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R103 m1_14509_3712# a_12884_317# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R104 a_472_317# m1_3338_649# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X77 VCC_IO a_4805_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
X78 a_11618_2763# a_11618_2763# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R105 m1_3363_7831# a_3382_7806# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R106 a_9941_4189# m1_14480_4306# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R107 a_472_1857# m1_5939_1881# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R108 a_472_471# m1_3334_496# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X79 a_472_6420# a_3382_6574# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X80 a_3382_6266# a_6517_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X81 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R109 a_472_1395# m1_3334_1420# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R110 a_7373_4189# m1_14480_5230# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R111 a_11618_3379# m1_14484_3608# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R112 a_6517_4189# m1_11613_5500# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
X82 a_472_7344# a_3382_7498# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R113 a_472_1549# m1_3338_1624# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R114 m1_14509_2172# a_12884_1857# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R115 m1_14509_4922# a_12884_7036# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R116 a_472_317# m1_467_1047# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R117 a_7373_4189# m1_11613_4884# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R118 a_472_317# m1_5681_734# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R119 m1_3363_6291# a_3382_6266# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R120 a_11618_3379# m1_14480_3404# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R121 m1_14509_5846# a_12884_6112# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R122 m1_14509_3096# a_12884_933# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R123 m1_10958_1112# a_472_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R124 a_11618_2763# m1_14480_2788# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R125 a_9085_4189# m1_14484_4818# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X83 a_472_317# a_9961_2295# a_472_317# a_336_26# sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.98 ps=7.28 w=7 l=4
X84 a_472_317# a_472_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R126 a_7373_4189# m1_14484_5383# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R127 a_472_317# m1_3338_957# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X85 IN IN a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R128 a_9085_4189# m1_14480_4614# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R129 m1_3363_804# a_3382_779# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X86 VCC_IO a_9085_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
X87 a_472_6728# a_3382_6882# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
X88 a_3382_6574# a_7373_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R130 a_472_1549# m1_3334_1728# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X89 a_472_317# a_12884_1241# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R131 a_472_6112# m1_3338_6136# sky130_fd_pr__res_generic_m1 w=0.29 l=0.31
R132 a_6517_4189# m1_14480_5538# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X90 VCC_IO a_1381_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
X91 a_11618_2147# a_11618_2147# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R133 a_472_1857# m1_3338_1932# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R134 m1_3363_1420# a_3382_1395# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R135 a_472_1087# m1_467_1076# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R136 a_11618_3687# m1_14484_3916# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X92 a_3382_7498# a_9941_4189# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
X93 VCC_IO a_9941_4189# VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.653 ps=4.85 w=6.12 l=4
R137 a_472_317# m1_467_1355# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R138 a_7373_4189# m1_11612_5169# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
X94 a_11618_3071# a_11618_3071# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=14
R139 a_11618_3687# m1_14480_3712# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
R140 a_472_317# m1_467_740# sky130_fd_pr__res_generic_m1 w=0.65 l=10m
R141 m1_3363_188# a_3382_163# sky130_fd_pr__res_generic_m1 w=0.26 l=10m
X95 a_472_317# a_12884_317# a_336_26# sky130_fd_pr__res_generic_nd w=0.5 l=47
R142 a_11618_2147# m1_14484_2376# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
R143 a_6517_4189# m1_14484_5691# sky130_fd_pr__res_generic_m1 w=0.26 l=0.31
.ends

.subckt sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2 w_415_600# a_4969_1552# a_2303_1380#
+ a_5961_1552# a_13777_1380# a_8817_1380# a_4287_1380# a_10921_1552# a_7945_1552#
+ a_12905_1552# a_7263_1380# a_12223_1380# a_9929_1552# a_9247_1380# a_2865_1380#
+ a_1993_1552# a_5841_1380# a_4849_1380# a_10801_1380# a_14135_1380# a_1311_1380#
+ a_3977_1552# a_12785_1380# a_7825_1380# a_3295_1380# a_6953_1552# a_9809_1380# a_11913_1552#
+ a_1001_1552# a_6271_1380# a_5279_1380# a_11231_1380# a_10239_1380# a_13897_1552#
+ a_8937_1552# a_8255_1380# a_1873_1380# a_13215_1380# a_3857_1380# a_2985_1552# a_11793_1380#
+ a_881_1380# a_6833_1380#
X0 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X1 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X2 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X3 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X4 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X5 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X6 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X7 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X8 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X9 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X10 a_4969_1552# a_4849_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X11 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X12 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X13 w_415_600# a_10239_1380# a_9929_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X14 a_8937_1552# a_8817_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X15 w_415_600# a_3295_1380# a_2985_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X16 w_415_600# a_2303_1380# a_1993_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X17 w_415_600# a_7263_1380# a_6953_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X18 a_12905_1552# a_12785_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X19 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X20 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X21 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X22 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X23 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X24 a_3977_1552# a_3857_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X25 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X26 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X27 a_7945_1552# a_7825_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X28 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X29 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X30 w_415_600# a_13215_1380# a_12905_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X31 w_415_600# a_1311_1380# a_1001_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X32 w_415_600# a_6271_1380# a_5961_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X33 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X34 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X35 w_415_600# a_5279_1380# a_4969_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X36 a_11913_1552# a_11793_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X37 a_10921_1552# a_10801_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X38 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X39 w_415_600# a_9247_1380# a_8937_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X40 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X41 a_1001_1552# a_881_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=4.32 ps=11.7 w=5 l=0.6
X42 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X43 a_2985_1552# a_2865_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X44 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X45 a_6953_1552# a_6833_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X46 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X47 w_415_600# a_12223_1380# a_11913_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X48 a_13897_1552# a_13777_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=2.97 pd=6.19 as=3.78 ps=11.5 w=5 l=0.6
X49 a_9929_1552# a_9809_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X50 a_1993_1552# a_1873_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X51 w_415_600# a_4287_1380# a_3977_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X52 w_415_600# a_14135_1380# a_13897_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=4.3 pd=11.7 as=2.97 ps=6.19 w=5 l=0.6
X53 w_415_600# a_8255_1380# a_7945_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
X54 a_5961_1552# a_5841_1380# w_415_600# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.88 pd=6.55 as=3.78 ps=11.5 w=5 l=0.6
X55 w_415_600# a_11231_1380# a_10921_1552# w_415_600# sky130_fd_pr__pfet_g5v0d10v5 ad=3.78 pd=11.5 as=3.88 ps=6.55 w=5 l=0.6
.ends

.subckt sky130_fd_io__gpio_pudrvr_strong_axres4v2 PU_H_N[3] PU_H_N[2] TIE_HI_ESD sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ VNB sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552# li_11868_461#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ a_14575_48# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
Xsky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0 sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/w_415_600#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_4969_1552# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_5961_1552#
+ m1_14229_1478# m1_8837_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_10921_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_7945_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_12905_1552#
+ PU_H_N[3] m1_11745_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_9929_1552#
+ m1_8837_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1993_1552#
+ PU_H_N[3] PU_H_N[3] m1_10391_1478# m1_14229_1478# PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_3977_1552#
+ PU_H_N[2] PU_H_N[3] PU_H_N[2] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_6953_1552#
+ m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_11913_1552# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_1001_1552#
+ PU_H_N[3] PU_H_N[3] m1_11745_1478# m1_10391_1478# sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_13897_1552#
+ sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_8937_1552# m1_8837_1478# PU_H_N[2]
+ m1_13667_1478# PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0/a_2985_1552#
+ m1_11745_1478# PU_H_N[2] PU_H_N[3] sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2
R0 m1_14229_1478# m2_14532_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R1 m1_13667_1478# m2_13593_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R2 TIE_HI_ESD a_14575_48# sky130_fd_pr__res_generic_po w=0.5 l=10.2
R3 PU_H_N[2] m2_9839_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R4 m1_10391_1478# m2_10945_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R5 PU_H_N[2] m2_11422_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R6 m1_13667_1478# m2_14075_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R7 m2_12267_n279# m1_11745_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R8 m1_11745_1478# m2_12510_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R9 m1_8837_1478# m2_9605_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R10 TIE_HI_ESD m2_10945_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R11 m1_8837_1478# m2_9363_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R12 m1_10391_1478# m2_11422_92# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R13 PU_H_N[3] m2_9605_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R14 PU_H_N[3] m2_12510_n280# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R15 PU_H_N[2] m2_14769_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R16 PU_H_N[3] m2_11186_n208# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R17 PU_H_N[3] m2_13837_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R18 TIE_HI_ESD m2_14286_658# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R19 PU_H_N[3] m2_14532_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R20 m2_11186_n208# m1_10391_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R21 TIE_HI_ESD m2_13593_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R22 PU_H_N[2] m2_12751_n280# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R23 m2_13837_658# m1_13667_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R24 m1_14229_1478# m2_14769_958# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R25 m1_11745_1478# m2_12751_21# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R26 TIE_HI_ESD m2_9363_n209# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R27 TIE_HI_ESD m2_12267_n279# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R28 m2_9839_n208# m1_8837_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R29 m2_14286_658# m1_14229_1478# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
R30 PU_H_N[2] m2_14075_657# sky130_fd_pr__res_generic_m2 w=0.65 l=10m
.ends

.subckt sky130_fd_io__top_xres4v2 XRES_H_N FILT_IN_H ENABLE_VDDIO TIE_WEAK_HI_H ENABLE_H
+ PULLUP_H EN_VDDIO_SIG_H TIE_LO_ESD TIE_HI_ESD DISABLE_PULLUP_H INP_SEL_H VSSA AMUXBUS_B
+ AMUXBUS_A VDDIO_Q VSWITCH VDDA VCCD VCCHIB VSSIO_Q VDDIO VSSD VSSIO PAD PAD_A_ESD_H
Xsky130_fd_io__com_res_weak_v2_0 PULLUP_H a_5670_7125# sky130_fd_io__com_res_weak_v2
Xsky130_fd_io__com_res_weak_0 sky130_fd_io__com_res_weak_0/RB VDDIO li_7794_26629#
+ li_9658_25954# li_12154_26629# li_8568_25954# li_11000_25954# sky130_fd_io__com_res_weak
Xsky130_fd_io__hvsbt_inv_x4_1 sky130_fd_io__hvsbt_inv_x4_1/IN XRES_H_N VDDIO_Q VSSD
+ VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__hvsbt_inv_x4_0 sky130_fd_io__hvsbt_inv_x4_1/IN XRES_H_N VDDIO_Q VSSD
+ VSSD VDDIO_Q sky130_fd_io__hvsbt_inv_x4
Xsky130_fd_io__xres4v2_in_buf_0 sky130_fd_io__xres4v2_in_buf_0/IN_H EN_VDDIO_SIG_H
+ sky130_fd_io__hvsbt_inv_x2_0/OUT sky130_fd_io__xres4v2_in_buf_0/PAD ENABLE_H sky130_fd_io__xres4v2_in_buf_0/IN_H_N
+ ENABLE_VDDIO VDDIO_Q m1_3250_3609# EN_VDDIO_SIG_H m1_1351_2970# VSSD VCCHIB VSSD
+ sky130_fd_io__xres4v2_in_buf
Xsky130_fd_io__hvsbt_inv_x2_0 VDDIO_Q VSSD EN_VDDIO_SIG_H sky130_fd_io__hvsbt_inv_x2_0/OUT
+ VDDIO_Q VSSD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_inv_x2_1 VDDIO VSSD sky130_fd_io__hvsbt_inv_x2_1/IN sky130_fd_io__hvsbt_inv_x2_1/OUT
+ VDDIO VSSD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_inv_x2_2 VDDIO VSSD DISABLE_PULLUP_H sky130_fd_io__hvsbt_inv_x2_1/IN
+ VDDIO VSSD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__hvsbt_inv_x2_3 VDDIO_Q VSSD INP_SEL_H sky130_fd_io__hvsbt_inv_x2_3/OUT
+ VDDIO_Q VSSD sky130_fd_io__hvsbt_inv_x2
Xsky130_fd_io__xres_inv_hysv2_0 sky130_fd_io__xres_inv_hysv2_0/OUT_H VSSD m1_6377_8979#
+ li_6043_2944# li_5552_2976# VDDIO_Q sky130_fd_io__xres_inv_hysv2
Xsky130_fd_io__gpio_buf_localesdv2_0 VSSD sky130_fd_io__xres4v2_in_buf_0/PAD sky130_fd_io__gpio_buf_localesdv2_0/OUT_VT
+ PAD VSSD VDDIO sky130_fd_io__gpio_buf_localesdv2
Xsky130_fd_io__gpio_pddrvr_strong_xres4v2_0 sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3] sky130_fd_io__gpio_pddrvr_strong_xres4v2_0/PD_H[3]
+ VSSIO PAD PAD PAD PAD PAD PAD PAD PAD VSSIO PAD PAD PAD PAD PAD m1_915_33059# PAD
+ VDDIO sky130_fd_io__gpio_pddrvr_strong_xres4v2
Xsky130_fd_io__tk_tie_r_out_esd_0 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__tk_tie_r_out_esd_1 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
Xsky130_fd_io__res250only_small_0 TIE_WEAK_HI_H sky130_fd_io__com_res_weak_0/RB sky130_fd_io__res250only_small
Xsky130_fd_io__hvsbt_inv_x1_0 sky130_fd_io__hvsbt_inv_x4_1/IN VDDIO_Q VSSD VDDIO_Q
+ sky130_fd_io__xres_inv_hysv2_0/OUT_H VSSD sky130_fd_io__hvsbt_inv_x1
Xsky130_fd_io__res250only_small_1 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
Xsky130_fd_io__xres2v2_rcfilter_lpfv2_0 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN
+ m1_10468_10072# m1_6377_8979# m1_10468_9216# m1_10468_4936# m1_10468_3224# m1_10468_1512#
+ m1_10468_4936# m1_10468_9216# m1_10468_3224# m1_10468_9216# m1_10468_6648# m1_10468_4080#
+ VSSD VSSD m1_10468_1512# m1_10468_7504# m1_10468_7504# m1_10468_10928# m1_10468_5792#
+ m1_10468_4080# m1_6377_8979# m1_10468_5792# m1_10468_10928# m1_10468_10072# VDDIO_Q
+ m1_10468_6648# sky130_fd_io__xres2v2_rcfilter_lpfv2
Xsky130_fd_io__gpio_pudrvr_strong_axres4v2_0 sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3] sky130_fd_io__gpio_pudrvr_strong_axres4v2_0/PU_H_N[3]
+ PAD PAD PAD PAD PAD PAD PAD PAD PAD VSSD PAD VSSD PAD PAD VDDIO PAD VDDIO PAD sky130_fd_io__gpio_pudrvr_strong_axres4v2
X0 a_5670_7125# sky130_fd_io__hvsbt_inv_x2_1/OUT VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=1.33 ps=10.5 w=5 l=0.5
X1 FILT_IN_H sky130_fd_io__hvsbt_inv_x2_3/OUT sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X2 VDDIO sky130_fd_io__hvsbt_inv_x2_1/OUT a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=1.33 pd=10.5 as=0.7 ps=5.28 w=5 l=0.5
X3 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN sky130_fd_io__hvsbt_inv_x2_3/OUT sky130_fd_io__xres4v2_in_buf_0/IN_H VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X4 VDDIO sky130_fd_io__hvsbt_inv_x2_1/OUT a_5670_7125# VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X5 a_5670_7125# sky130_fd_io__hvsbt_inv_x2_1/OUT VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 ad=0.7 pd=5.28 as=0.7 ps=5.28 w=5 l=0.5
X6 FILT_IN_H INP_SEL_H sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
X7 sky130_fd_io__xres2v2_rcfilter_lpfv2_0/IN INP_SEL_H sky130_fd_io__xres4v2_in_buf_0/IN_H VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 ad=0.84 pd=6.56 as=0.84 ps=6.56 w=3 l=0.5
.ends

.subckt chip_io_openframe vddio vssio_pad vdda_pad vccd2 vccd vdda vdda1 vdda2 vccd1
+ resetb_pad porb_h porb_l por_l resetb_h resetb_l mask_rev[31] mask_rev[30] mask_rev[29]
+ mask_rev[28] mask_rev[27] mask_rev[26] mask_rev[25] mask_rev[24] mask_rev[23] mask_rev[22]
+ mask_rev[21] mask_rev[20] mask_rev[19] mask_rev[18] mask_rev[17] mask_rev[16] mask_rev[15]
+ mask_rev[14] mask_rev[13] mask_rev[12] mask_rev[11] mask_rev[10] mask_rev[9] mask_rev[8]
+ mask_rev[7] mask_rev[6] mask_rev[5] mask_rev[4] mask_rev[3] mask_rev[2] mask_rev[1]
+ mask_rev[0] gpio[39] gpio[32] gpio[19] gpio_out[43] gpio_out[40] gpio_out[39] gpio_out[38]
+ gpio_out[37] gpio_out[36] gpio_out[28] gpio_out[27] gpio_out[26] gpio_out[25] gpio_out[19]
+ gpio_out[18] gpio_out[17] gpio_out[16] gpio_out[15] gpio_out[14] gpio_out[13] gpio_out[12]
+ gpio_out[11] gpio_out[10] gpio_out[0] gpio_oeb[43] gpio_oeb[42] gpio_oeb[41] gpio_oeb[40]
+ gpio_oeb[39] gpio_oeb[34] gpio_oeb[33] gpio_oeb[29] gpio_oeb[28] gpio_oeb[27] gpio_oeb[26]
+ gpio_oeb[25] gpio_oeb[23] gpio_oeb[22] gpio_oeb[21] gpio_oeb[20] gpio_oeb[17] gpio_oeb[16]
+ gpio_oeb[11] gpio_oeb[7] gpio_oeb[6] gpio_oeb[1] gpio_inp_dis[39] gpio_inp_dis[37]
+ gpio_inp_dis[35] gpio_inp_dis[34] gpio_inp_dis[33] gpio_inp_dis[30] gpio_inp_dis[29]
+ gpio_inp_dis[22] gpio_inp_dis[21] gpio_inp_dis[20] gpio_inp_dis[18] gpio_inp_dis[17]
+ gpio_inp_dis[16] gpio_inp_dis[13] gpio_inp_dis[12] gpio_inp_dis[9] gpio_inp_dis[5]
+ gpio_inp_dis[1] gpio_ib_mode_sel[43] gpio_ib_mode_sel[42] gpio_ib_mode_sel[41] gpio_ib_mode_sel[40]
+ gpio_ib_mode_sel[39] gpio_ib_mode_sel[38] gpio_ib_mode_sel[37] gpio_ib_mode_sel[34]
+ gpio_ib_mode_sel[32] gpio_ib_mode_sel[31] gpio_ib_mode_sel[26] gpio_ib_mode_sel[25]
+ gpio_ib_mode_sel[24] gpio_ib_mode_sel[23] gpio_ib_mode_sel[22] gpio_ib_mode_sel[21]
+ gpio_ib_mode_sel[20] gpio_ib_mode_sel[16] gpio_ib_mode_sel[13] gpio_ib_mode_sel[10]
+ gpio_ib_mode_sel[9] gpio_ib_mode_sel[7] gpio_ib_mode_sel[4] gpio_ib_mode_sel[1]
+ gpio_vtrip_sel[43] gpio_vtrip_sel[42] gpio_vtrip_sel[37] gpio_vtrip_sel[36] gpio_vtrip_sel[35]
+ gpio_vtrip_sel[28] gpio_vtrip_sel[27] gpio_vtrip_sel[26] gpio_vtrip_sel[25] gpio_vtrip_sel[24]
+ gpio_vtrip_sel[23] gpio_vtrip_sel[22] gpio_vtrip_sel[19] gpio_vtrip_sel[18] gpio_vtrip_sel[17]
+ gpio_vtrip_sel[16] gpio_vtrip_sel[15] gpio_vtrip_sel[14] gpio_vtrip_sel[13] gpio_vtrip_sel[12]
+ gpio_vtrip_sel[11] gpio_vtrip_sel[10] gpio_vtrip_sel[5] gpio_vtrip_sel[4] gpio_vtrip_sel[3]
+ gpio_vtrip_sel[2] gpio_vtrip_sel[1] gpio_vtrip_sel[0] gpio_slow_sel[43] gpio_slow_sel[34]
+ gpio_slow_sel[32] gpio_slow_sel[31] gpio_slow_sel[30] gpio_slow_sel[28] gpio_slow_sel[27]
+ gpio_slow_sel[26] gpio_slow_sel[22] gpio_slow_sel[21] gpio_slow_sel[17] gpio_slow_sel[15]
+ gpio_slow_sel[14] gpio_slow_sel[13] gpio_slow_sel[12] gpio_slow_sel[10] gpio_slow_sel[9]
+ gpio_slow_sel[8] gpio_slow_sel[5] gpio_slow_sel[4] gpio_slow_sel[0] gpio_holdover[42]
+ gpio_holdover[41] gpio_holdover[37] gpio_holdover[32] gpio_holdover[31] gpio_holdover[30]
+ gpio_holdover[29] gpio_holdover[26] gpio_holdover[25] gpio_holdover[22] gpio_holdover[21]
+ gpio_holdover[15] gpio_holdover[14] gpio_holdover[13] gpio_holdover[12] gpio_holdover[11]
+ gpio_holdover[10] gpio_holdover[9] gpio_holdover[8] gpio_holdover[7] gpio_holdover[6]
+ gpio_holdover[5] gpio_holdover[3] gpio_holdover[2] gpio_holdover[1] gpio_analog_en[41]
+ gpio_analog_en[40] gpio_analog_en[38] gpio_analog_en[37] gpio_analog_en[36] gpio_analog_en[35]
+ gpio_analog_en[34] gpio_analog_en[33] gpio_analog_en[32] gpio_analog_en[31] gpio_analog_en[30]
+ gpio_analog_en[29] gpio_analog_en[19] gpio_analog_en[18] gpio_analog_en[17] gpio_analog_en[16]
+ gpio_analog_en[8] gpio_analog_en[7] gpio_analog_en[6] gpio_analog_en[5] gpio_analog_en[4]
+ gpio_analog_en[3] gpio_analog_en[2] gpio_analog_en[1] gpio_analog_en[0] gpio_analog_sel[39]
+ gpio_analog_sel[38] gpio_analog_sel[36] gpio_analog_sel[35] gpio_analog_sel[34]
+ gpio_analog_sel[31] gpio_analog_sel[30] gpio_analog_sel[26] gpio_analog_sel[19]
+ gpio_analog_sel[18] gpio_analog_sel[16] gpio_analog_sel[15] gpio_analog_sel[14]
+ gpio_analog_sel[11] gpio_analog_sel[10] gpio_analog_sel[9] gpio_analog_sel[8] gpio_analog_sel[5]
+ gpio_analog_sel[4] gpio_analog_sel[0] gpio_analog_pol[43] gpio_analog_pol[39] gpio_analog_pol[38]
+ gpio_analog_pol[37] gpio_analog_pol[34] gpio_analog_pol[33] gpio_analog_pol[32]
+ gpio_analog_pol[29] gpio_analog_pol[25] gpio_analog_pol[19] gpio_analog_pol[18]
+ gpio_analog_pol[17] gpio_analog_pol[14] gpio_analog_pol[13] gpio_analog_pol[8] gpio_analog_pol[7]
+ gpio_analog_pol[6] gpio_analog_pol[3] gpio_analog_pol[2] gpio_dm0[39] gpio_dm0[30]
+ gpio_dm0[28] gpio_dm0[27] gpio_dm0[24] gpio_dm0[23] gpio_dm0[20] gpio_dm0[19] gpio_dm0[13]
+ gpio_dm0[12] gpio_dm0[11] gpio_dm0[10] gpio_dm0[8] gpio_dm0[7] gpio_dm0[3] gpio_dm1[41]
+ gpio_dm1[40] gpio_dm1[39] gpio_dm1[34] gpio_dm1[30] gpio_dm1[29] gpio_dm1[28] gpio_dm1[27]
+ gpio_dm1[26] gpio_dm1[25] gpio_dm1[24] gpio_dm1[23] gpio_dm1[21] gpio_dm1[20] gpio_dm1[19]
+ gpio_dm1[16] gpio_dm1[15] gpio_dm1[11] gpio_dm1[2] gpio_dm1[1] gpio_dm1[0] gpio_dm2[39]
+ gpio_dm2[37] gpio_dm2[35] gpio_dm2[34] gpio_dm2[31] gpio_dm2[30] gpio_dm2[27] gpio_dm2[23]
+ gpio_dm2[19] gpio_dm2[17] gpio_dm2[16] gpio_dm2[15] gpio_dm2[12] gpio_dm2[11] gpio_dm2[9]
+ gpio_dm2[8] gpio_dm2[7] gpio_dm2[6] gpio_dm2[4] gpio_dm2[3] gpio_dm2[0] gpio_in[39]
+ gpio_in[38] gpio_in[37] gpio_in[35] gpio_in[34] gpio_in[33] gpio_in[32] gpio_in[31]
+ gpio_in[30] gpio_in[27] gpio_in[26] gpio_in[23] gpio_in[18] gpio_in[17] gpio_in[16]
+ gpio_in[15] gpio_in[14] gpio_in[12] gpio_in[11] gpio_in[8] gpio_in[5] gpio_in_h[42]
+ gpio_in_h[39] gpio_in_h[37] gpio_in_h[34] gpio_in_h[33] gpio_in_h[32] gpio_in_h[29]
+ gpio_in_h[24] gpio_in_h[20] gpio_in_h[17] gpio_in_h[16] gpio_in_h[15] gpio_in_h[12]
+ gpio_in_h[11] gpio_in_h[10] gpio_in_h[7] gpio_in_h[6] gpio_in_h[2] gpio_in_h[1]
+ gpio_loopback_zero[43] gpio_loopback_zero[42] gpio_loopback_zero[41] gpio_loopback_zero[40]
+ gpio_loopback_zero[39] gpio_loopback_zero[38] gpio_loopback_one[43] gpio_loopback_one[42]
+ gpio_loopback_one[41] gpio_loopback_one[40] gpio_loopback_one[39] gpio_loopback_one[35]
+ gpio_loopback_one[31] gpio_loopback_one[29] gpio_loopback_one[28] gpio_loopback_one[27]
+ gpio_loopback_one[25] gpio_loopback_one[24] gpio_loopback_one[23] gpio_loopback_one[21]
+ gpio_loopback_one[20] gpio_loopback_one[17] gpio_loopback_one[13] gpio_loopback_one[9]
+ gpio_loopback_one[6] analog_io[43] analog_io[41] analog_io[39] analog_io[38] analog_io[35]
+ analog_io[34] analog_io[33] analog_io[30] analog_io[24] analog_io[20] analog_io[19]
+ analog_io[18] analog_io[16] analog_io[15] analog_io[14] analog_io[10] analog_io[9]
+ analog_io[8] analog_io[3] gpio[42] gpio[28] gpio[27] gpio[26] gpio[25] gpio[23]
+ gpio[1] gpio[0] gpio_analog_pol[20] w_694469_865869# w_23367_407274# w_694469_100152#
+ w_23367_534874# w_137274_1012253# gpio_out[1] w_188674_1014469# gpio_dm0[15] w_404752_21253#
+ w_459552_23367# w_485565_1014469# w_291674_1014469# w_638765_1014469# w_23367_280765#
+ gpio_out[2] w_692253_776670# w_23367_710765# gpio_holdover[16] gpio_inp_dis[25]
+ w_692355_547952# w_23367_537965# w_21151_364074# gpio_holdover[33] w_21253_966965#
+ gpio_out[3] w_694469_145352# w_459552_21253# w_692355_593152# w_485565_1012355#
+ w_694469_951752# w_694469_190352# w_638765_1012355# gpio_analog_pol[41] w_349952_23367#
+ gpio_analog_sel[40] gpio_out[4] w_692355_325552# w_189869_23367# gpio_inp_dis[41]
+ w_21151_794074# w_694469_235552# w_692355_683352# gpio_analog_sel[21] w_21253_194365#
+ w_694469_280552# w_85874_1014469# gpio_out[5] gpio_in_h[40] analog_io[40] gpio_loopback_one[2]
+ gpio_inp_dis[42] gpio_dm0[34] w_21253_624365# w_482474_1012253# w_295152_23367#
+ w_635674_1012253# w_349952_21253# gpio_in[20] gpio_analog_pol[24] w_23367_578074#
+ w_692253_551270# gpio_dm1[3] gpio_out[6] w_694469_370752# w_189869_21253# gpio_dm1[7]
+ gpio_in_h[23] gpio_in[2] gpio_out[7] gpio_oeb[0] gpio_slow_sel[37] w_21151_277674#
+ w_692253_641470# w_692253_955070# analog_io[23] w_295152_21253# w_294765_1014469#
+ gpio_inp_dis[6] gpio_analog_en[9] w_21151_707674# w_23367_234474# w_692355_100152#
+ w_694469_776669# gpio_analog_en[20] gpio_out[8] w_393474_1014469# w_21151_963874#
+ gpio_ib_mode_sel[29] gpio_holdover[39] gpio_inp_dis[2] gpio_dm0[16] w_692253_596470#
+ gpio_oeb[10] gpio_ib_mode_sel[28] gpio_dm1[12] gpio_analog_en[21] w_692253_731670#
+ w_21253_280765# analog_io[28] gpio_out[9] analog_io[29] w_692253_328870# gpio_holdover[17]
+ gpio_analog_en[22] w_23367_410365# w_21253_710765# gpio_loopback_one[10] gpio_inp_dis[26]
+ w_294765_1012355# gpio_holdover[34] w_462869_23367# w_23367_237565# gpio_in_h[28]
+ w_21253_537965# gpio_dm2[20] w_23367_664474# w_692253_686670# gpio_analog_en[23]
+ w_21151_191274# analog_io[2] gpio_in_h[0] gpio_analog_sel[25] w_692253_374070# gpio_oeb[5]
+ gpio_ib_mode_sel[11] gpio_dm2[24] w_21151_621274# w_692355_145352# gpio_analog_en[24]
+ gpio_analog_sel[20] gpio_out[41] w_692355_951752# w_692355_190352# w_694469_862552#
+ gpio_oeb[32] w_88965_1014469# gpio_analog_pol[28] gpio_loopback_one[14] gpio_dm2[28]
+ gpio_analog_pol[42] gpio_analog_en[25] w_188674_1012253# analog_io[7] gpio_analog_pol[23]
+ gpio_in[9] w_291674_1012253# gpio_oeb[15] w_462869_21253# w_23367_667565# gpio_in_h[22]
+ gpio_dm0[0] w_692355_235552# gpio_analog_en[26] w_694469_551269# gpio_dm0[31] gpio_vtrip_sel[39]
+ w_23367_320874# gpio_loopback_one[32] w_692355_280552# gpio_slow_sel[20] gpio_slow_sel[36]
+ gpio_in[24] gpio_slow_sel[38] gpio_dm0[4] gpio_analog_en[27] gpio_dm0[35] gpio_analog_en[42]
+ gpio_dm1[31] gpio_analog_sel[43] gpio_loopback_one[3] gpio_analog_sel[3] gpio_loopback_one[18]
+ analog_io[22] w_88965_1012355# gpio_ib_mode_sel[2] gpio_slow_sel[41] w_692253_103470#
+ gpio_in_h[5] w_140365_1014469# gpio_analog_en[28] w_694469_641469# w_694469_955069#
+ gpio_dm1[4] gpio_dm1[35] gpio_ib_mode_sel[14] w_692355_370752# gpio_slow_sel[3]
+ gpio_in[6] gpio_analog_sel[41] gpio_loopback_one[36] w_23367_323965# w_23367_750874#
+ gpio_vtrip_sel[38] gpio_dm1[8] gpio_oeb[37] w_396565_1014469# gpio_analog_pol[1]
+ w_240074_1014469# analog_io[27] gpio_analog_en[43] w_694469_596469# gpio_ib_mode_sel[35]
+ gpio_inp_dis[7] w_23367_581165# gpio_loopback_one[7] gpio_in[21] w_694469_731669#
+ gpio_analog_pol[12] w_21151_407274# w_186552_23367# gpio_in_h[27] w_517669_23367#
+ w_21151_534874# w_85874_1012253# w_694469_328869# w_140365_1012355# gpio_slow_sel[25]
+ gpio_oeb[4] gpio_inp_dis[3] gpio_analog_sel[29] analog_io[1] gpio_dm0[21] w_692253_148670#
+ w_23367_753965# gpio_in[3] w_694469_686669# gpio_dm0[17] w_692253_193670# gpio_analog_sel[24]
+ gpio_inp_dis[14] gpio_dm1[13] analog_io[13] gpio_in_h[43] gpio_oeb[31] w_694469_374069#
+ gpio_ib_mode_sel[5] gpio_dm0[25] gpio_holdover[18] w_396565_1012355# gpio_inp_dis[31]
+ gpio_inp_dis[27] gpio_ib_mode_sel[17] w_21253_410365# gpio_holdover[35] gpio_dm1[17]
+ w_694469_638152# gpio_inp_dis[10] gpio_dm2[13] gpio_oeb[14] analog_io[6] gpio_analog_pol[27]
+ gpio_in_h[21] w_186552_21253# w_517669_21253# gpio_inp_dis[43] gpio_loopback_one[11]
+ w_21253_237565# w_692253_238870# w_23367_364074# gpio_dm0[40] gpio_inp_dis[23] gpio_dm2[21]
+ w_692253_283870# gpio_slow_sel[19] gpio_slow_sel[35] w_533874_1014469# gpio_analog_pol[22]
+ gpio_in[42] gpio_holdover[27] gpio_dm2[25] gpio_out[42] gpio_in[0] gpio_inp_dis[19]
+ gpio_slow_sel[18] w_694469_728352# gpio_holdover[43] gpio_analog_sel[7] w_692355_862552#
+ gpio_in_h[4] w_393474_1012253# gpio_holdover[23] w_694469_773352# gpio_oeb[9] analog_io[21]
+ gpio_analog_sel[2] gpio_loopback_one[0] gpio_slow_sel[2] gpio_dm2[40] gpio_loopback_one[15]
+ gpio_ib_mode_sel[30] w_23367_367165# w_21253_667565# gpio_in_h[31] w_23367_794074#
+ w_694469_103469# gpio_holdover[19] analog_io[42] gpio_dm0[41] gpio_analog_sel[13]
+ gpio_in[28] gpio_oeb[36] gpio_dm0[1] gpio_dm0[32] w_137274_1014469# w_353269_23367#
+ gpio_ib_mode_sel[8] gpio_slow_sel[29] gpio_oeb[38] gpio_analog_pol[5] gpio_analog_en[10]
+ gpio_loopback_one[33] gpio_in_h[14] gpio_dm0[5] analog_io[26] gpio_dm0[36] gpio_in_h[26]
+ gpio_in[40] gpio_dm1[32] gpio_analog_pol[0] w_21151_578074# gpio_analog_pol[16]
+ gpio_analog_en[11] gpio_loopback_one[4] gpio_slow_sel[24] gpio_oeb[3] w_243165_1014469#
+ gpio_dm0[9] gpio_ib_mode_sel[0] gpio_analog_pol[11] gpio_dm1[5] gpio[14] gpio[8]
+ gpio_dm1[36] gpio_dm2[41] gpio_analog_sel[33] gpio_dm2[1] gpio_dm2[32] w_23367_797165#
+ gpio_analog_en[12] analog_io[0] gpio_ib_mode_sel[12] w_21253_323965# gpio_vtrip_sel[41]
+ gpio_oeb[30] gpio[2] gpio_analog_sel[28] w_353269_21253# gpio_dm1[9] gpio_loopback_one[22]
+ gpio_in[25] gpio_in_h[9] gpio_analog_sel[42] gpio_loopback_one[37] analog_io[32]
+ gpio_dm2[5] analog_io[12] gpio_inp_dis[8] gpio_dm2[36] gpio_analog_en[13] gpio_analog_en[39]
+ w_23367_277674# w_694469_148669# gpio_slow_sel[42] gpio_analog_pol[36] gpio_slow_sel[7]
+ gpio_analog_sel[23] gpio_in[29] w_21253_581165# w_694469_193669# gpio_oeb[13] gpio_ib_mode_sel[33]
+ gpio_in_h[36] w_23367_707674# gpio_analog_pol[40] gpio_out[29] gpio[3] gpio_in[43]
+ gpio_analog_en[14] gpio_loopback_one[8] gpio_analog_pol[31] w_21151_234474# analog_io[5]
+ gpio_inp_dis[4] gpio_in_h[38] gpio_inp_dis[36] w_243165_1012355# gpio_dm0[14] gpio_in[7]
+ w_23367_963874# gpio_in[41] gpio_dm1[10] gpio_analog_pol[26] gpio_analog_en[15]
+ analog_io[37] analog_io[17] gpio_dm0[22] gpio_inp_dis[15] gpio_in_h[41] w_694469_238869#
+ gpio[10] w_21253_753965# gpio_loopback_one[26] gpio_inp_dis[0] gpio_out[30] gpio_dm0[18]
+ w_694469_283869# gpio_analog_pol[21] gpio_inp_dis[32] gpio_dm1[14] w_692253_865870#
+ gpio_inp_dis[28] gpio_in_h[3] gpio[15] gpio_dm2[10] gpio_holdover[4] gpio_in[22]
+ w_536965_1014469# gpio_oeb[8] gpio_dm0[26] gpio_holdover[36] gpio_ib_mode_sel[3]
+ gpio_dm1[22] w_298469_23367# gpio_inp_dis[11] w_191765_1014469# gpio_slow_sel[1]
+ w_694469_547952# w_482474_1014469# gpio_analog_sel[6] w_692355_638152# gpio_slow_sel[40]
+ gpio_dm1[18] w_635674_1014469# gpio_ib_mode_sel[15] gpio_in_h[30] gpio_inp_dis[38]
+ gpio_dm2[14] gpio_inp_dis[24] gpio_out[20] gpio_out[31] w_21151_664474# gpio_slow_sel[39]
+ gpio_holdover[0] gpio_oeb[19] gpio_oeb[35] gpio[4] w_23367_191274# w_23367_966965#
+ gpio_analog_sel[1] vssd_pad gpio_holdover[28] gpio_analog_sel[17] w_240074_1012253#
+ gpio_dm2[22] w_408069_23367# gpio_loopback_one[12] gpio_in[4] gpio[12] gpio_vtrip_sel[6]
+ gpio_dm2[18] w_694469_593152# gpio_vtrip_sel[29] gpio_in_h[13] w_23367_621274# gpio_analog_pol[9]
+ gpio_analog_sel[12] gpio[35] gpio_oeb[18] gpio[16] gpio_ib_mode_sel[36] gpio_inp_dis[40]
+ gpio_in[13] gpio_in_h[25] gpio_dm2[26] gpio_out[21] gpio_out[32] gpio_slow_sel[11]
+ gpio_holdover[38] gpio_holdover[24] analog_io[25] w_692355_728352# gpio_vtrip_sel[40]
+ gpio_analog_pol[4] gpio_vtrip_sel[7] gpio_vtrip_sel[30] w_514352_23367# gpio_loopback_one[30]
+ w_694469_325552# gpio_dm0[43] gpio_slow_sel[23] w_536965_1012355# gpio_oeb[2] gpio_in[19]
+ w_692355_773352# gpio[31] gpio[41] w_298469_21253# w_191765_1012355# gpio_dm0[29]
+ gpio_analog_pol[15] gpio[38] gpio[33] gpio_analog_sel[37] gpio_vtrip_sel[8] gpio_holdover[20]
+ gpio_dm0[42] gpio[20] gpio_vtrip_sel[31] gpio[13] w_694469_683352# w_21253_367165#
+ gpio_out[22] gpio_out[33] gpio_dm1[38] gpio_loopback_one[1] gpio_holdover[40] xres_buf_0/VGND
+ w_23367_194365# w_21151_320874# gpio_dm1[43] gpio[11] gpio_in[36] gpio_loopback_one[16]
+ gpio[21] gpio_in_h[8] gpio_analog_pol[10] gpio_dm0[2] gpio_analog_sel[32] w_408069_21253#
+ gpio_dm0[33] gpio[30] gpio_vtrip_sel[9] gpio_ib_mode_sel[27] gpio_vtrip_sel[32]
+ w_23367_624365# gpio_ib_mode_sel[6] gpio[37] gpio_in[1] gpio[24] gpio_slow_sel[6]
+ analog_io[31] gpio_dm1[42] gpio[6] analog_io[11] gpio_dm0[38] gpio_oeb[12] gpio_dm2[43]
+ gpio_vtrip_sel[20] gpio_analog_sel[27] gpio_loopback_one[19] gpio_in_h[19] gpio[5]
+ gpio[29] gpio_ib_mode_sel[18] gpio_in_h[35] gpio_dm0[6] gpio[9] gpio_out[23] gpio_out[34]
+ gpio_loopback_one[34] gpio_in[10] gpio_dm0[37] gpio_oeb[24] gpio_vtrip_sel[33] gpio_dm1[33]
+ gpio_loopback_one[38] gpio[40] gpio_dm2[29] w_514352_21253# gpio_analog_pol[35]
+ gpio[34] w_533874_1012253# gpio[36] gpio_slow_sel[33] gpio_analog_sel[22] gpio[18]
+ gpio_dm2[42] gpio_vtrip_sel[21] analog_io[4] gpio_dm2[38] w_404752_23367# gpio_in_h[18]
+ gpio_ib_mode_sel[19] gpio_dm1[6] gpio_loopback_one[5] gpio[43] gpio[7] gpio_analog_pol[30]
+ gpio_vtrip_sel[34] gpio_dm1[37] vssa_pad gpio_dm2[2] w_21253_797165# gpio_dm2[33]
+ w_21151_750874# gpio_out[24] gpio[17] gpio_out[35] analog_io[36] gpio[22] gpio_slow_sel[16]
+ SUB
Xclock_pad gpio_in_h[38] analog_io[38] clock_pad/PAD_A_ESD_1_H gpio_dm2[38] gpio_dm0[38]
+ gpio_dm1[38] gpio_in[38] gpio_inp_dis[38] gpio_ib_mode_sel[38] porb_h porb_h clock_pad/TIE_LO_ESD
+ gpio_oeb[38] clock_pad/HLD_H_N clock_pad/TIE_LO_ESD gpio_slow_sel[38] gpio_vtrip_sel[38]
+ gpio_holdover[38] gpio_analog_en[38] gpio_analog_sel[38] gpio_loopback_one[38] clock_pad/TIE_LO_ESD
+ gpio_analog_pol[38] gpio_out[38] vddio w_189869_21253# clock_pad/HLD_H_N SUB w_186552_21253#
+ vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda w_186552_23367# vddio SUB
+ w_189869_23367# gpio[38] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[17\] gpio_in_h[36] analog_io[36] mprj_pads.area2_io_pad\[17\]/PAD_A_ESD_1_H
+ gpio_dm2[36] gpio_dm1[36] gpio_dm0[36] gpio_in[36] gpio_inp_dis[36] gpio_ib_mode_sel[36]
+ porb_h porb_h mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD gpio_oeb[36] mprj_pads.area2_io_pad\[17\]/HLD_H_N
+ mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD gpio_slow_sel[36] gpio_vtrip_sel[36] gpio_holdover[36]
+ gpio_analog_en[36] gpio_analog_sel[36] gpio_loopback_one[36] mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD
+ gpio_analog_pol[36] gpio_out[36] vddio w_21151_234474# mprj_pads.area2_io_pad\[17\]/HLD_H_N
+ SUB w_21253_237565# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_237565#
+ vddio SUB w_23367_234474# gpio[36] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vccd_lvclamp_pad vdda vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vccd vccd vddio
+ vddio vddio SUB SUB sky130_ef_io__vccd_lvc_clamped_pad
Xmprj_pads.area2_io_pad\[7\] gpio_in_h[26] analog_io[26] mprj_pads.area2_io_pad\[7\]/PAD_A_ESD_1_H
+ gpio_dm2[26] gpio_dm1[26] gpio_dm0[26] gpio_in[26] gpio_inp_dis[26] gpio_ib_mode_sel[26]
+ porb_h porb_h mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD gpio_oeb[26] mprj_pads.area2_io_pad\[7\]/HLD_H_N
+ mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD gpio_slow_sel[26] gpio_vtrip_sel[26] gpio_holdover[26]
+ gpio_analog_en[26] gpio_analog_sel[26] gpio_loopback_one[26] mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD
+ gpio_analog_pol[26] gpio_out[26] vddio w_21151_750874# mprj_pads.area2_io_pad\[7\]/HLD_H_N
+ SUB w_21253_753965# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_753965#
+ vddio SUB w_23367_750874# gpio[26] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_2 gpio_loopback_zero[41] vccd gpio_loopback_one[41] SUB constant_block
Xmprj_pads.area1_io_pad\[7\] gpio_in_h[7] analog_io[7] mprj_pads.area1_io_pad\[7\]/PAD_A_ESD_1_H
+ gpio_dm2[7] gpio_dm1[7] gpio_dm0[7] gpio_in[7] gpio_inp_dis[7] gpio_ib_mode_sel[7]
+ porb_h porb_h mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD gpio_oeb[7] mprj_pads.area1_io_pad\[7\]/HLD_H_N
+ mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD gpio_slow_sel[7] gpio_vtrip_sel[7] gpio_holdover[7]
+ gpio_analog_en[7] gpio_analog_sel[7] gpio_loopback_one[7] mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD
+ gpio_analog_pol[7] gpio_out[7] vddio w_694469_551269# mprj_pads.area1_io_pad\[7\]/HLD_H_N
+ SUB w_694469_547952# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_547952#
+ vddio SUB w_692253_551270# gpio[7] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_3 gpio_loopback_zero[40] vccd gpio_loopback_one[40] SUB constant_block
Xmprj_pads.area1_io_pad\[11\] gpio_in_h[11] analog_io[11] mprj_pads.area1_io_pad\[11\]/PAD_A_ESD_1_H
+ gpio_dm2[11] gpio_dm1[11] gpio_dm0[11] gpio_in[11] gpio_inp_dis[11] gpio_ib_mode_sel[11]
+ porb_h porb_h mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD gpio_oeb[11] mprj_pads.area1_io_pad\[11\]/HLD_H_N
+ mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD gpio_slow_sel[11] gpio_vtrip_sel[11] gpio_holdover[11]
+ gpio_analog_en[11] gpio_analog_sel[11] gpio_loopback_one[11] mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD
+ gpio_analog_pol[11] gpio_out[11] vddio w_694469_731669# mprj_pads.area1_io_pad\[11\]/HLD_H_N
+ SUB w_694469_728352# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_728352#
+ vddio SUB w_692253_731670# gpio[11] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_4 gpio_loopback_zero[39] vccd gpio_loopback_one[39] SUB constant_block
Xmprj_pads.area2_io_pad\[15\] gpio_in_h[34] analog_io[34] mprj_pads.area2_io_pad\[15\]/PAD_A_ESD_1_H
+ gpio_dm2[34] gpio_dm1[34] gpio_dm0[34] gpio_in[34] gpio_inp_dis[34] gpio_ib_mode_sel[34]
+ porb_h porb_h mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD gpio_oeb[34] mprj_pads.area2_io_pad\[15\]/HLD_H_N
+ mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD gpio_slow_sel[34] gpio_vtrip_sel[34] gpio_holdover[34]
+ gpio_analog_en[34] gpio_analog_sel[34] gpio_loopback_one[34] mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD
+ gpio_analog_pol[34] gpio_out[34] vddio w_21151_320874# mprj_pads.area2_io_pad\[15\]/HLD_H_N
+ SUB w_21253_323965# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_323965#
+ vddio SUB w_23367_320874# gpio[34] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_5 gpio_loopback_zero[38] vccd gpio_loopback_one[38] SUB constant_block
Xsimple_por_0 vddio vccd porb_h por_l porb_l SUB SUB simple_por
Xmprj_pads.area2_io_pad\[5\] gpio_in_h[24] analog_io[24] mprj_pads.area2_io_pad\[5\]/PAD_A_ESD_1_H
+ gpio_dm2[24] gpio_dm1[24] gpio_dm0[24] gpio_in[24] gpio_inp_dis[24] gpio_ib_mode_sel[24]
+ porb_h porb_h mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD gpio_oeb[24] mprj_pads.area2_io_pad\[5\]/HLD_H_N
+ mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD gpio_slow_sel[24] gpio_vtrip_sel[24] gpio_holdover[24]
+ gpio_analog_en[24] gpio_analog_sel[24] gpio_loopback_one[24] mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD
+ gpio_analog_pol[24] gpio_out[24] vddio w_21151_963874# mprj_pads.area2_io_pad\[5\]/HLD_H_N
+ SUB w_21253_966965# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_966965#
+ vddio SUB w_23367_963874# gpio[24] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area1_io_pad\[5\] gpio_in_h[5] analog_io[5] mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_1_H
+ gpio_dm2[5] gpio_dm1[5] gpio_dm0[5] gpio_in[5] gpio_inp_dis[5] gpio_ib_mode_sel[5]
+ porb_h porb_h mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD gpio_oeb[5] mprj_pads.area1_io_pad\[5\]/HLD_H_N
+ mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD gpio_slow_sel[5] gpio_vtrip_sel[5] gpio_holdover[5]
+ gpio_analog_en[5] gpio_analog_sel[5] gpio_loopback_one[5] mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD
+ gpio_analog_pol[5] gpio_out[5] vddio w_694469_328869# mprj_pads.area1_io_pad\[5\]/HLD_H_N
+ SUB w_694469_325552# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_325552#
+ vddio SUB w_692253_328870# gpio[5] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_6 constant_block_6/zero vccd constant_block_6/one SUB constant_block
Xconstant_block_7 SUB vccd gpio_loopback_one[36] SUB constant_block
Xmgmt_vddio_hvclamp_pad\[0\] SUB vdda SUB SUB vddio gpio_pad/AMUXBUS_B vddio gpio_pad/AMUXBUS_A
+ vccd vccd vddio SUB sky130_ef_io__vddio_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[13\] gpio_in_h[32] analog_io[32] mprj_pads.area2_io_pad\[13\]/PAD_A_ESD_1_H
+ gpio_dm2[32] gpio_dm1[32] gpio_dm0[32] gpio_in[32] gpio_inp_dis[32] gpio_ib_mode_sel[32]
+ porb_h porb_h mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD gpio_oeb[32] mprj_pads.area2_io_pad\[13\]/HLD_H_N
+ mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD gpio_slow_sel[32] gpio_vtrip_sel[32] gpio_holdover[32]
+ gpio_analog_en[32] gpio_analog_sel[32] gpio_loopback_one[32] mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD
+ gpio_analog_pol[32] gpio_out[32] vddio w_21151_407274# mprj_pads.area2_io_pad\[13\]/HLD_H_N
+ SUB w_21253_410365# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_410365#
+ vddio SUB w_23367_407274# gpio[32] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_8 SUB vccd gpio_loopback_one[37] SUB constant_block
Xmgmt_vssio_hvclamp_pad\[1\] vdda2 SUB SUB gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A SUB
+ vddio vddio SUB vddio vccd vccd sky130_ef_io__vssio_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[3\] gpio_in_h[22] analog_io[22] mprj_pads.area2_io_pad\[3\]/PAD_A_ESD_1_H
+ gpio_dm2[22] gpio_dm1[22] gpio_dm0[22] gpio_in[22] gpio_inp_dis[22] gpio_ib_mode_sel[22]
+ porb_h porb_h mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD gpio_oeb[22] mprj_pads.area2_io_pad\[3\]/HLD_H_N
+ mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD gpio_slow_sel[22] gpio_vtrip_sel[22] gpio_holdover[22]
+ gpio_analog_en[22] gpio_analog_sel[22] gpio_loopback_one[22] mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD
+ gpio_analog_pol[22] gpio_out[22] vddio w_137274_1014469# mprj_pads.area2_io_pad\[3\]/HLD_H_N
+ SUB w_140365_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_140365_1012355#
+ vddio SUB w_137274_1012253# gpio[22] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_9 SUB vccd gpio_loopback_one[22] SUB constant_block
Xmprj_pads.area1_io_pad\[3\] gpio_in_h[3] analog_io[3] mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_1_H
+ gpio_dm2[3] gpio_dm1[3] gpio_dm0[3] gpio_in[3] gpio_inp_dis[3] gpio_ib_mode_sel[3]
+ porb_h porb_h mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD gpio_oeb[3] mprj_pads.area1_io_pad\[3\]/HLD_H_N
+ mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD gpio_slow_sel[3] gpio_vtrip_sel[3] gpio_holdover[3]
+ gpio_analog_en[3] gpio_analog_sel[3] gpio_loopback_one[3] mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD
+ gpio_analog_pol[3] gpio_out[3] vddio w_694469_238869# mprj_pads.area1_io_pad\[3\]/HLD_H_N
+ SUB w_694469_235552# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_235552#
+ vddio SUB w_692253_238870# gpio[3] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser2_vdda_hvclamp_pad SUB vdda2 SUB vccd vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vddio vccd vdda2 SUB SUB vddio sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[18\] gpio_in_h[18] analog_io[18] mprj_pads.area1_io_pad\[18\]/PAD_A_ESD_1_H
+ gpio_dm2[18] gpio_dm1[18] gpio_dm0[18] gpio_in[18] gpio_inp_dis[18] gpio_ib_mode_sel[18]
+ porb_h porb_h mprj_pads.area1_io_pad\[18\]/TIE_LO_ESD gpio_oeb[18] mprj_pads.area1_io_pad\[18\]/HLD_H_N
+ mprj_pads.area1_io_pad\[18\]/TIE_LO_ESD gpio_slow_sel[18] gpio_vtrip_sel[18] gpio_holdover[18]
+ gpio_analog_en[18] gpio_analog_sel[18] gpio_loopback_one[18] mprj_pads.area1_io_pad\[18\]/TIE_LO_ESD
+ gpio_analog_pol[18] gpio_out[18] vddio w_393474_1014469# mprj_pads.area1_io_pad\[18\]/HLD_H_N
+ SUB w_396565_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_396565_1012355#
+ vddio SUB w_393474_1012253# gpio[18] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[11\] gpio_in_h[30] analog_io[30] mprj_pads.area2_io_pad\[11\]/PAD_A_ESD_1_H
+ gpio_dm2[30] gpio_dm1[30] gpio_dm0[30] gpio_in[30] gpio_inp_dis[30] gpio_ib_mode_sel[30]
+ porb_h porb_h mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD gpio_oeb[30] mprj_pads.area2_io_pad\[11\]/HLD_H_N
+ mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD gpio_slow_sel[30] gpio_vtrip_sel[30] gpio_holdover[30]
+ gpio_analog_en[30] gpio_analog_sel[30] gpio_loopback_one[30] mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD
+ gpio_analog_pol[30] gpio_out[30] vddio w_21151_578074# mprj_pads.area2_io_pad\[11\]/HLD_H_N
+ SUB w_21253_581165# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_581165#
+ vddio SUB w_23367_578074# gpio[30] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[1\] gpio_in_h[20] analog_io[20] mprj_pads.area2_io_pad\[1\]/PAD_A_ESD_1_H
+ gpio_dm2[20] gpio_dm1[20] gpio_dm0[20] gpio_in[20] gpio_inp_dis[20] gpio_ib_mode_sel[20]
+ porb_h porb_h mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD gpio_oeb[20] mprj_pads.area2_io_pad\[1\]/HLD_H_N
+ mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD gpio_slow_sel[20] gpio_vtrip_sel[20] gpio_holdover[20]
+ gpio_analog_en[20] gpio_analog_sel[20] gpio_loopback_one[20] mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD
+ gpio_analog_pol[20] gpio_out[20] vddio w_240074_1014469# mprj_pads.area2_io_pad\[1\]/HLD_H_N
+ SUB w_243165_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_243165_1012355#
+ vddio SUB w_240074_1012253# gpio[20] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area1_io_pad\[1\] gpio_in_h[1] analog_io[1] mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_1_H
+ gpio_dm2[1] gpio_dm1[1] gpio_dm0[1] gpio_in[1] gpio_inp_dis[1] gpio_ib_mode_sel[1]
+ porb_h porb_h mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD gpio_oeb[1] mprj_pads.area1_io_pad\[1\]/HLD_H_N
+ mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD gpio_slow_sel[1] gpio_vtrip_sel[1] gpio_holdover[1]
+ gpio_analog_en[1] gpio_analog_sel[1] gpio_loopback_one[1] mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD
+ gpio_analog_pol[1] gpio_out[1] vddio w_694469_148669# mprj_pads.area1_io_pad\[1\]/HLD_H_N
+ SUB w_694469_145352# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_145352#
+ vddio SUB w_692253_148670# gpio[1] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vssd_lvclamp_pad SUB vdda1 vddio SUB vccd1 SUB vddio vccd vccd gpio_pad/AMUXBUS_B
+ vddio gpio_pad/AMUXBUS_A SUB sky130_ef_io__vssd_lvc_clamped3_pad
Xgpio_pad gpio_in_h[43] analog_io[43] gpio_pad/PAD_A_ESD_1_H gpio_dm2[43] gpio_dm1[43]
+ gpio_dm0[43] gpio_in[43] gpio_inp_dis[43] gpio_ib_mode_sel[43] porb_h porb_h gpio_pad/TIE_LO_ESD
+ gpio_oeb[43] gpio_pad/HLD_H_N gpio_pad/TIE_LO_ESD gpio_slow_sel[43] gpio_vtrip_sel[43]
+ gpio_holdover[43] gpio_analog_en[43] gpio_analog_sel[43] gpio_loopback_one[43] gpio_pad/TIE_LO_ESD
+ gpio_analog_pol[43] gpio_out[43] vddio w_517669_21253# gpio_pad/HLD_H_N SUB w_514352_21253#
+ vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda w_514352_23367# vddio SUB
+ w_517669_23367# gpio[43] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area1_io_pad\[16\] gpio_in_h[16] analog_io[16] mprj_pads.area1_io_pad\[16\]/PAD_A_ESD_1_H
+ gpio_dm2[16] gpio_dm1[16] gpio_dm0[16] gpio_in[16] gpio_inp_dis[16] gpio_ib_mode_sel[16]
+ porb_h porb_h mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD gpio_oeb[16] mprj_pads.area1_io_pad\[16\]/HLD_H_N
+ mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD gpio_slow_sel[16] gpio_vtrip_sel[16] gpio_holdover[16]
+ gpio_analog_en[16] gpio_analog_sel[16] gpio_loopback_one[16] mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD
+ gpio_analog_pol[16] gpio_out[16] vddio w_533874_1014469# mprj_pads.area1_io_pad\[16\]/HLD_H_N
+ SUB w_536965_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_536965_1012355#
+ vddio SUB w_533874_1012253# gpio[16] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[0\] SUB vdda1 SUB vccd vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vddio vccd vdda1 SUB SUB vddio sky130_ef_io__vdda_hvc_clamped_pad
Xmgmt_vssd_lvclamp_pad vdda vddio vssd_pad vddio vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vddio vccd SUB SUB sky130_ef_io__vssd_lvc_clamped_pad
Xuser2_vccd_lvclamp_pad vdda2 vccd vddio vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vccd vccd2 vccd2 SUB SUB vddio SUB sky130_ef_io__vccd_lvc_clamped3_pad
Xxres_buf_0 resetb_h resetb_l xres_buf_0/LVPWR xres_buf_0/LVGND xres_buf_0/VPWR xres_buf_0/VGND
+ xres_buf
Xmgmt_vssa_hvclamp_pad SUB vddio vssa_pad SUB vccd vddio SUB vddio vdda vccd SUB gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B sky130_ef_io__vssa_hvc_clamped_pad
Xuser1_vssa_hvclamp_pad\[1\] SUB vddio SUB SUB vccd vddio SUB vddio vdda1 vccd SUB
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[14\] gpio_in_h[14] analog_io[14] mprj_pads.area1_io_pad\[14\]/PAD_A_ESD_1_H
+ gpio_dm2[14] gpio_dm1[14] gpio_dm0[14] gpio_in[14] gpio_inp_dis[14] gpio_ib_mode_sel[14]
+ porb_h porb_h mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD gpio_oeb[14] mprj_pads.area1_io_pad\[14\]/HLD_H_N
+ mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD gpio_slow_sel[14] gpio_vtrip_sel[14] gpio_holdover[14]
+ gpio_analog_en[14] gpio_analog_sel[14] gpio_loopback_one[14] mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD
+ gpio_analog_pol[14] gpio_out[14] vddio w_694469_955069# mprj_pads.area1_io_pad\[14\]/HLD_H_N
+ SUB w_694469_951752# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_951752#
+ vddio SUB w_692253_955070# gpio[14] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser_id_programming_0 mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[14]
+ mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20]
+ mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27]
+ mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5]
+ mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[28] mask_rev[13] SUB vccd
+ user_id_programming
Xmprj_pads.area2_io_pad\[18\] gpio_in_h[37] analog_io[37] mprj_pads.area2_io_pad\[18\]/PAD_A_ESD_1_H
+ gpio_dm2[37] gpio_dm1[37] gpio_dm0[37] gpio_in[37] gpio_inp_dis[37] gpio_ib_mode_sel[37]
+ porb_h porb_h mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD gpio_oeb[37] mprj_pads.area2_io_pad\[18\]/HLD_H_N
+ mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD gpio_slow_sel[37] gpio_vtrip_sel[37] gpio_holdover[37]
+ gpio_analog_en[37] gpio_analog_sel[37] gpio_loopback_one[37] mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD
+ gpio_analog_pol[37] gpio_out[37] vddio w_21151_191274# mprj_pads.area2_io_pad\[18\]/HLD_H_N
+ SUB w_21253_194365# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_194365#
+ vddio SUB w_23367_191274# gpio[37] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[8\] gpio_in_h[27] analog_io[27] mprj_pads.area2_io_pad\[8\]/PAD_A_ESD_1_H
+ gpio_dm2[27] gpio_dm1[27] gpio_dm0[27] gpio_in[27] gpio_inp_dis[27] gpio_ib_mode_sel[27]
+ porb_h porb_h mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD gpio_oeb[27] mprj_pads.area2_io_pad\[8\]/HLD_H_N
+ mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD gpio_slow_sel[27] gpio_vtrip_sel[27] gpio_holdover[27]
+ gpio_analog_en[27] gpio_analog_sel[27] gpio_loopback_one[27] mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD
+ gpio_analog_pol[27] gpio_out[27] vddio w_21151_707674# mprj_pads.area2_io_pad\[8\]/HLD_H_N
+ SUB w_21253_710765# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_710765#
+ vddio SUB w_23367_707674# gpio[27] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area1_io_pad\[8\] gpio_in_h[8] analog_io[8] mprj_pads.area1_io_pad\[8\]/PAD_A_ESD_1_H
+ gpio_dm2[8] gpio_dm1[8] gpio_dm0[8] gpio_in[8] gpio_inp_dis[8] gpio_ib_mode_sel[8]
+ porb_h porb_h mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD gpio_oeb[8] mprj_pads.area1_io_pad\[8\]/HLD_H_N
+ mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD gpio_slow_sel[8] gpio_vtrip_sel[8] gpio_holdover[8]
+ gpio_analog_en[8] gpio_analog_sel[8] gpio_loopback_one[8] mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD
+ gpio_analog_pol[8] gpio_out[8] vddio w_694469_596469# mprj_pads.area1_io_pad\[8\]/HLD_H_N
+ SUB w_694469_593152# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_593152#
+ vddio SUB w_692253_596470# gpio[8] vccd sky130_ef_io__gpiov2_pad_wrapped
Xresetb_pad resetb_h xres_vss_loop constant_block_6/one xresloop porb_h xres_vss_loop
+ xres_vss_loop xres_vss_loop resetb_pad/TIE_HI_ESD xres_vss_loop xres_vss_loop SUB
+ gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vddio vdda vccd vccd SUB vddio SUB SUB
+ resetb_pad xresloop sky130_fd_io__top_xres4v2
Xconstant_block_40 SUB vccd gpio_loopback_one[5] SUB constant_block
Xmprj_pads.area1_io_pad\[12\] gpio_in_h[12] analog_io[12] mprj_pads.area1_io_pad\[12\]/PAD_A_ESD_1_H
+ gpio_dm2[12] gpio_dm1[12] gpio_dm0[12] gpio_in[12] gpio_inp_dis[12] gpio_ib_mode_sel[12]
+ porb_h porb_h mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD gpio_oeb[12] mprj_pads.area1_io_pad\[12\]/HLD_H_N
+ mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD gpio_slow_sel[12] gpio_vtrip_sel[12] gpio_holdover[12]
+ gpio_analog_en[12] gpio_analog_sel[12] gpio_loopback_one[12] mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD
+ gpio_analog_pol[12] gpio_out[12] vddio w_694469_776669# mprj_pads.area1_io_pad\[12\]/HLD_H_N
+ SUB w_694469_773352# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_773352#
+ vddio SUB w_692253_776670# gpio[12] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_30 SUB vccd gpio_loopback_one[28] SUB constant_block
Xconstant_block_41 SUB vccd gpio_loopback_one[4] SUB constant_block
Xmprj_pads.area2_io_pad\[16\] gpio_in_h[35] analog_io[35] mprj_pads.area2_io_pad\[16\]/PAD_A_ESD_1_H
+ gpio_dm2[35] gpio_dm1[35] gpio_dm0[35] gpio_in[35] gpio_inp_dis[35] gpio_ib_mode_sel[35]
+ porb_h porb_h mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD gpio_oeb[35] mprj_pads.area2_io_pad\[16\]/HLD_H_N
+ mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD gpio_slow_sel[35] gpio_vtrip_sel[35] gpio_holdover[35]
+ gpio_analog_en[35] gpio_analog_sel[35] gpio_loopback_one[35] mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD
+ gpio_analog_pol[35] gpio_out[35] vddio w_21151_277674# mprj_pads.area2_io_pad\[16\]/HLD_H_N
+ SUB w_21253_280765# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_280765#
+ vddio SUB w_23367_277674# gpio[35] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_20 SUB vccd gpio_loopback_one[13] SUB constant_block
Xmprj_pads.area2_io_pad\[6\] gpio_in_h[25] analog_io[25] mprj_pads.area2_io_pad\[6\]/PAD_A_ESD_1_H
+ gpio_dm2[25] gpio_dm1[25] gpio_dm0[25] gpio_in[25] gpio_inp_dis[25] gpio_ib_mode_sel[25]
+ porb_h porb_h mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD gpio_oeb[25] mprj_pads.area2_io_pad\[6\]/HLD_H_N
+ mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD gpio_slow_sel[25] gpio_vtrip_sel[25] gpio_holdover[25]
+ gpio_analog_en[25] gpio_analog_sel[25] gpio_loopback_one[25] mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD
+ gpio_analog_pol[25] gpio_out[25] vddio w_21151_794074# mprj_pads.area2_io_pad\[6\]/HLD_H_N
+ SUB w_21253_797165# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_797165#
+ vddio SUB w_23367_794074# gpio[25] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_31 SUB vccd gpio_loopback_one[27] SUB constant_block
Xconstant_block_42 SUB vccd gpio_loopback_one[3] SUB constant_block
Xflash_csb_pad gpio_in_h[39] analog_io[39] flash_csb_pad/PAD_A_ESD_1_H gpio_dm2[39]
+ gpio_dm1[39] gpio_dm0[39] gpio_in[39] gpio_inp_dis[39] gpio_ib_mode_sel[39] porb_h
+ porb_h flash_csb_pad/TIE_LO_ESD gpio_oeb[39] flash_csb_pad/HLD_H_N flash_csb_pad/TIE_LO_ESD
+ gpio_slow_sel[39] gpio_vtrip_sel[39] gpio_holdover[39] gpio_analog_en[39] gpio_analog_sel[39]
+ gpio_loopback_one[39] flash_csb_pad/TIE_LO_ESD gpio_analog_pol[39] gpio_out[39]
+ vddio w_298469_21253# flash_csb_pad/HLD_H_N SUB w_295152_21253# vccd gpio_pad/AMUXBUS_B
+ gpio_pad/AMUXBUS_A vddio vdda w_295152_23367# vddio SUB w_298469_23367# gpio[40]
+ vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area1_io_pad\[6\] gpio_in_h[6] analog_io[6] mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_1_H
+ gpio_dm2[6] gpio_dm1[6] gpio_dm0[6] gpio_in[6] gpio_inp_dis[6] gpio_ib_mode_sel[6]
+ porb_h porb_h mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD gpio_oeb[6] mprj_pads.area1_io_pad\[6\]/HLD_H_N
+ mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD gpio_slow_sel[6] gpio_vtrip_sel[6] gpio_holdover[6]
+ gpio_analog_en[6] gpio_analog_sel[6] gpio_loopback_one[6] mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD
+ gpio_analog_pol[6] gpio_out[6] vddio w_694469_374069# mprj_pads.area1_io_pad\[6\]/HLD_H_N
+ SUB w_694469_370752# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_370752#
+ vddio SUB w_692253_374070# gpio[6] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_10 SUB vccd gpio_loopback_one[21] SUB constant_block
Xconstant_block_21 SUB vccd gpio_loopback_one[11] SUB constant_block
Xconstant_block_32 SUB vccd gpio_loopback_one[26] SUB constant_block
Xconstant_block_43 SUB vccd gpio_loopback_one[2] SUB constant_block
Xmprj_pads.area1_io_pad\[10\] gpio_in_h[10] analog_io[10] mprj_pads.area1_io_pad\[10\]/PAD_A_ESD_1_H
+ gpio_dm2[10] gpio_dm1[10] gpio_dm0[10] gpio_in[10] gpio_inp_dis[10] gpio_ib_mode_sel[10]
+ porb_h porb_h mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD gpio_oeb[10] mprj_pads.area1_io_pad\[10\]/HLD_H_N
+ mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD gpio_slow_sel[10] gpio_vtrip_sel[10] gpio_holdover[10]
+ gpio_analog_en[10] gpio_analog_sel[10] gpio_loopback_one[10] mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD
+ gpio_analog_pol[10] gpio_out[10] vddio w_694469_686669# mprj_pads.area1_io_pad\[10\]/HLD_H_N
+ SUB w_694469_683352# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_683352#
+ vddio SUB w_692253_686670# gpio[10] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_11 SUB vccd gpio_loopback_one[20] SUB constant_block
Xconstant_block_22 SUB vccd gpio_loopback_one[23] SUB constant_block
Xconstant_block_33 SUB vccd gpio_loopback_one[25] SUB constant_block
Xconstant_block_44 SUB vccd gpio_loopback_one[1] SUB constant_block
Xflash_io1_pad gpio_in_h[42] analog_io[42] flash_io1_pad/PAD_A_ESD_1_H gpio_dm2[42]
+ gpio_dm1[42] gpio_dm0[42] gpio_in[42] gpio_inp_dis[42] gpio_ib_mode_sel[42] porb_h
+ porb_h flash_io1_pad/TIE_LO_ESD gpio_oeb[42] flash_io1_pad/HLD_H_N flash_io1_pad/TIE_LO_ESD
+ gpio_slow_sel[42] gpio_vtrip_sel[42] gpio_holdover[42] gpio_analog_en[42] gpio_analog_sel[42]
+ gpio_loopback_one[42] flash_io1_pad/TIE_LO_ESD gpio_analog_pol[42] gpio_out[42]
+ vddio w_462869_21253# flash_io1_pad/HLD_H_N SUB w_459552_21253# vccd gpio_pad/AMUXBUS_B
+ gpio_pad/AMUXBUS_A vddio vdda w_459552_23367# vddio SUB w_462869_23367# gpio[42]
+ vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vddio_hvclamp_pad\[1\] SUB vdda2 SUB SUB vddio gpio_pad/AMUXBUS_B vddio gpio_pad/AMUXBUS_A
+ vccd vccd vddio SUB sky130_ef_io__vddio_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[14\] gpio_in_h[33] analog_io[33] mprj_pads.area2_io_pad\[14\]/PAD_A_ESD_1_H
+ gpio_dm2[33] gpio_dm1[33] gpio_dm0[33] gpio_in[33] gpio_inp_dis[33] gpio_ib_mode_sel[33]
+ porb_h porb_h mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD gpio_oeb[33] mprj_pads.area2_io_pad\[14\]/HLD_H_N
+ mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD gpio_slow_sel[33] gpio_vtrip_sel[33] gpio_holdover[33]
+ gpio_analog_en[33] gpio_analog_sel[33] gpio_loopback_one[33] mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD
+ gpio_analog_pol[33] gpio_out[33] vddio w_21151_364074# mprj_pads.area2_io_pad\[14\]/HLD_H_N
+ SUB w_21253_367165# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_367165#
+ vddio SUB w_23367_364074# gpio[33] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_12 SUB vccd gpio_loopback_one[19] SUB constant_block
Xconstant_block_34 SUB vccd gpio_loopback_one[24] SUB constant_block
Xconstant_block_23 SUB vccd gpio_loopback_one[35] SUB constant_block
Xmprj_pads.area2_io_pad\[4\] gpio_in_h[23] analog_io[23] mprj_pads.area2_io_pad\[4\]/PAD_A_ESD_1_H
+ gpio_dm2[23] gpio_dm1[23] gpio_dm0[23] gpio_in[23] gpio_inp_dis[23] gpio_ib_mode_sel[23]
+ porb_h porb_h mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD gpio_oeb[23] mprj_pads.area2_io_pad\[4\]/HLD_H_N
+ mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD gpio_slow_sel[23] gpio_vtrip_sel[23] gpio_holdover[23]
+ gpio_analog_en[23] gpio_analog_sel[23] gpio_loopback_one[23] mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD
+ gpio_analog_pol[23] gpio_out[23] vddio w_85874_1014469# mprj_pads.area2_io_pad\[4\]/HLD_H_N
+ SUB w_88965_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_88965_1012355#
+ vddio SUB w_85874_1012253# gpio[23] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_13 SUB vccd gpio_loopback_one[18] SUB constant_block
Xconstant_block_35 SUB vccd gpio_loopback_one[10] SUB constant_block
Xconstant_block_24 SUB vccd gpio_loopback_one[34] SUB constant_block
Xmprj_pads.area1_io_pad\[4\] gpio_in_h[4] analog_io[4] mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_1_H
+ gpio_dm2[4] gpio_dm1[4] gpio_dm0[4] gpio_in[4] gpio_inp_dis[4] gpio_ib_mode_sel[4]
+ porb_h porb_h mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD gpio_oeb[4] mprj_pads.area1_io_pad\[4\]/HLD_H_N
+ mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD gpio_slow_sel[4] gpio_vtrip_sel[4] gpio_holdover[4]
+ gpio_analog_en[4] gpio_analog_sel[4] gpio_loopback_one[4] mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD
+ gpio_analog_pol[4] gpio_out[4] vddio w_694469_283869# mprj_pads.area1_io_pad\[4\]/HLD_H_N
+ SUB w_694469_280552# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_280552#
+ vddio SUB w_692253_283870# gpio[4] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_14 SUB vccd gpio_loopback_one[17] SUB constant_block
Xconstant_block_36 SUB vccd gpio_loopback_one[9] SUB constant_block
Xconstant_block_25 SUB vccd gpio_loopback_one[33] SUB constant_block
Xuser2_vssd_lvclamp_pad SUB vdda2 vddio SUB vccd2 SUB vddio vccd vccd gpio_pad/AMUXBUS_B
+ vddio gpio_pad/AMUXBUS_A SUB sky130_ef_io__vssd_lvc_clamped3_pad
Xconstant_block_15 SUB vccd gpio_loopback_one[16] SUB constant_block
Xconstant_block_37 SUB vccd gpio_loopback_one[8] SUB constant_block
Xmprj_pads.area2_io_pad\[12\] gpio_in_h[31] analog_io[31] mprj_pads.area2_io_pad\[12\]/PAD_A_ESD_1_H
+ gpio_dm2[31] gpio_dm1[31] gpio_dm0[31] gpio_in[31] gpio_inp_dis[31] gpio_ib_mode_sel[31]
+ porb_h porb_h mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD gpio_oeb[31] mprj_pads.area2_io_pad\[12\]/HLD_H_N
+ mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD gpio_slow_sel[31] gpio_vtrip_sel[31] gpio_holdover[31]
+ gpio_analog_en[31] gpio_analog_sel[31] gpio_loopback_one[31] mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD
+ gpio_analog_pol[31] gpio_out[31] vddio w_21151_534874# mprj_pads.area2_io_pad\[12\]/HLD_H_N
+ SUB w_21253_537965# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_537965#
+ vddio SUB w_23367_534874# gpio[31] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_26 SUB vccd gpio_loopback_one[32] SUB constant_block
Xmgmt_vssio_hvclamp_pad\[0\] vdda SUB SUB gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vssio_pad
+ vddio vddio SUB vddio vccd vccd sky130_ef_io__vssio_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[2\] gpio_in_h[21] analog_io[21] mprj_pads.area2_io_pad\[2\]/PAD_A_ESD_1_H
+ gpio_dm2[21] gpio_dm1[21] gpio_dm0[21] gpio_in[21] gpio_inp_dis[21] gpio_ib_mode_sel[21]
+ porb_h porb_h mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD gpio_oeb[21] mprj_pads.area2_io_pad\[2\]/HLD_H_N
+ mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD gpio_slow_sel[21] gpio_vtrip_sel[21] gpio_holdover[21]
+ gpio_analog_en[21] gpio_analog_sel[21] gpio_loopback_one[21] mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD
+ gpio_analog_pol[21] gpio_out[21] vddio w_188674_1014469# mprj_pads.area2_io_pad\[2\]/HLD_H_N
+ SUB w_191765_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_191765_1012355#
+ vddio SUB w_188674_1012253# gpio[21] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_38 SUB vccd gpio_loopback_one[7] SUB constant_block
Xconstant_block_27 SUB vccd gpio_loopback_one[31] SUB constant_block
Xconstant_block_16 SUB vccd gpio_loopback_one[0] SUB constant_block
Xuser2_vssa_hvclamp_pad SUB vddio SUB SUB vccd vddio SUB vddio vdda2 vccd SUB gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[2\] gpio_in_h[2] analog_io[2] mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_1_H
+ gpio_dm2[2] gpio_dm1[2] gpio_dm0[2] gpio_in[2] gpio_inp_dis[2] gpio_ib_mode_sel[2]
+ porb_h porb_h mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD gpio_oeb[2] mprj_pads.area1_io_pad\[2\]/HLD_H_N
+ mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD gpio_slow_sel[2] gpio_vtrip_sel[2] gpio_holdover[2]
+ gpio_analog_en[2] gpio_analog_sel[2] gpio_loopback_one[2] mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD
+ gpio_analog_pol[2] gpio_out[2] vddio w_694469_193669# mprj_pads.area1_io_pad\[2\]/HLD_H_N
+ SUB w_694469_190352# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_190352#
+ vddio SUB w_692253_193670# gpio[2] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_17 SUB vccd gpio_loopback_one[15] SUB constant_block
Xconstant_block_28 SUB vccd gpio_loopback_one[30] SUB constant_block
Xconstant_block_39 SUB vccd gpio_loopback_one[6] SUB constant_block
Xmprj_pads.area1_io_pad\[17\] gpio_in_h[17] analog_io[17] mprj_pads.area1_io_pad\[17\]/PAD_A_ESD_1_H
+ gpio_dm2[17] gpio_dm1[17] gpio_dm0[17] gpio_in[17] gpio_inp_dis[17] gpio_ib_mode_sel[17]
+ porb_h porb_h mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD gpio_oeb[17] mprj_pads.area1_io_pad\[17\]/HLD_H_N
+ mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD gpio_slow_sel[17] gpio_vtrip_sel[17] gpio_holdover[17]
+ gpio_analog_en[17] gpio_analog_sel[17] gpio_loopback_one[17] mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD
+ gpio_analog_pol[17] gpio_out[17] vddio w_482474_1014469# mprj_pads.area1_io_pad\[17\]/HLD_H_N
+ SUB w_485565_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_485565_1012355#
+ vddio SUB w_482474_1012253# gpio[17] vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[1\] SUB vdda1 SUB vccd vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vddio vccd vdda1 SUB SUB vddio sky130_ef_io__vdda_hvc_clamped_pad
Xconstant_block_18 SUB vccd gpio_loopback_one[14] SUB constant_block
Xconstant_block_29 SUB vccd gpio_loopback_one[29] SUB constant_block
Xmprj_pads.area2_io_pad\[10\] gpio_in_h[29] analog_io[29] mprj_pads.area2_io_pad\[10\]/PAD_A_ESD_1_H
+ gpio_dm2[29] gpio_dm1[29] gpio_dm0[29] gpio_in[29] gpio_inp_dis[29] gpio_ib_mode_sel[29]
+ porb_h porb_h mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD gpio_oeb[29] mprj_pads.area2_io_pad\[10\]/HLD_H_N
+ mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD gpio_slow_sel[29] gpio_vtrip_sel[29] gpio_holdover[29]
+ gpio_analog_en[29] gpio_analog_sel[29] gpio_loopback_one[29] mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD
+ gpio_analog_pol[29] gpio_out[29] vddio w_21151_621274# mprj_pads.area2_io_pad\[10\]/HLD_H_N
+ SUB w_21253_624365# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_624365#
+ vddio SUB w_23367_621274# gpio[29] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[0\] gpio_in_h[19] analog_io[19] mprj_pads.area2_io_pad\[0\]/PAD_A_ESD_1_H
+ gpio_dm2[19] gpio_dm1[19] gpio_dm0[19] gpio_in[19] gpio_inp_dis[19] gpio_ib_mode_sel[19]
+ porb_h porb_h mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD gpio_oeb[19] mprj_pads.area2_io_pad\[0\]/HLD_H_N
+ mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD gpio_slow_sel[19] gpio_vtrip_sel[19] gpio_holdover[19]
+ gpio_analog_en[19] gpio_analog_sel[19] gpio_loopback_one[19] mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD
+ gpio_analog_pol[19] gpio_out[19] vddio w_291674_1014469# mprj_pads.area2_io_pad\[0\]/HLD_H_N
+ SUB w_294765_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_294765_1012355#
+ vddio SUB w_291674_1012253# gpio[19] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_19 SUB vccd gpio_loopback_one[12] SUB constant_block
Xmprj_pads.area1_io_pad\[0\] gpio_in_h[0] analog_io[0] mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_1_H
+ gpio_dm2[0] gpio_dm1[0] gpio_dm0[0] gpio_in[0] gpio_inp_dis[0] gpio_ib_mode_sel[0]
+ porb_h porb_h mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD gpio_oeb[0] mprj_pads.area1_io_pad\[0\]/HLD_H_N
+ mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD gpio_slow_sel[0] gpio_vtrip_sel[0] gpio_holdover[0]
+ gpio_analog_en[0] gpio_analog_sel[0] gpio_loopback_one[0] mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD
+ gpio_analog_pol[0] gpio_out[0] vddio w_694469_103469# mprj_pads.area1_io_pad\[0\]/HLD_H_N
+ SUB w_694469_100152# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_100152#
+ vddio SUB w_692253_103470# gpio[0] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmgmt_vdda_hvclamp_pad SUB vdda_pad SUB vccd vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vddio vccd vdda SUB SUB vddio sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[15\] gpio_in_h[15] analog_io[15] mprj_pads.area1_io_pad\[15\]/PAD_A_ESD_1_H
+ gpio_dm2[15] gpio_dm1[15] gpio_dm0[15] gpio_in[15] gpio_inp_dis[15] gpio_ib_mode_sel[15]
+ porb_h porb_h mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD gpio_oeb[15] mprj_pads.area1_io_pad\[15\]/HLD_H_N
+ mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD gpio_slow_sel[15] gpio_vtrip_sel[15] gpio_holdover[15]
+ gpio_analog_en[15] gpio_analog_sel[15] gpio_loopback_one[15] mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD
+ gpio_analog_pol[15] gpio_out[15] vddio w_635674_1014469# mprj_pads.area1_io_pad\[15\]/HLD_H_N
+ SUB w_638765_1014469# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_638765_1012355#
+ vddio SUB w_635674_1012253# gpio[15] vccd sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[9\] gpio_in_h[28] analog_io[28] mprj_pads.area2_io_pad\[9\]/PAD_A_ESD_1_H
+ gpio_dm2[28] gpio_dm1[28] gpio_dm0[28] gpio_in[28] gpio_inp_dis[28] gpio_ib_mode_sel[28]
+ porb_h porb_h mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD gpio_oeb[28] mprj_pads.area2_io_pad\[9\]/HLD_H_N
+ mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD gpio_slow_sel[28] gpio_vtrip_sel[28] gpio_holdover[28]
+ gpio_analog_en[28] gpio_analog_sel[28] gpio_loopback_one[28] mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD
+ gpio_analog_pol[28] gpio_out[28] vddio w_21151_664474# mprj_pads.area2_io_pad\[9\]/HLD_H_N
+ SUB w_21253_667565# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda2 w_23367_667565#
+ vddio SUB w_23367_664474# gpio[28] vccd sky130_ef_io__gpiov2_pad_wrapped
Xflash_io0_pad gpio_in_h[41] analog_io[41] flash_io0_pad/PAD_A_ESD_1_H gpio_dm2[41]
+ gpio_dm1[41] gpio_dm0[41] gpio_in[41] gpio_inp_dis[41] gpio_ib_mode_sel[41] porb_h
+ porb_h flash_io0_pad/TIE_LO_ESD gpio_oeb[41] flash_io0_pad/HLD_H_N flash_io0_pad/TIE_LO_ESD
+ gpio_slow_sel[41] gpio_vtrip_sel[41] gpio_holdover[41] gpio_analog_en[41] gpio_analog_sel[41]
+ gpio_loopback_one[41] flash_io0_pad/TIE_LO_ESD gpio_analog_pol[41] gpio_out[41]
+ vddio w_408069_21253# flash_io0_pad/HLD_H_N SUB w_404752_21253# vccd gpio_pad/AMUXBUS_B
+ gpio_pad/AMUXBUS_A vddio vdda w_404752_23367# vddio SUB w_408069_23367# gpio[41]
+ vccd sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vssa_hvclamp_pad\[0\] SUB vddio SUB SUB vccd vddio SUB vddio vdda1 vccd SUB
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[9\] gpio_in_h[9] analog_io[9] mprj_pads.area1_io_pad\[9\]/PAD_A_ESD_1_H
+ gpio_dm2[9] gpio_dm1[9] gpio_dm0[9] gpio_in[9] gpio_inp_dis[9] gpio_ib_mode_sel[9]
+ porb_h porb_h mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD gpio_oeb[9] mprj_pads.area1_io_pad\[9\]/HLD_H_N
+ mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD gpio_slow_sel[9] gpio_vtrip_sel[9] gpio_holdover[9]
+ gpio_analog_en[9] gpio_analog_sel[9] gpio_loopback_one[9] mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD
+ gpio_analog_pol[9] gpio_out[9] vddio w_694469_641469# mprj_pads.area1_io_pad\[9\]/HLD_H_N
+ SUB w_694469_638152# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_638152#
+ vddio SUB w_692253_641470# gpio[9] vccd sky130_ef_io__gpiov2_pad_wrapped
Xflash_clk_pad gpio_in_h[40] analog_io[40] flash_clk_pad/PAD_A_ESD_1_H gpio_dm2[40]
+ gpio_dm1[40] gpio_dm0[40] gpio_in[40] gpio_inp_dis[40] gpio_ib_mode_sel[40] porb_h
+ porb_h flash_clk_pad/TIE_LO_ESD gpio_oeb[40] flash_clk_pad/HLD_H_N flash_clk_pad/TIE_LO_ESD
+ gpio_slow_sel[40] gpio_vtrip_sel[40] gpio_holdover[40] gpio_analog_en[40] gpio_analog_sel[40]
+ gpio_loopback_one[40] flash_clk_pad/TIE_LO_ESD gpio_analog_pol[40] gpio_out[40]
+ vddio w_353269_21253# flash_clk_pad/HLD_H_N SUB w_349952_21253# vccd gpio_pad/AMUXBUS_B
+ gpio_pad/AMUXBUS_A vddio vdda w_349952_23367# vddio SUB w_353269_23367# gpio[39]
+ vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_0 gpio_loopback_zero[43] vccd gpio_loopback_one[43] SUB constant_block
Xuser1_vccd_lvclamp_pad vdda1 vccd vddio vddio gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A
+ vccd vccd1 vccd1 SUB SUB vddio SUB sky130_ef_io__vccd_lvc_clamped3_pad
Xmprj_pads.area1_io_pad\[13\] gpio_in_h[13] analog_io[13] mprj_pads.area1_io_pad\[13\]/PAD_A_ESD_1_H
+ gpio_dm2[13] gpio_dm1[13] gpio_dm0[13] gpio_in[13] gpio_inp_dis[13] gpio_ib_mode_sel[13]
+ porb_h porb_h mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD gpio_oeb[13] mprj_pads.area1_io_pad\[13\]/HLD_H_N
+ mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD gpio_slow_sel[13] gpio_vtrip_sel[13] gpio_holdover[13]
+ gpio_analog_en[13] gpio_analog_sel[13] gpio_loopback_one[13] mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD
+ gpio_analog_pol[13] gpio_out[13] vddio w_694469_865869# mprj_pads.area1_io_pad\[13\]/HLD_H_N
+ SUB w_694469_862552# vccd gpio_pad/AMUXBUS_B gpio_pad/AMUXBUS_A vddio vdda1 w_692355_862552#
+ vddio SUB w_692253_865870# gpio[13] vccd sky130_ef_io__gpiov2_pad_wrapped
Xconstant_block_1 gpio_loopback_zero[42] vccd gpio_loopback_one[42] SUB constant_block
.ends

.subckt caravel_openframe vddio_2 vssio vssd1 vdda vssa vccd vssd vdda1_2 vccd1 vccd2
+ gpio[0] gpio[1] gpio[2] gpio[3] gpio[4] gpio[5] gpio[6] gpio[7] gpio[8] gpio[9]
+ gpio[10] gpio[11] gpio[12] gpio[13] gpio[14] gpio[15] gpio[16] gpio[17] gpio[18]
+ gpio[19] gpio[20] gpio[21] gpio[22] gpio[23] gpio[24] gpio[25] gpio[26] gpio[27]
+ gpio[28] gpio[29] gpio[30] gpio[31] gpio[32] gpio[33] gpio[34] gpio[35] gpio[36]
+ gpio[37] gpio[38] gpio[39] gpio[40] gpio[41] gpio[42] gpio[43] resetb vdda2
Xchip_io_openframe_0 vddio_2 vssio vdda vccd2 vccd chip_io_openframe_0/vdda vdda1_2
+ vdda2 vccd1 resetb chip_io_openframe_0/porb_h chip_io_openframe_0/porb_l chip_io_openframe_0/por_l
+ chip_io_openframe_0/resetb_h chip_io_openframe_0/resetb_l chip_io_openframe_0/mask_rev[31]
+ chip_io_openframe_0/mask_rev[30] chip_io_openframe_0/mask_rev[29] chip_io_openframe_0/mask_rev[28]
+ chip_io_openframe_0/mask_rev[27] chip_io_openframe_0/mask_rev[26] chip_io_openframe_0/mask_rev[25]
+ chip_io_openframe_0/mask_rev[24] chip_io_openframe_0/mask_rev[23] chip_io_openframe_0/mask_rev[22]
+ chip_io_openframe_0/mask_rev[21] chip_io_openframe_0/mask_rev[20] chip_io_openframe_0/mask_rev[19]
+ chip_io_openframe_0/mask_rev[18] chip_io_openframe_0/mask_rev[17] chip_io_openframe_0/mask_rev[16]
+ chip_io_openframe_0/mask_rev[15] chip_io_openframe_0/mask_rev[14] chip_io_openframe_0/mask_rev[13]
+ chip_io_openframe_0/mask_rev[12] chip_io_openframe_0/mask_rev[11] chip_io_openframe_0/mask_rev[10]
+ chip_io_openframe_0/mask_rev[9] chip_io_openframe_0/mask_rev[8] chip_io_openframe_0/mask_rev[7]
+ chip_io_openframe_0/mask_rev[6] chip_io_openframe_0/mask_rev[5] chip_io_openframe_0/mask_rev[4]
+ chip_io_openframe_0/mask_rev[3] chip_io_openframe_0/mask_rev[2] chip_io_openframe_0/mask_rev[1]
+ chip_io_openframe_0/mask_rev[0] gpio[39] gpio[32] gpio[19] chip_io_openframe_0/gpio_out[43]
+ chip_io_openframe_0/gpio_out[40] chip_io_openframe_0/gpio_out[39] chip_io_openframe_0/gpio_out[38]
+ chip_io_openframe_0/gpio_out[37] chip_io_openframe_0/gpio_out[36] chip_io_openframe_0/gpio_out[28]
+ chip_io_openframe_0/gpio_out[27] chip_io_openframe_0/gpio_out[26] chip_io_openframe_0/gpio_out[25]
+ chip_io_openframe_0/gpio_out[19] chip_io_openframe_0/gpio_out[18] chip_io_openframe_0/gpio_out[17]
+ chip_io_openframe_0/gpio_out[16] chip_io_openframe_0/gpio_out[15] chip_io_openframe_0/gpio_out[14]
+ chip_io_openframe_0/gpio_out[13] chip_io_openframe_0/gpio_out[12] chip_io_openframe_0/gpio_out[11]
+ chip_io_openframe_0/gpio_out[10] chip_io_openframe_0/gpio_out[0] chip_io_openframe_0/gpio_oeb[43]
+ chip_io_openframe_0/gpio_oeb[42] chip_io_openframe_0/gpio_oeb[41] chip_io_openframe_0/gpio_oeb[40]
+ chip_io_openframe_0/gpio_oeb[39] chip_io_openframe_0/gpio_oeb[34] chip_io_openframe_0/gpio_oeb[33]
+ chip_io_openframe_0/gpio_oeb[29] chip_io_openframe_0/gpio_oeb[28] chip_io_openframe_0/gpio_oeb[27]
+ chip_io_openframe_0/gpio_oeb[26] chip_io_openframe_0/gpio_oeb[25] chip_io_openframe_0/gpio_oeb[23]
+ chip_io_openframe_0/gpio_oeb[22] chip_io_openframe_0/gpio_oeb[21] chip_io_openframe_0/gpio_oeb[20]
+ chip_io_openframe_0/gpio_oeb[17] chip_io_openframe_0/gpio_oeb[16] chip_io_openframe_0/gpio_oeb[11]
+ chip_io_openframe_0/gpio_oeb[7] chip_io_openframe_0/gpio_oeb[6] chip_io_openframe_0/gpio_oeb[1]
+ chip_io_openframe_0/gpio_inp_dis[39] chip_io_openframe_0/gpio_inp_dis[37] chip_io_openframe_0/gpio_inp_dis[35]
+ chip_io_openframe_0/gpio_inp_dis[34] chip_io_openframe_0/gpio_inp_dis[33] chip_io_openframe_0/gpio_inp_dis[30]
+ chip_io_openframe_0/gpio_inp_dis[29] chip_io_openframe_0/gpio_inp_dis[22] chip_io_openframe_0/gpio_inp_dis[21]
+ chip_io_openframe_0/gpio_inp_dis[20] chip_io_openframe_0/gpio_inp_dis[18] chip_io_openframe_0/gpio_inp_dis[17]
+ chip_io_openframe_0/gpio_inp_dis[16] chip_io_openframe_0/gpio_inp_dis[13] chip_io_openframe_0/gpio_inp_dis[12]
+ chip_io_openframe_0/gpio_inp_dis[9] chip_io_openframe_0/gpio_inp_dis[5] chip_io_openframe_0/gpio_inp_dis[1]
+ chip_io_openframe_0/gpio_ib_mode_sel[43] chip_io_openframe_0/gpio_ib_mode_sel[42]
+ chip_io_openframe_0/gpio_ib_mode_sel[41] chip_io_openframe_0/gpio_ib_mode_sel[40]
+ chip_io_openframe_0/gpio_ib_mode_sel[39] chip_io_openframe_0/gpio_ib_mode_sel[38]
+ chip_io_openframe_0/gpio_ib_mode_sel[37] chip_io_openframe_0/gpio_ib_mode_sel[34]
+ chip_io_openframe_0/gpio_ib_mode_sel[32] chip_io_openframe_0/gpio_ib_mode_sel[31]
+ chip_io_openframe_0/gpio_ib_mode_sel[26] chip_io_openframe_0/gpio_ib_mode_sel[25]
+ chip_io_openframe_0/gpio_ib_mode_sel[24] chip_io_openframe_0/gpio_ib_mode_sel[23]
+ chip_io_openframe_0/gpio_ib_mode_sel[22] chip_io_openframe_0/gpio_ib_mode_sel[21]
+ chip_io_openframe_0/gpio_ib_mode_sel[20] chip_io_openframe_0/gpio_ib_mode_sel[16]
+ chip_io_openframe_0/gpio_ib_mode_sel[13] chip_io_openframe_0/gpio_ib_mode_sel[10]
+ chip_io_openframe_0/gpio_ib_mode_sel[9] chip_io_openframe_0/gpio_ib_mode_sel[7]
+ chip_io_openframe_0/gpio_ib_mode_sel[4] chip_io_openframe_0/gpio_ib_mode_sel[1]
+ chip_io_openframe_0/gpio_vtrip_sel[43] chip_io_openframe_0/gpio_vtrip_sel[42] chip_io_openframe_0/gpio_vtrip_sel[37]
+ chip_io_openframe_0/gpio_vtrip_sel[36] chip_io_openframe_0/gpio_vtrip_sel[35] chip_io_openframe_0/gpio_vtrip_sel[28]
+ chip_io_openframe_0/gpio_vtrip_sel[27] chip_io_openframe_0/gpio_vtrip_sel[26] chip_io_openframe_0/gpio_vtrip_sel[25]
+ chip_io_openframe_0/gpio_vtrip_sel[24] chip_io_openframe_0/gpio_vtrip_sel[23] chip_io_openframe_0/gpio_vtrip_sel[22]
+ chip_io_openframe_0/gpio_vtrip_sel[19] chip_io_openframe_0/gpio_vtrip_sel[18] chip_io_openframe_0/gpio_vtrip_sel[17]
+ chip_io_openframe_0/gpio_vtrip_sel[16] chip_io_openframe_0/gpio_vtrip_sel[15] chip_io_openframe_0/gpio_vtrip_sel[14]
+ chip_io_openframe_0/gpio_vtrip_sel[13] chip_io_openframe_0/gpio_vtrip_sel[12] chip_io_openframe_0/gpio_vtrip_sel[11]
+ chip_io_openframe_0/gpio_vtrip_sel[10] chip_io_openframe_0/gpio_vtrip_sel[5] chip_io_openframe_0/gpio_vtrip_sel[4]
+ chip_io_openframe_0/gpio_vtrip_sel[3] chip_io_openframe_0/gpio_vtrip_sel[2] chip_io_openframe_0/gpio_vtrip_sel[1]
+ chip_io_openframe_0/gpio_vtrip_sel[0] chip_io_openframe_0/gpio_slow_sel[43] chip_io_openframe_0/gpio_slow_sel[34]
+ chip_io_openframe_0/gpio_slow_sel[32] chip_io_openframe_0/gpio_slow_sel[31] chip_io_openframe_0/gpio_slow_sel[30]
+ chip_io_openframe_0/gpio_slow_sel[28] chip_io_openframe_0/gpio_slow_sel[27] chip_io_openframe_0/gpio_slow_sel[26]
+ chip_io_openframe_0/gpio_slow_sel[22] chip_io_openframe_0/gpio_slow_sel[21] chip_io_openframe_0/gpio_slow_sel[17]
+ chip_io_openframe_0/gpio_slow_sel[15] chip_io_openframe_0/gpio_slow_sel[14] chip_io_openframe_0/gpio_slow_sel[13]
+ chip_io_openframe_0/gpio_slow_sel[12] chip_io_openframe_0/gpio_slow_sel[10] chip_io_openframe_0/gpio_slow_sel[9]
+ chip_io_openframe_0/gpio_slow_sel[8] chip_io_openframe_0/gpio_slow_sel[5] chip_io_openframe_0/gpio_slow_sel[4]
+ chip_io_openframe_0/gpio_slow_sel[0] chip_io_openframe_0/gpio_holdover[42] chip_io_openframe_0/gpio_holdover[41]
+ chip_io_openframe_0/gpio_holdover[37] chip_io_openframe_0/gpio_holdover[32] chip_io_openframe_0/gpio_holdover[31]
+ chip_io_openframe_0/gpio_holdover[30] chip_io_openframe_0/gpio_holdover[29] chip_io_openframe_0/gpio_holdover[26]
+ chip_io_openframe_0/gpio_holdover[25] chip_io_openframe_0/gpio_holdover[22] chip_io_openframe_0/gpio_holdover[21]
+ chip_io_openframe_0/gpio_holdover[15] chip_io_openframe_0/gpio_holdover[14] chip_io_openframe_0/gpio_holdover[13]
+ chip_io_openframe_0/gpio_holdover[12] chip_io_openframe_0/gpio_holdover[11] chip_io_openframe_0/gpio_holdover[10]
+ chip_io_openframe_0/gpio_holdover[9] chip_io_openframe_0/gpio_holdover[8] chip_io_openframe_0/gpio_holdover[7]
+ chip_io_openframe_0/gpio_holdover[6] chip_io_openframe_0/gpio_holdover[5] chip_io_openframe_0/gpio_holdover[3]
+ chip_io_openframe_0/gpio_holdover[2] chip_io_openframe_0/gpio_holdover[1] chip_io_openframe_0/gpio_analog_en[41]
+ chip_io_openframe_0/gpio_analog_en[40] chip_io_openframe_0/gpio_analog_en[38] chip_io_openframe_0/gpio_analog_en[37]
+ chip_io_openframe_0/gpio_analog_en[36] chip_io_openframe_0/gpio_analog_en[35] chip_io_openframe_0/gpio_analog_en[34]
+ chip_io_openframe_0/gpio_analog_en[33] chip_io_openframe_0/gpio_analog_en[32] chip_io_openframe_0/gpio_analog_en[31]
+ chip_io_openframe_0/gpio_analog_en[30] chip_io_openframe_0/gpio_analog_en[29] chip_io_openframe_0/gpio_analog_en[19]
+ chip_io_openframe_0/gpio_analog_en[18] chip_io_openframe_0/gpio_analog_en[17] chip_io_openframe_0/gpio_analog_en[16]
+ chip_io_openframe_0/gpio_analog_en[8] chip_io_openframe_0/gpio_analog_en[7] chip_io_openframe_0/gpio_analog_en[6]
+ chip_io_openframe_0/gpio_analog_en[5] chip_io_openframe_0/gpio_analog_en[4] chip_io_openframe_0/gpio_analog_en[3]
+ chip_io_openframe_0/gpio_analog_en[2] chip_io_openframe_0/gpio_analog_en[1] chip_io_openframe_0/gpio_analog_en[0]
+ chip_io_openframe_0/gpio_analog_sel[39] chip_io_openframe_0/gpio_analog_sel[38]
+ chip_io_openframe_0/gpio_analog_sel[36] chip_io_openframe_0/gpio_analog_sel[35]
+ chip_io_openframe_0/gpio_analog_sel[34] chip_io_openframe_0/gpio_analog_sel[31]
+ chip_io_openframe_0/gpio_analog_sel[30] chip_io_openframe_0/gpio_analog_sel[26]
+ chip_io_openframe_0/gpio_analog_sel[19] chip_io_openframe_0/gpio_analog_sel[18]
+ chip_io_openframe_0/gpio_analog_sel[16] chip_io_openframe_0/gpio_analog_sel[15]
+ chip_io_openframe_0/gpio_analog_sel[14] chip_io_openframe_0/gpio_analog_sel[11]
+ chip_io_openframe_0/gpio_analog_sel[10] chip_io_openframe_0/gpio_analog_sel[9] chip_io_openframe_0/gpio_analog_sel[8]
+ chip_io_openframe_0/gpio_analog_sel[5] chip_io_openframe_0/gpio_analog_sel[4] chip_io_openframe_0/gpio_analog_sel[0]
+ chip_io_openframe_0/gpio_analog_pol[43] chip_io_openframe_0/gpio_analog_pol[39]
+ chip_io_openframe_0/gpio_analog_pol[38] chip_io_openframe_0/gpio_analog_pol[37]
+ chip_io_openframe_0/gpio_analog_pol[34] chip_io_openframe_0/gpio_analog_pol[33]
+ chip_io_openframe_0/gpio_analog_pol[32] chip_io_openframe_0/gpio_analog_pol[29]
+ chip_io_openframe_0/gpio_analog_pol[25] chip_io_openframe_0/gpio_analog_pol[19]
+ chip_io_openframe_0/gpio_analog_pol[18] chip_io_openframe_0/gpio_analog_pol[17]
+ chip_io_openframe_0/gpio_analog_pol[14] chip_io_openframe_0/gpio_analog_pol[13]
+ chip_io_openframe_0/gpio_analog_pol[8] chip_io_openframe_0/gpio_analog_pol[7] chip_io_openframe_0/gpio_analog_pol[6]
+ chip_io_openframe_0/gpio_analog_pol[3] chip_io_openframe_0/gpio_analog_pol[2] chip_io_openframe_0/gpio_dm0[39]
+ chip_io_openframe_0/gpio_dm0[30] chip_io_openframe_0/gpio_dm0[28] chip_io_openframe_0/gpio_dm0[27]
+ chip_io_openframe_0/gpio_dm0[24] chip_io_openframe_0/gpio_dm0[23] chip_io_openframe_0/gpio_dm0[20]
+ chip_io_openframe_0/gpio_dm0[19] chip_io_openframe_0/gpio_dm0[13] chip_io_openframe_0/gpio_dm0[12]
+ chip_io_openframe_0/gpio_dm0[11] chip_io_openframe_0/gpio_dm0[10] chip_io_openframe_0/gpio_dm0[8]
+ chip_io_openframe_0/gpio_dm0[7] chip_io_openframe_0/gpio_dm0[3] chip_io_openframe_0/gpio_dm1[41]
+ chip_io_openframe_0/gpio_dm1[40] chip_io_openframe_0/gpio_dm1[39] chip_io_openframe_0/gpio_dm1[34]
+ chip_io_openframe_0/gpio_dm1[30] chip_io_openframe_0/gpio_dm1[29] chip_io_openframe_0/gpio_dm1[28]
+ chip_io_openframe_0/gpio_dm1[27] chip_io_openframe_0/gpio_dm1[26] chip_io_openframe_0/gpio_dm1[25]
+ chip_io_openframe_0/gpio_dm1[24] chip_io_openframe_0/gpio_dm1[23] chip_io_openframe_0/gpio_dm1[21]
+ chip_io_openframe_0/gpio_dm1[20] chip_io_openframe_0/gpio_dm1[19] chip_io_openframe_0/gpio_dm1[16]
+ chip_io_openframe_0/gpio_dm1[15] chip_io_openframe_0/gpio_dm1[11] chip_io_openframe_0/gpio_dm1[2]
+ chip_io_openframe_0/gpio_dm1[1] chip_io_openframe_0/gpio_dm1[0] chip_io_openframe_0/gpio_dm2[39]
+ chip_io_openframe_0/gpio_dm2[37] chip_io_openframe_0/gpio_dm2[35] chip_io_openframe_0/gpio_dm2[34]
+ chip_io_openframe_0/gpio_dm2[31] chip_io_openframe_0/gpio_dm2[30] chip_io_openframe_0/gpio_dm2[27]
+ chip_io_openframe_0/gpio_dm2[23] chip_io_openframe_0/gpio_dm2[19] chip_io_openframe_0/gpio_dm2[17]
+ chip_io_openframe_0/gpio_dm2[16] chip_io_openframe_0/gpio_dm2[15] chip_io_openframe_0/gpio_dm2[12]
+ chip_io_openframe_0/gpio_dm2[11] chip_io_openframe_0/gpio_dm2[9] chip_io_openframe_0/gpio_dm2[8]
+ chip_io_openframe_0/gpio_dm2[7] chip_io_openframe_0/gpio_dm2[6] chip_io_openframe_0/gpio_dm2[4]
+ chip_io_openframe_0/gpio_dm2[3] chip_io_openframe_0/gpio_dm2[0] chip_io_openframe_0/gpio_in[39]
+ chip_io_openframe_0/gpio_in[38] chip_io_openframe_0/gpio_in[37] chip_io_openframe_0/gpio_in[35]
+ chip_io_openframe_0/gpio_in[34] chip_io_openframe_0/gpio_in[33] chip_io_openframe_0/gpio_in[32]
+ chip_io_openframe_0/gpio_in[31] chip_io_openframe_0/gpio_in[30] chip_io_openframe_0/gpio_in[27]
+ chip_io_openframe_0/gpio_in[26] chip_io_openframe_0/gpio_in[23] chip_io_openframe_0/gpio_in[18]
+ chip_io_openframe_0/gpio_in[17] chip_io_openframe_0/gpio_in[16] chip_io_openframe_0/gpio_in[15]
+ chip_io_openframe_0/gpio_in[14] chip_io_openframe_0/gpio_in[12] chip_io_openframe_0/gpio_in[11]
+ chip_io_openframe_0/gpio_in[8] chip_io_openframe_0/gpio_in[5] chip_io_openframe_0/gpio_in_h[42]
+ chip_io_openframe_0/gpio_in_h[39] chip_io_openframe_0/gpio_in_h[37] chip_io_openframe_0/gpio_in_h[34]
+ chip_io_openframe_0/gpio_in_h[33] chip_io_openframe_0/gpio_in_h[32] chip_io_openframe_0/gpio_in_h[29]
+ chip_io_openframe_0/gpio_in_h[24] chip_io_openframe_0/gpio_in_h[20] chip_io_openframe_0/gpio_in_h[17]
+ chip_io_openframe_0/gpio_in_h[16] chip_io_openframe_0/gpio_in_h[15] chip_io_openframe_0/gpio_in_h[12]
+ chip_io_openframe_0/gpio_in_h[11] chip_io_openframe_0/gpio_in_h[10] chip_io_openframe_0/gpio_in_h[7]
+ chip_io_openframe_0/gpio_in_h[6] chip_io_openframe_0/gpio_in_h[2] chip_io_openframe_0/gpio_in_h[1]
+ chip_io_openframe_0/gpio_loopback_zero[43] chip_io_openframe_0/gpio_loopback_zero[42]
+ chip_io_openframe_0/gpio_loopback_zero[41] chip_io_openframe_0/gpio_loopback_zero[40]
+ chip_io_openframe_0/gpio_loopback_zero[39] chip_io_openframe_0/gpio_loopback_zero[38]
+ chip_io_openframe_0/gpio_loopback_one[43] chip_io_openframe_0/gpio_loopback_one[42]
+ chip_io_openframe_0/gpio_loopback_one[41] chip_io_openframe_0/gpio_loopback_one[40]
+ chip_io_openframe_0/gpio_loopback_one[39] chip_io_openframe_0/gpio_loopback_one[35]
+ chip_io_openframe_0/gpio_loopback_one[31] chip_io_openframe_0/gpio_loopback_one[29]
+ chip_io_openframe_0/gpio_loopback_one[28] chip_io_openframe_0/gpio_loopback_one[27]
+ chip_io_openframe_0/gpio_loopback_one[25] chip_io_openframe_0/gpio_loopback_one[24]
+ chip_io_openframe_0/gpio_loopback_one[23] chip_io_openframe_0/gpio_loopback_one[21]
+ chip_io_openframe_0/gpio_loopback_one[20] chip_io_openframe_0/gpio_loopback_one[17]
+ chip_io_openframe_0/gpio_loopback_one[13] chip_io_openframe_0/gpio_loopback_one[9]
+ chip_io_openframe_0/gpio_loopback_one[6] chip_io_openframe_0/analog_io[43] chip_io_openframe_0/analog_io[41]
+ chip_io_openframe_0/analog_io[39] chip_io_openframe_0/analog_io[38] chip_io_openframe_0/analog_io[35]
+ chip_io_openframe_0/analog_io[34] chip_io_openframe_0/analog_io[33] chip_io_openframe_0/analog_io[30]
+ chip_io_openframe_0/analog_io[24] chip_io_openframe_0/analog_io[20] chip_io_openframe_0/analog_io[19]
+ chip_io_openframe_0/analog_io[18] chip_io_openframe_0/analog_io[16] chip_io_openframe_0/analog_io[15]
+ chip_io_openframe_0/analog_io[14] chip_io_openframe_0/analog_io[10] chip_io_openframe_0/analog_io[9]
+ chip_io_openframe_0/analog_io[8] chip_io_openframe_0/analog_io[3] gpio[42] gpio[28]
+ gpio[27] gpio[26] gpio[25] gpio[23] gpio[1] gpio[0] chip_io_openframe_0/gpio_analog_pol[20]
+ w_694469_865869# w_23367_407274# w_694469_100152# w_23367_534874# w_137274_1012253#
+ chip_io_openframe_0/gpio_out[1] w_188674_1014469# chip_io_openframe_0/gpio_dm0[15]
+ w_404752_21253# w_459552_23367# w_485565_1014469# w_291674_1014469# w_638765_1014469#
+ w_23367_280765# chip_io_openframe_0/gpio_out[2] w_692253_776670# w_23367_710765#
+ chip_io_openframe_0/gpio_holdover[16] chip_io_openframe_0/gpio_inp_dis[25] w_692355_547952#
+ w_23367_537965# w_21151_364074# chip_io_openframe_0/gpio_holdover[33] w_21253_966965#
+ chip_io_openframe_0/gpio_out[3] w_694469_145352# w_459552_21253# w_692355_593152#
+ w_485565_1012355# w_694469_951752# w_694469_190352# w_638765_1012355# chip_io_openframe_0/gpio_analog_pol[41]
+ w_349952_23367# chip_io_openframe_0/gpio_analog_sel[40] chip_io_openframe_0/gpio_out[4]
+ w_692355_325552# w_189869_23367# chip_io_openframe_0/gpio_inp_dis[41] w_21151_794074#
+ w_694469_235552# w_692355_683352# chip_io_openframe_0/gpio_analog_sel[21] w_21253_194365#
+ w_694469_280552# w_85874_1014469# chip_io_openframe_0/gpio_out[5] chip_io_openframe_0/gpio_in_h[40]
+ chip_io_openframe_0/analog_io[40] chip_io_openframe_0/gpio_loopback_one[2] chip_io_openframe_0/gpio_inp_dis[42]
+ chip_io_openframe_0/gpio_dm0[34] w_21253_624365# w_482474_1012253# w_295152_23367#
+ w_635674_1012253# w_349952_21253# chip_io_openframe_0/gpio_in[20] chip_io_openframe_0/gpio_analog_pol[24]
+ w_23367_578074# w_692253_551270# chip_io_openframe_0/gpio_dm1[3] chip_io_openframe_0/gpio_out[6]
+ w_694469_370752# w_189869_21253# chip_io_openframe_0/gpio_dm1[7] chip_io_openframe_0/gpio_in_h[23]
+ chip_io_openframe_0/gpio_in[2] chip_io_openframe_0/gpio_out[7] chip_io_openframe_0/gpio_oeb[0]
+ chip_io_openframe_0/gpio_slow_sel[37] w_21151_277674# w_692253_641470# w_692253_955070#
+ chip_io_openframe_0/analog_io[23] w_295152_21253# w_294765_1014469# chip_io_openframe_0/gpio_inp_dis[6]
+ chip_io_openframe_0/gpio_analog_en[9] w_21151_707674# w_23367_234474# w_692355_100152#
+ w_694469_776669# chip_io_openframe_0/gpio_analog_en[20] chip_io_openframe_0/gpio_out[8]
+ w_393474_1014469# w_21151_963874# chip_io_openframe_0/gpio_ib_mode_sel[29] chip_io_openframe_0/gpio_holdover[39]
+ chip_io_openframe_0/gpio_inp_dis[2] chip_io_openframe_0/gpio_dm0[16] w_692253_596470#
+ chip_io_openframe_0/gpio_oeb[10] chip_io_openframe_0/gpio_ib_mode_sel[28] chip_io_openframe_0/gpio_dm1[12]
+ chip_io_openframe_0/gpio_analog_en[21] w_692253_731670# w_21253_280765# chip_io_openframe_0/analog_io[28]
+ chip_io_openframe_0/gpio_out[9] chip_io_openframe_0/analog_io[29] w_692253_328870#
+ chip_io_openframe_0/gpio_holdover[17] chip_io_openframe_0/gpio_analog_en[22] w_23367_410365#
+ w_21253_710765# chip_io_openframe_0/gpio_loopback_one[10] chip_io_openframe_0/gpio_inp_dis[26]
+ w_294765_1012355# chip_io_openframe_0/gpio_holdover[34] w_462869_23367# w_23367_237565#
+ chip_io_openframe_0/gpio_in_h[28] w_21253_537965# chip_io_openframe_0/gpio_dm2[20]
+ w_23367_664474# w_692253_686670# chip_io_openframe_0/gpio_analog_en[23] w_21151_191274#
+ chip_io_openframe_0/analog_io[2] chip_io_openframe_0/gpio_in_h[0] chip_io_openframe_0/gpio_analog_sel[25]
+ w_692253_374070# chip_io_openframe_0/gpio_oeb[5] chip_io_openframe_0/gpio_ib_mode_sel[11]
+ chip_io_openframe_0/gpio_dm2[24] w_21151_621274# w_692355_145352# chip_io_openframe_0/gpio_analog_en[24]
+ chip_io_openframe_0/gpio_analog_sel[20] chip_io_openframe_0/gpio_out[41] w_692355_951752#
+ w_692355_190352# w_694469_862552# chip_io_openframe_0/gpio_oeb[32] w_88965_1014469#
+ chip_io_openframe_0/gpio_analog_pol[28] chip_io_openframe_0/gpio_loopback_one[14]
+ chip_io_openframe_0/gpio_dm2[28] chip_io_openframe_0/gpio_analog_pol[42] chip_io_openframe_0/gpio_analog_en[25]
+ w_188674_1012253# chip_io_openframe_0/analog_io[7] chip_io_openframe_0/gpio_analog_pol[23]
+ chip_io_openframe_0/gpio_in[9] w_291674_1012253# chip_io_openframe_0/gpio_oeb[15]
+ w_462869_21253# w_23367_667565# chip_io_openframe_0/gpio_in_h[22] chip_io_openframe_0/gpio_dm0[0]
+ w_692355_235552# chip_io_openframe_0/gpio_analog_en[26] w_694469_551269# chip_io_openframe_0/gpio_dm0[31]
+ chip_io_openframe_0/gpio_vtrip_sel[39] w_23367_320874# chip_io_openframe_0/gpio_loopback_one[32]
+ w_692355_280552# chip_io_openframe_0/gpio_slow_sel[20] chip_io_openframe_0/gpio_slow_sel[36]
+ chip_io_openframe_0/gpio_in[24] chip_io_openframe_0/gpio_slow_sel[38] chip_io_openframe_0/gpio_dm0[4]
+ chip_io_openframe_0/gpio_analog_en[27] chip_io_openframe_0/gpio_dm0[35] chip_io_openframe_0/gpio_analog_en[42]
+ chip_io_openframe_0/gpio_dm1[31] chip_io_openframe_0/gpio_analog_sel[43] chip_io_openframe_0/gpio_loopback_one[3]
+ chip_io_openframe_0/gpio_analog_sel[3] chip_io_openframe_0/gpio_loopback_one[18]
+ chip_io_openframe_0/analog_io[22] w_88965_1012355# chip_io_openframe_0/gpio_ib_mode_sel[2]
+ chip_io_openframe_0/gpio_slow_sel[41] w_692253_103470# chip_io_openframe_0/gpio_in_h[5]
+ w_140365_1014469# chip_io_openframe_0/gpio_analog_en[28] w_694469_641469# w_694469_955069#
+ chip_io_openframe_0/gpio_dm1[4] chip_io_openframe_0/gpio_dm1[35] chip_io_openframe_0/gpio_ib_mode_sel[14]
+ w_692355_370752# chip_io_openframe_0/gpio_slow_sel[3] chip_io_openframe_0/gpio_in[6]
+ chip_io_openframe_0/gpio_analog_sel[41] chip_io_openframe_0/gpio_loopback_one[36]
+ w_23367_323965# w_23367_750874# chip_io_openframe_0/gpio_vtrip_sel[38] chip_io_openframe_0/gpio_dm1[8]
+ chip_io_openframe_0/gpio_oeb[37] w_396565_1014469# chip_io_openframe_0/gpio_analog_pol[1]
+ w_240074_1014469# chip_io_openframe_0/analog_io[27] chip_io_openframe_0/gpio_analog_en[43]
+ w_694469_596469# chip_io_openframe_0/gpio_ib_mode_sel[35] chip_io_openframe_0/gpio_inp_dis[7]
+ w_23367_581165# chip_io_openframe_0/gpio_loopback_one[7] chip_io_openframe_0/gpio_in[21]
+ w_694469_731669# chip_io_openframe_0/gpio_analog_pol[12] w_21151_407274# w_186552_23367#
+ chip_io_openframe_0/gpio_in_h[27] w_517669_23367# w_21151_534874# w_85874_1012253#
+ w_694469_328869# w_140365_1012355# chip_io_openframe_0/gpio_slow_sel[25] chip_io_openframe_0/gpio_oeb[4]
+ chip_io_openframe_0/gpio_inp_dis[3] chip_io_openframe_0/gpio_analog_sel[29] chip_io_openframe_0/analog_io[1]
+ chip_io_openframe_0/gpio_dm0[21] w_692253_148670# w_23367_753965# chip_io_openframe_0/gpio_in[3]
+ w_694469_686669# chip_io_openframe_0/gpio_dm0[17] w_692253_193670# chip_io_openframe_0/gpio_analog_sel[24]
+ chip_io_openframe_0/gpio_inp_dis[14] chip_io_openframe_0/gpio_dm1[13] chip_io_openframe_0/analog_io[13]
+ chip_io_openframe_0/gpio_in_h[43] chip_io_openframe_0/gpio_oeb[31] w_694469_374069#
+ chip_io_openframe_0/gpio_ib_mode_sel[5] chip_io_openframe_0/gpio_dm0[25] chip_io_openframe_0/gpio_holdover[18]
+ w_396565_1012355# chip_io_openframe_0/gpio_inp_dis[31] chip_io_openframe_0/gpio_inp_dis[27]
+ chip_io_openframe_0/gpio_ib_mode_sel[17] w_21253_410365# chip_io_openframe_0/gpio_holdover[35]
+ chip_io_openframe_0/gpio_dm1[17] w_694469_638152# chip_io_openframe_0/gpio_inp_dis[10]
+ chip_io_openframe_0/gpio_dm2[13] chip_io_openframe_0/gpio_oeb[14] chip_io_openframe_0/analog_io[6]
+ chip_io_openframe_0/gpio_analog_pol[27] chip_io_openframe_0/gpio_in_h[21] w_186552_21253#
+ w_517669_21253# chip_io_openframe_0/gpio_inp_dis[43] chip_io_openframe_0/gpio_loopback_one[11]
+ w_21253_237565# w_692253_238870# w_23367_364074# chip_io_openframe_0/gpio_dm0[40]
+ chip_io_openframe_0/gpio_inp_dis[23] chip_io_openframe_0/gpio_dm2[21] w_692253_283870#
+ chip_io_openframe_0/gpio_slow_sel[19] chip_io_openframe_0/gpio_slow_sel[35] w_533874_1014469#
+ chip_io_openframe_0/gpio_analog_pol[22] chip_io_openframe_0/gpio_in[42] chip_io_openframe_0/gpio_holdover[27]
+ chip_io_openframe_0/gpio_dm2[25] chip_io_openframe_0/gpio_out[42] chip_io_openframe_0/gpio_in[0]
+ chip_io_openframe_0/gpio_inp_dis[19] chip_io_openframe_0/gpio_slow_sel[18] w_694469_728352#
+ chip_io_openframe_0/gpio_holdover[43] chip_io_openframe_0/gpio_analog_sel[7] w_692355_862552#
+ chip_io_openframe_0/gpio_in_h[4] w_393474_1012253# chip_io_openframe_0/gpio_holdover[23]
+ w_694469_773352# chip_io_openframe_0/gpio_oeb[9] chip_io_openframe_0/analog_io[21]
+ chip_io_openframe_0/gpio_analog_sel[2] chip_io_openframe_0/gpio_loopback_one[0]
+ chip_io_openframe_0/gpio_slow_sel[2] chip_io_openframe_0/gpio_dm2[40] chip_io_openframe_0/gpio_loopback_one[15]
+ chip_io_openframe_0/gpio_ib_mode_sel[30] w_23367_367165# w_21253_667565# chip_io_openframe_0/gpio_in_h[31]
+ w_23367_794074# w_694469_103469# chip_io_openframe_0/gpio_holdover[19] chip_io_openframe_0/analog_io[42]
+ chip_io_openframe_0/gpio_dm0[41] chip_io_openframe_0/gpio_analog_sel[13] chip_io_openframe_0/gpio_in[28]
+ chip_io_openframe_0/gpio_oeb[36] chip_io_openframe_0/gpio_dm0[1] chip_io_openframe_0/gpio_dm0[32]
+ w_137274_1014469# w_353269_23367# chip_io_openframe_0/gpio_ib_mode_sel[8] chip_io_openframe_0/gpio_slow_sel[29]
+ chip_io_openframe_0/gpio_oeb[38] chip_io_openframe_0/gpio_analog_pol[5] chip_io_openframe_0/gpio_analog_en[10]
+ chip_io_openframe_0/gpio_loopback_one[33] chip_io_openframe_0/gpio_in_h[14] chip_io_openframe_0/gpio_dm0[5]
+ chip_io_openframe_0/analog_io[26] chip_io_openframe_0/gpio_dm0[36] chip_io_openframe_0/gpio_in_h[26]
+ chip_io_openframe_0/gpio_in[40] chip_io_openframe_0/gpio_dm1[32] chip_io_openframe_0/gpio_analog_pol[0]
+ w_21151_578074# chip_io_openframe_0/gpio_analog_pol[16] chip_io_openframe_0/gpio_analog_en[11]
+ chip_io_openframe_0/gpio_loopback_one[4] chip_io_openframe_0/gpio_slow_sel[24] chip_io_openframe_0/gpio_oeb[3]
+ w_243165_1014469# chip_io_openframe_0/gpio_dm0[9] chip_io_openframe_0/gpio_ib_mode_sel[0]
+ chip_io_openframe_0/gpio_analog_pol[11] chip_io_openframe_0/gpio_dm1[5] gpio[14]
+ gpio[8] chip_io_openframe_0/gpio_dm1[36] chip_io_openframe_0/gpio_dm2[41] chip_io_openframe_0/gpio_analog_sel[33]
+ chip_io_openframe_0/gpio_dm2[1] chip_io_openframe_0/gpio_dm2[32] w_23367_797165#
+ chip_io_openframe_0/gpio_analog_en[12] chip_io_openframe_0/analog_io[0] chip_io_openframe_0/gpio_ib_mode_sel[12]
+ w_21253_323965# chip_io_openframe_0/gpio_vtrip_sel[41] chip_io_openframe_0/gpio_oeb[30]
+ gpio[2] chip_io_openframe_0/gpio_analog_sel[28] w_353269_21253# chip_io_openframe_0/gpio_dm1[9]
+ chip_io_openframe_0/gpio_loopback_one[22] chip_io_openframe_0/gpio_in[25] chip_io_openframe_0/gpio_in_h[9]
+ chip_io_openframe_0/gpio_analog_sel[42] chip_io_openframe_0/gpio_loopback_one[37]
+ chip_io_openframe_0/analog_io[32] chip_io_openframe_0/gpio_dm2[5] chip_io_openframe_0/analog_io[12]
+ chip_io_openframe_0/gpio_inp_dis[8] chip_io_openframe_0/gpio_dm2[36] chip_io_openframe_0/gpio_analog_en[13]
+ chip_io_openframe_0/gpio_analog_en[39] w_23367_277674# w_694469_148669# chip_io_openframe_0/gpio_slow_sel[42]
+ chip_io_openframe_0/gpio_analog_pol[36] chip_io_openframe_0/gpio_slow_sel[7] chip_io_openframe_0/gpio_analog_sel[23]
+ chip_io_openframe_0/gpio_in[29] w_21253_581165# w_694469_193669# chip_io_openframe_0/gpio_oeb[13]
+ chip_io_openframe_0/gpio_ib_mode_sel[33] chip_io_openframe_0/gpio_in_h[36] w_23367_707674#
+ chip_io_openframe_0/gpio_analog_pol[40] chip_io_openframe_0/gpio_out[29] gpio[3]
+ chip_io_openframe_0/gpio_in[43] chip_io_openframe_0/gpio_analog_en[14] chip_io_openframe_0/gpio_loopback_one[8]
+ chip_io_openframe_0/gpio_analog_pol[31] w_21151_234474# chip_io_openframe_0/analog_io[5]
+ chip_io_openframe_0/gpio_inp_dis[4] chip_io_openframe_0/gpio_in_h[38] chip_io_openframe_0/gpio_inp_dis[36]
+ w_243165_1012355# chip_io_openframe_0/gpio_dm0[14] chip_io_openframe_0/gpio_in[7]
+ w_23367_963874# chip_io_openframe_0/gpio_in[41] chip_io_openframe_0/gpio_dm1[10]
+ chip_io_openframe_0/gpio_analog_pol[26] chip_io_openframe_0/gpio_analog_en[15] chip_io_openframe_0/analog_io[37]
+ chip_io_openframe_0/analog_io[17] chip_io_openframe_0/gpio_dm0[22] chip_io_openframe_0/gpio_inp_dis[15]
+ chip_io_openframe_0/gpio_in_h[41] w_694469_238869# gpio[10] w_21253_753965# chip_io_openframe_0/gpio_loopback_one[26]
+ chip_io_openframe_0/gpio_inp_dis[0] chip_io_openframe_0/gpio_out[30] chip_io_openframe_0/gpio_dm0[18]
+ w_694469_283869# chip_io_openframe_0/gpio_analog_pol[21] chip_io_openframe_0/gpio_inp_dis[32]
+ chip_io_openframe_0/gpio_dm1[14] w_692253_865870# chip_io_openframe_0/gpio_inp_dis[28]
+ chip_io_openframe_0/gpio_in_h[3] gpio[15] chip_io_openframe_0/gpio_dm2[10] chip_io_openframe_0/gpio_holdover[4]
+ chip_io_openframe_0/gpio_in[22] w_536965_1014469# chip_io_openframe_0/gpio_oeb[8]
+ chip_io_openframe_0/gpio_dm0[26] chip_io_openframe_0/gpio_holdover[36] chip_io_openframe_0/gpio_ib_mode_sel[3]
+ chip_io_openframe_0/gpio_dm1[22] w_298469_23367# chip_io_openframe_0/gpio_inp_dis[11]
+ w_191765_1014469# chip_io_openframe_0/gpio_slow_sel[1] w_694469_547952# w_482474_1014469#
+ chip_io_openframe_0/gpio_analog_sel[6] w_692355_638152# chip_io_openframe_0/gpio_slow_sel[40]
+ chip_io_openframe_0/gpio_dm1[18] w_635674_1014469# chip_io_openframe_0/gpio_ib_mode_sel[15]
+ chip_io_openframe_0/gpio_in_h[30] chip_io_openframe_0/gpio_inp_dis[38] chip_io_openframe_0/gpio_dm2[14]
+ chip_io_openframe_0/gpio_inp_dis[24] chip_io_openframe_0/gpio_out[20] chip_io_openframe_0/gpio_out[31]
+ w_21151_664474# chip_io_openframe_0/gpio_slow_sel[39] chip_io_openframe_0/gpio_holdover[0]
+ chip_io_openframe_0/gpio_oeb[19] chip_io_openframe_0/gpio_oeb[35] gpio[4] w_23367_191274#
+ w_23367_966965# chip_io_openframe_0/gpio_analog_sel[1] vssd chip_io_openframe_0/gpio_holdover[28]
+ chip_io_openframe_0/gpio_analog_sel[17] w_240074_1012253# chip_io_openframe_0/gpio_dm2[22]
+ w_408069_23367# chip_io_openframe_0/gpio_loopback_one[12] chip_io_openframe_0/gpio_in[4]
+ gpio[12] chip_io_openframe_0/gpio_vtrip_sel[6] chip_io_openframe_0/gpio_dm2[18]
+ w_694469_593152# chip_io_openframe_0/gpio_vtrip_sel[29] chip_io_openframe_0/gpio_in_h[13]
+ w_23367_621274# chip_io_openframe_0/gpio_analog_pol[9] chip_io_openframe_0/gpio_analog_sel[12]
+ gpio[35] chip_io_openframe_0/gpio_oeb[18] gpio[16] chip_io_openframe_0/gpio_ib_mode_sel[36]
+ chip_io_openframe_0/gpio_inp_dis[40] chip_io_openframe_0/gpio_in[13] chip_io_openframe_0/gpio_in_h[25]
+ chip_io_openframe_0/gpio_dm2[26] chip_io_openframe_0/gpio_out[21] chip_io_openframe_0/gpio_out[32]
+ chip_io_openframe_0/gpio_slow_sel[11] chip_io_openframe_0/gpio_holdover[38] chip_io_openframe_0/gpio_holdover[24]
+ chip_io_openframe_0/analog_io[25] w_692355_728352# chip_io_openframe_0/gpio_vtrip_sel[40]
+ chip_io_openframe_0/gpio_analog_pol[4] chip_io_openframe_0/gpio_vtrip_sel[7] chip_io_openframe_0/gpio_vtrip_sel[30]
+ w_514352_23367# chip_io_openframe_0/gpio_loopback_one[30] w_694469_325552# chip_io_openframe_0/gpio_dm0[43]
+ chip_io_openframe_0/gpio_slow_sel[23] w_536965_1012355# chip_io_openframe_0/gpio_oeb[2]
+ chip_io_openframe_0/gpio_in[19] w_692355_773352# gpio[31] gpio[41] w_298469_21253#
+ w_191765_1012355# chip_io_openframe_0/gpio_dm0[29] chip_io_openframe_0/gpio_analog_pol[15]
+ gpio[38] gpio[33] chip_io_openframe_0/gpio_analog_sel[37] chip_io_openframe_0/gpio_vtrip_sel[8]
+ chip_io_openframe_0/gpio_holdover[20] chip_io_openframe_0/gpio_dm0[42] gpio[20]
+ chip_io_openframe_0/gpio_vtrip_sel[31] gpio[13] w_694469_683352# w_21253_367165#
+ chip_io_openframe_0/gpio_out[22] chip_io_openframe_0/gpio_out[33] chip_io_openframe_0/gpio_dm1[38]
+ chip_io_openframe_0/gpio_loopback_one[1] chip_io_openframe_0/gpio_holdover[40] chip_io_openframe_0/xres_buf_0/VGND
+ w_23367_194365# w_21151_320874# chip_io_openframe_0/gpio_dm1[43] gpio[11] chip_io_openframe_0/gpio_in[36]
+ chip_io_openframe_0/gpio_loopback_one[16] gpio[21] chip_io_openframe_0/gpio_in_h[8]
+ chip_io_openframe_0/gpio_analog_pol[10] chip_io_openframe_0/gpio_dm0[2] chip_io_openframe_0/gpio_analog_sel[32]
+ w_408069_21253# chip_io_openframe_0/gpio_dm0[33] gpio[30] chip_io_openframe_0/gpio_vtrip_sel[9]
+ chip_io_openframe_0/gpio_ib_mode_sel[27] chip_io_openframe_0/gpio_vtrip_sel[32]
+ w_23367_624365# chip_io_openframe_0/gpio_ib_mode_sel[6] gpio[37] chip_io_openframe_0/gpio_in[1]
+ gpio[24] chip_io_openframe_0/gpio_slow_sel[6] chip_io_openframe_0/analog_io[31]
+ chip_io_openframe_0/gpio_dm1[42] gpio[6] chip_io_openframe_0/analog_io[11] chip_io_openframe_0/gpio_dm0[38]
+ chip_io_openframe_0/gpio_oeb[12] chip_io_openframe_0/gpio_dm2[43] chip_io_openframe_0/gpio_vtrip_sel[20]
+ chip_io_openframe_0/gpio_analog_sel[27] chip_io_openframe_0/gpio_loopback_one[19]
+ chip_io_openframe_0/gpio_in_h[19] gpio[5] gpio[29] chip_io_openframe_0/gpio_ib_mode_sel[18]
+ chip_io_openframe_0/gpio_in_h[35] chip_io_openframe_0/gpio_dm0[6] gpio[9] chip_io_openframe_0/gpio_out[23]
+ chip_io_openframe_0/gpio_out[34] chip_io_openframe_0/gpio_loopback_one[34] chip_io_openframe_0/gpio_in[10]
+ chip_io_openframe_0/gpio_dm0[37] chip_io_openframe_0/gpio_oeb[24] chip_io_openframe_0/gpio_vtrip_sel[33]
+ chip_io_openframe_0/gpio_dm1[33] chip_io_openframe_0/gpio_loopback_one[38] gpio[40]
+ chip_io_openframe_0/gpio_dm2[29] w_514352_21253# chip_io_openframe_0/gpio_analog_pol[35]
+ gpio[34] w_533874_1012253# gpio[36] chip_io_openframe_0/gpio_slow_sel[33] chip_io_openframe_0/gpio_analog_sel[22]
+ gpio[18] chip_io_openframe_0/gpio_dm2[42] chip_io_openframe_0/gpio_vtrip_sel[21]
+ chip_io_openframe_0/analog_io[4] chip_io_openframe_0/gpio_dm2[38] w_404752_23367#
+ chip_io_openframe_0/gpio_in_h[18] chip_io_openframe_0/gpio_ib_mode_sel[19] chip_io_openframe_0/gpio_dm1[6]
+ chip_io_openframe_0/gpio_loopback_one[5] gpio[43] gpio[7] chip_io_openframe_0/gpio_analog_pol[30]
+ chip_io_openframe_0/gpio_vtrip_sel[34] chip_io_openframe_0/gpio_dm1[37] vssa chip_io_openframe_0/gpio_dm2[2]
+ w_21253_797165# chip_io_openframe_0/gpio_dm2[33] w_21151_750874# chip_io_openframe_0/gpio_out[24]
+ gpio[17] chip_io_openframe_0/gpio_out[35] chip_io_openframe_0/analog_io[36] gpio[22]
+ chip_io_openframe_0/gpio_slow_sel[16] vssd1 chip_io_openframe
.ends

