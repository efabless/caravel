module gpio_defaults_block (VPWR,
    VGND,
    gpio_defaults);
 input VPWR;
 input VGND;
 output [12:0] gpio_defaults;

 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_low[1] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;

 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign gpio_defaults[10] = \gpio_defaults_high[10] ;
 assign gpio_defaults[1] = \gpio_defaults_high[1] ;
 assign gpio_defaults[0] = \gpio_defaults_low[0] ;
 assign gpio_defaults[11] = \gpio_defaults_low[11] ;
 assign gpio_defaults[12] = \gpio_defaults_low[12] ;
 assign gpio_defaults[2] = \gpio_defaults_low[2] ;
 assign gpio_defaults[3] = \gpio_defaults_low[3] ;
 assign gpio_defaults[4] = \gpio_defaults_low[4] ;
 assign gpio_defaults[5] = \gpio_defaults_low[5] ;
 assign gpio_defaults[6] = \gpio_defaults_low[6] ;
 assign gpio_defaults[7] = \gpio_defaults_low[7] ;
 assign gpio_defaults[8] = \gpio_defaults_low[8] ;
 assign gpio_defaults[9] = \gpio_defaults_low[9] ;
endmodule
