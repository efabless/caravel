magic
tech sky130A
magscale 1 2
timestamp 1665519328
<< fillblock >>
rect -262 -266 35048 2764
rect -140 -5140 37048 -1424
rect 26 -10348 17310 -5358
use font_2E  font_2E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786878
transform 1 0 13680 0 1 0
box 0 0 720 720
use font_6B  font_6B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766293
transform 1 0 11520 0 1 -4000
box 0 0 1080 2520
use font_4B  font_4B_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766293
transform 1 0 34200 0 1 -4000
box 0 0 1080 2520
use font_6C  font_6C_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766404
transform 1 0 5760 0 1 -4000
box 0 0 1080 2520
use font_6E  font_6E_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598766739
transform 1 0 28080 0 1 -4000
box 0 0 1440 2520
use font_6F  font_6F_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598767855
transform 1 0 1440 0 1 -4000
box 0 0 1080 2520
use font_6F  font_6F_1
timestamp 1598767855
transform 1 0 2880 0 1 -4000
box 0 0 1080 2520
use font_6F  font_6F_2
timestamp 1598767855
transform 1 0 23760 0 1 -4000
box 0 0 1080 2520
use font_6C  font_6C_1
timestamp 1598776550
transform 1 0 8640 0 1 0
box 0 0 360 2520
use font_6C  font_6C_2
timestamp 1598776550
transform 1 0 28440 0 1 0
box 0 0 360 2520
use font_6C  font_6C_3
timestamp 1598776550
transform 1 0 5400 0 1 -8000
box 0 0 360 2520
use font_20  font_20_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598785497
transform 1 0 9360 0 1 0
box 0 0 1 1
use font_20  font_20_1
timestamp 1598785497
transform 1 0 16200 0 1 0
box 0 0 1 1
use font_20  font_20_2
timestamp 1598785497
transform 1 0 21240 0 1 0
box 0 0 1 1
use font_20  font_20_3
timestamp 1598785497
transform 1 0 33480 0 1 0
box 0 0 1 1
use font_20  font_20_4
timestamp 1598785497
transform 1 0 22320 0 1 -4000
box 0 0 1 1
use font_20  font_20_5
timestamp 1598785497
transform 1 0 29880 0 1 -4000
box 0 0 1 1
use font_20  font_20_6
timestamp 1598785497
transform 1 0 35640 0 1 -4000
box 0 0 1 1
use font_20  font_20_7
timestamp 1598785497
transform 1 0 6120 0 1 -8000
box 0 0 1 1
use font_28  font_28_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1606780629
transform 1 0 17640 0 1 0
box 0 0 720 2520
use font_29  font_29_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786350
transform 1 0 20160 0 1 0
box 0 0 720 2520
use font_30  font_30_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598786981
transform 1 0 14760 0 1 0
box 0 0 1080 2520
use font_30  font_30_1
timestamp 1598786981
transform 1 0 9000 0 1 -8000
box 0 0 1080 2520
use font_32  font_32_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787041
transform 1 0 7560 0 1 -8000
box 0 0 1080 2520
use font_32  font_32_1
timestamp 1598787041
transform 1 0 10440 0 1 -8000
box 0 0 1080 2520
use font_33  font_33_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787077
transform 1 0 11880 0 1 -8000
box 0 0 1080 2520
use font_36  font_36_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598787225
transform 1 0 12240 0 1 0
box 0 0 1080 2520
use font_61  font_61_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763107
transform 1 0 16560 0 1 -4000
box 0 0 1080 2520
use font_41  font_41_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763107
transform 1 0 0 0 1 -8000
box 0 0 1080 2520
use font_43  font_43_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763351
transform 1 0 0 0 1 0
box 0 0 1080 2520
use font_43  font_43_1
timestamp 1598763351
transform 1 0 18720 0 1 0
box 0 0 1080 2520
use font_44  font_44_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598763661
transform 1 0 32760 0 1 -4000
box 0 0 1080 2520
use font_65  font_65_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765099
transform 1 0 6500 0 1 -4000
box 0 0 1080 2520
use font_65  font_65_1
timestamp 1598765099
transform 1 0 19440 0 1 -4000
box 0 0 1080 2520
use font_65  font_65_2
timestamp 1598765099
transform 1 0 26640 0 1 -4000
box 0 0 1080 2520
use font_47  font_47_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765398
transform 1 0 0 0 1 -4000
box 0 0 1080 2520
use font_67  font_67_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598765398
transform 1 0 4320 0 1 -4000
box 0 0 1080 2520
use font_70  font_70_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 25200 0 1 -4000
box 0 0 1080 2520
use font_50  font_50_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768087
transform 1 0 31320 0 1 -4000
box 0 0 1080 2520
use font_70  font_70_1
timestamp 1598768087
transform 1 0 1440 0 1 -8000
box 0 0 1080 2520
use font_2D  font_2D_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768325
transform 1 0 8140 0 1 -4000
box 0 0 1080 2520
use font_72  font_72_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768719
transform 1 0 20880 0 1 -4000
box 0 0 1080 2520
use font_53  font_53_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768855
transform 1 0 10080 0 1 -4000
box 0 0 1080 2520
use font_74  font_74_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598768910
transform 1 0 18000 0 1 -4000
box 0 0 1080 2520
use font_56  font_56_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769117
transform 1 0 10800 0 1 0
box 0 0 1080 2520
use font_57  font_57_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769216
transform 1 0 14400 0 1 -4000
box 0 0 1800 2520
use font_79  font_79_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598769811
transform 1 0 12960 0 1 -4000
box 0 0 1080 2520
use font_61  font_61_1
timestamp 1598775307
transform 1 0 1440 0 1 0
box 0 0 1080 1800
use font_61  font_61_2
timestamp 1598775307
transform 1 0 4320 0 1 0
box 0 0 1080 1800
use font_61  font_61_3
timestamp 1598775307
transform 1 0 25560 0 1 0
box 0 0 1080 1800
use font_62  font_62_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775406
transform 1 0 27000 0 1 0
box 0 0 1080 2520
use font_65  font_65_3
timestamp 1598775915
transform 1 0 7200 0 1 0
box 0 0 1080 1800
use font_65  font_65_4
timestamp 1598775915
transform 1 0 22680 0 1 0
box 0 0 1080 1800
use font_65  font_65_5
timestamp 1598775915
transform 1 0 29160 0 1 0
box 0 0 1080 1800
use font_66  font_66_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598775974
transform 1 0 24120 0 1 0
box 0 0 1080 2520
use font_69  font_69_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598776260
transform 1 0 4320 0 1 -8000
box 0 0 720 2520
use font_72  font_72_1
timestamp 1598777237
transform 1 0 2880 0 1 0
box 0 0 1080 1800
use font_72  font_72_2
timestamp 1598777237
transform 1 0 2880 0 1 -8000
box 0 0 1080 1800
use font_73  font_73_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777283
transform 1 0 30600 0 1 0
box 0 0 1080 1800
use font_73  font_73_1
timestamp 1598777283
transform 1 0 32040 0 1 0
box 0 0 1080 1800
use font_76  font_76_0 $PDKPATH/libs.ref/sky130_ml_xx_hd/mag
timestamp 1598777472
transform 1 0 5760 0 1 0
box 0 0 1080 1800
<< end >>
