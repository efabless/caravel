* NGSPICE file created from housekeeping_alt.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_2 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_1 abstract view
.subckt sky130_fd_sc_hd__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_4 abstract view
.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping_alt VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0]
+ irq[1] irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_79_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3691__A2 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__A1 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6914_ _7264_/CLK _6914_/D fanout690/X VGND VGND VPWR VPWR _6914_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_70_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6845_ _6869_/A _6872_/B VGND VGND VPWR VPWR _6845_/X sky130_fd_sc_hd__and2_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6776_ _6930_/Q _6776_/A2 _6774_/Y _6775_/X VGND VGND VPWR VPWR _6776_/X sky130_fd_sc_hd__a22o_1
XFILLER_167_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3988_ _3988_/A _3988_/B _3988_/C _3988_/D VGND VGND VPWR VPWR _3995_/C sky130_fd_sc_hd__nor4_1
XANTENNA_fanout427_A _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5727_ _5727_/A0 _5952_/A1 _5730_/S VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3746__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6145__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5658_ _5955_/A1 _5658_/A1 _5658_/S VGND VGND VPWR VPWR _5658_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4156__A0 _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4609_ _4879_/D _4747_/B _4887_/B _4945_/A _4772_/B VGND VGND VPWR VPWR _4909_/A
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__6696__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5589_ _5589_/A0 _5645_/A0 _5589_/S VGND VGND VPWR VPWR _5589_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5705__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold340 _6900_/Q VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7328_ _7329_/CLK _7328_/D fanout704/X VGND VGND VPWR VPWR _7328_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_104_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold351 hold351/A VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold362 hold362/A VGND VGND VPWR VPWR _7328_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold373 hold373/A VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold384 hold384/A VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7259_ _7578_/CLK _7259_/D fanout745/X VGND VGND VPWR VPWR _7259_/Q sky130_fd_sc_hd__dfrtp_4
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5656__A0 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1611_A _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5120__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4845__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1040 _5786_/X VGND VGND VPWR VPWR _7391_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1051 hold3077/X VGND VGND VPWR VPWR hold3078/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1062 hold2967/X VGND VGND VPWR VPWR hold1062/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input127_A wb_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1073 hold1073/A VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1084 hold2972/X VGND VGND VPWR VPWR hold2973/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5959__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 hold3167/X VGND VGND VPWR VPWR _7559_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6620__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A3 _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4580__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_38_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5187__A2 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input92_A spimemio_flash_io3_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6687__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5895__A0 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6439__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5647__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7201__RESET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4905__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6611__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4960_ _4960_/A _4960_/B VGND VGND VPWR VPWR _5252_/B sky130_fd_sc_hd__nor2_1
X_3911_ _6912_/Q _5612_/B _5947_/A _3657_/X _6958_/Q VGND VGND VPWR VPWR _3911_/X
+ sky130_fd_sc_hd__a32o_4
X_4891_ _5222_/B _5222_/C _4970_/C _4891_/D VGND VGND VPWR VPWR _4891_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3976__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6630_ _7574_/Q _6424_/X _6628_/X _6629_/X VGND VGND VPWR VPWR _6630_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5178__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3842_ _7505_/Q _5983_/A _4376_/B _3841_/X VGND VGND VPWR VPWR _3842_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5032__D1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4386__A0 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6561_ _7371_/Q _6561_/A2 _6769_/A3 _6468_/X _7411_/Q VGND VGND VPWR VPWR _6561_/X
+ sky130_fd_sc_hd__a32o_1
X_3773_ _7490_/Q _5893_/A _3765_/X _3772_/X VGND VGND VPWR VPWR _3773_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3728__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5512_ _5512_/A _5575_/A _5548_/A _5512_/D VGND VGND VPWR VPWR _5512_/Y sky130_fd_sc_hd__nand4_1
XFILLER_157_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6127__A1 _7496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6492_ _7312_/Q _6419_/D _6452_/X _7344_/Q VGND VGND VPWR VPWR _6492_/X sky130_fd_sc_hd__a22o_1
XFILLER_145_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6678__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5443_ _4601_/Y _4956_/B _4659_/Y VGND VGND VPWR VPWR _5541_/D sky130_fd_sc_hd__a21o_1
X_5374_ _5480_/A1 _4846_/Y _4428_/B _5373_/X VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3553__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7113_ _7186_/CLK _7113_/D fanout725/X VGND VGND VPWR VPWR _7113_/Q sky130_fd_sc_hd__dfrtp_4
X_4325_ _4548_/A0 _4325_/A1 _4327_/S VGND VGND VPWR VPWR _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5638__A0 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7044_ _7201_/CLK _7044_/D fanout726/X VGND VGND VPWR VPWR _7044_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4256_ _4256_/A0 _5998_/A1 _4258_/S VGND VGND VPWR VPWR _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4187_ _4187_/A0 _7640_/Q _4429_/B VGND VGND VPWR VPWR _4187_/X sky130_fd_sc_hd__mux2_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6063__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6602__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout544_A _4447_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3967__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6828_ _6828_/A1 _7107_/Q _6798_/C VGND VGND VPWR VPWR _6828_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5169__A2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6366__A1 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4831__C _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3719__A3 _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6759_ _7015_/Q _4105_/B _6459_/B _6467_/X _7156_/Q VGND VGND VPWR VPWR _6759_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_183_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6669__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6120__A _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold170 hold170/A VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold192 hold192/A VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout661 fanout661/A VGND VGND VPWR VPWR _5107_/C sky130_fd_sc_hd__buf_6
XANTENNA__4301__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout672 _5134_/A VGND VGND VPWR VPWR _5059_/A sky130_fd_sc_hd__buf_6
XANTENNA__4575__A _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout683 _4840_/D VGND VGND VPWR VPWR _4747_/B sky130_fd_sc_hd__buf_12
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout694 fanout750/X VGND VGND VPWR VPWR fanout694/X sky130_fd_sc_hd__buf_6
XANTENNA__4852__A1 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A3 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3591__A1 input59/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3654__A _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3894__A2 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4110_ _4427_/C _4084_/X _4425_/B VGND VGND VPWR VPWR _7110_/D sky130_fd_sc_hd__a21o_1
XFILLER_96_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5090_ _4774_/Y _4960_/A _5089_/Y _5088_/Y VGND VGND VPWR VPWR _5090_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_150_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1809 _7520_/Q VGND VGND VPWR VPWR hold395/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6293__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4041_ _4041_/A1 _4040_/D _4040_/A _4044_/A1 VGND VGND VPWR VPWR _4042_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__4485__A _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5992_ _5992_/A hold40/X _5992_/C _5992_/D VGND VGND VPWR VPWR _6000_/S sky130_fd_sc_hd__and4_4
X_4943_ _5248_/B _4943_/B VGND VGND VPWR VPWR _4944_/C sky130_fd_sc_hd__nand2_1
XFILLER_178_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3949__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4932__B _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7662_ _7662_/A VGND VGND VPWR VPWR _7662_/X sky130_fd_sc_hd__clkbuf_2
X_4874_ _4984_/B _4984_/A _4668_/C _5100_/A VGND VGND VPWR VPWR _5203_/B sky130_fd_sc_hd__a2bb2o_2
X_6613_ _7317_/Q _6419_/D _6424_/X _7573_/Q _6612_/X VGND VGND VPWR VPWR _6613_/X
+ sky130_fd_sc_hd__a221o_1
X_3825_ _7174_/Q _3931_/B _4364_/B _5581_/A _7211_/Q VGND VGND VPWR VPWR _3825_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7593_ _7594_/CLK _7593_/D fanout692/X VGND VGND VPWR VPWR _7593_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_137_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6544_ _6544_/A _6544_/B _6544_/C _6544_/D VGND VGND VPWR VPWR _6545_/C sky130_fd_sc_hd__nor4_2
XFILLER_146_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3756_ _7554_/Q _3508_/X _4422_/S input46/X _3755_/X VGND VGND VPWR VPWR _3759_/C
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_5_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_5_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_134_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6475_ _7448_/Q _6467_/A _6574_/C _6408_/B _7376_/Q VGND VGND VPWR VPWR _6475_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5859__A0 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3687_ _7176_/Q _5866_/B _3576_/X _3537_/X _7427_/Q VGND VGND VPWR VPWR _3687_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3564__A _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5426_ _5158_/A _5342_/B _5038_/B _5339_/A VGND VGND VPWR VPWR _5426_/X sky130_fd_sc_hd__o211a_1
Xoutput220 _7658_/X VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
XANTENNA__5323__A2 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput231 _7668_/X VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput242 _7652_/X VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
Xoutput253 _4132_/A VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
Xoutput264 _7228_/Q VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
X_5357_ _4870_/A _4907_/B _5346_/X _5102_/B wire658/X VGND VGND VPWR VPWR _5357_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout494_A _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput275 _6918_/Q VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
Xoutput286 _6928_/Q VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XANTENNA__3885__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput297 _7246_/Q VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_99_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4308_ _4308_/A0 _5736_/A1 _4308_/S VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5288_ _4847_/X _5061_/X _5286_/X _5123_/X VGND VGND VPWR VPWR _5288_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_141_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7027_ _7035_/CLK _7027_/D fanout723/X VGND VGND VPWR VPWR _7027_/Q sky130_fd_sc_hd__dfrtp_4
X_4239_ _4239_/A0 _4238_/X _4249_/S VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5938__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire347 _3810_/Y VGND VGND VPWR VPWR _3855_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input55_A mgmt_gpio_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3876__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5078__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3628__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout480 _6561_/A2 VGND VGND VPWR VPWR _6459_/B sky130_fd_sc_hd__buf_8
XANTENNA__4736__C _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout491 _6447_/C VGND VGND VPWR VPWR _6600_/B sky130_fd_sc_hd__buf_6
XFILLER_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4455__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__A _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4244__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3610_ _7356_/Q _5803_/A hold90/A _3494_/X _7476_/Q VGND VGND VPWR VPWR _3610_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_80_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4590_ _4674_/A _4825_/A VGND VGND VPWR VPWR _4591_/B sky130_fd_sc_hd__and2b_4
XANTENNA__6750__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3541_ _5938_/B _3860_/D VGND VGND VPWR VPWR _3541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold906 _5792_/X VGND VGND VPWR VPWR _7397_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold917 hold917/A VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold928 hold928/A VGND VGND VPWR VPWR _7357_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold939 hold939/A VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6260_ _6649_/S _6260_/A2 _6258_/X _6259_/X _6573_/S VGND VGND VPWR VPWR _6260_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4108__A3 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3472_ _4551_/A _3507_/A _3576_/C VGND VGND VPWR VPWR _3472_/X sky130_fd_sc_hd__and3_2
XFILLER_170_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5211_ _4716_/Y _4886_/Y _4906_/B VGND VGND VPWR VPWR _5224_/A sky130_fd_sc_hd__o21ai_1
Xhold3008 _5957_/X VGND VGND VPWR VPWR hold3008/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6191_ _6649_/S _7604_/Q _6573_/S _6190_/X VGND VGND VPWR VPWR _6191_/X sky130_fd_sc_hd__a211o_1
Xhold3019 _7455_/Q VGND VGND VPWR VPWR hold3019/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_1_1__f_user_clock clkbuf_0_user_clock/X VGND VGND VPWR VPWR _4161_/A1 sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_7_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3867__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2307 hold593/X VGND VGND VPWR VPWR _5608_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5142_ _4956_/A _4690_/Y _4713_/X _4720_/Y _4706_/Y VGND VGND VPWR VPWR _5143_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2318 _7501_/Q VGND VGND VPWR VPWR hold747/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2329 _7310_/Q VGND VGND VPWR VPWR hold603/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1606 _5607_/X VGND VGND VPWR VPWR hold129/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1617 _5982_/X VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4419__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1628 _6905_/Q VGND VGND VPWR VPWR _4028_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5073_ _5073_/A _5073_/B VGND VGND VPWR VPWR _5081_/A sky130_fd_sc_hd__nand2_8
Xhold1639 hold163/X VGND VGND VPWR VPWR _7469_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4024_ _4024_/A1 _4040_/A _4023_/X VGND VGND VPWR VPWR _6906_/D sky130_fd_sc_hd__o21a_1
XANTENNA__3550__C _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4292__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4943__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5758__B hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5975_ _5975_/A0 _5975_/A1 _5982_/S VGND VGND VPWR VPWR _5975_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4154__S _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4926_ _4997_/B _4954_/C _4933_/A _5260_/D VGND VGND VPWR VPWR _4927_/B sky130_fd_sc_hd__and4_1
XFILLER_33_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4857_ _4856_/A _5072_/B _5058_/D VGND VGND VPWR VPWR _4857_/X sky130_fd_sc_hd__and3b_4
X_7645_ _4164_/A1 _7645_/D fanout751/X VGND VGND VPWR VPWR _7645_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3808_ _7305_/Q _5686_/A _5704_/A _7321_/Q _3807_/X VGND VGND VPWR VPWR _3808_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7576_ _7576_/CLK _7576_/D fanout718/X VGND VGND VPWR VPWR _7576_/Q sky130_fd_sc_hd__dfstp_2
X_4788_ _4790_/C _5089_/B _4788_/C VGND VGND VPWR VPWR _5096_/A sky130_fd_sc_hd__and3_4
XANTENNA__5544__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6741__B2 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6527_ _7370_/Q _6561_/A2 _6769_/A3 _6455_/X _7458_/Q VGND VGND VPWR VPWR _6527_/X
+ sky130_fd_sc_hd__a32o_1
X_3739_ _7290_/Q _5956_/B _4352_/A _4322_/A _7004_/Q VGND VGND VPWR VPWR _3739_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6458_ _7431_/Q _6747_/B _6747_/C _6457_/X _7471_/Q VGND VGND VPWR VPWR _6458_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5409_ _4687_/Y _5406_/Y _4761_/Y _5140_/X _5303_/D VGND VGND VPWR VPWR _5569_/A
+ sky130_fd_sc_hd__o311a_1
X_6389_ _7030_/Q _6099_/X _6111_/X _7040_/Q _6388_/X VGND VGND VPWR VPWR _6389_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_133_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2830 _7654_/A VGND VGND VPWR VPWR hold2830/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2841 _5815_/X VGND VGND VPWR VPWR hold2841/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2852 _4349_/X VGND VGND VPWR VPWR hold2852/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2863 _7237_/Q VGND VGND VPWR VPWR hold2863/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2874 _7482_/Q VGND VGND VPWR VPWR hold2874/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2885 hold2885/A VGND VGND VPWR VPWR _5599_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2896 _5861_/X VGND VGND VPWR VPWR hold2896/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5480__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5480__B2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3491__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5668__B _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5232__A1 _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3546__A1 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3546__B2 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A2 _3549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4747__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6248__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3651__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4239__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6799__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6799__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6263__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4663__B1_N _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5471__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5760_ _5994_/A1 _5760_/A1 hold27/X VGND VGND VPWR VPWR _5760_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ _4753_/C _4767_/B VGND VGND VPWR VPWR _5404_/B sky130_fd_sc_hd__and2_2
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5691_ _5952_/A1 _5691_/A1 _5694_/S VGND VGND VPWR VPWR _5691_/X sky130_fd_sc_hd__mux2_1
X_7430_ _7579_/CLK hold34/X fanout731/X VGND VGND VPWR VPWR _7430_/Q sky130_fd_sc_hd__dfrtp_4
X_4642_ _4675_/A _4675_/B _4643_/C _4645_/D VGND VGND VPWR VPWR _4648_/A sky130_fd_sc_hd__nand4_4
XFILLER_147_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7361_ _7537_/CLK _7361_/D fanout707/X VGND VGND VPWR VPWR _7361_/Q sky130_fd_sc_hd__dfrtp_4
X_4573_ _5058_/D _4888_/B _4888_/C VGND VGND VPWR VPWR _4667_/B sky130_fd_sc_hd__nand3_4
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold703 hold703/A VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold714 _5757_/X VGND VGND VPWR VPWR _7366_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6312_ _7042_/Q _6089_/X _6308_/X _6309_/X _6311_/X VGND VGND VPWR VPWR _6312_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3545__C _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3524_ _3524_/A _3524_/B _3524_/C _3524_/D VGND VGND VPWR VPWR _3570_/B sky130_fd_sc_hd__nor4_2
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7292_ _7334_/CLK _7292_/D fanout710/X VGND VGND VPWR VPWR _7292_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold736 hold736/A VGND VGND VPWR VPWR _7010_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold747 hold747/A VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold758 _5592_/X VGND VGND VPWR VPWR _7225_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6487__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6243_ _7381_/Q _6089_/X _6239_/X _6240_/X _6242_/X VGND VGND VPWR VPWR _6243_/X
+ sky130_fd_sc_hd__a2111o_1
X_3455_ _6904_/Q hold246/X _4007_/B VGND VGND VPWR VPWR _3455_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6174_ _7378_/Q _6089_/X _6144_/C _6173_/X VGND VGND VPWR VPWR _6174_/X sky130_fd_sc_hd__a31o_1
Xhold2104 _4220_/X VGND VGND VPWR VPWR hold530/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2115 _7188_/Q VGND VGND VPWR VPWR hold322/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2126 hold477/X VGND VGND VPWR VPWR _4232_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3561__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6239__B1 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2137 _7002_/Q VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5125_ _4851_/Y _5294_/A _5064_/Y _4968_/X _5124_/X VGND VGND VPWR VPWR _5125_/Y
+ sky130_fd_sc_hd__a221oi_1
Xhold1403 _7287_/Q VGND VGND VPWR VPWR _5669_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2148 _4366_/X VGND VGND VPWR VPWR hold406/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4149__S _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2159 hold407/X VGND VGND VPWR VPWR _4505_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1414 _7258_/Q VGND VGND VPWR VPWR hold1414/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1425 hold15/X VGND VGND VPWR VPWR _4197_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1436 hold1436/A VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1447 _4085_/A2 VGND VGND VPWR VPWR _4179_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5056_ _5056_/A _5056_/B _5056_/C VGND VGND VPWR VPWR _5060_/C sky130_fd_sc_hd__nand3_1
Xhold1458 _5899_/X VGND VGND VPWR VPWR hold131/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1469 _7556_/Q VGND VGND VPWR VPWR hold186/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4007_ _4062_/A _4007_/B VGND VGND VPWR VPWR _4040_/D sky130_fd_sc_hd__nand2_4
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout457_A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7219__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6411__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout624_A _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5958_ _5958_/A0 _5985_/A1 _5964_/S VGND VGND VPWR VPWR _5958_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3776__A1 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4909_ _4909_/A _4924_/B _4909_/C _4909_/D VGND VGND VPWR VPWR _4915_/C sky130_fd_sc_hd__and4_2
XANTENNA__4973__B1 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5889_ _5889_/A0 _5979_/A0 hold91/X VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5708__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7628_ _7646_/CLK _7628_/D fanout751/X VGND VGND VPWR VPWR _7628_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3528__A1 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__B2 _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6190__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6112__B _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7559_ _7561_/CLK _7559_/D fanout738/X VGND VGND VPWR VPWR _7559_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input157_A wb_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3350 _7221_/Q VGND VGND VPWR VPWR _3573_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3361 _6892_/Q VGND VGND VPWR VPWR _4064_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3372 _6890_/Q VGND VGND VPWR VPWR _4123_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3700__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2660 hold729/X VGND VGND VPWR VPWR _4339_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2671 hold691/X VGND VGND VPWR VPWR _4375_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2682 _5819_/X VGND VGND VPWR VPWR hold924/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2693 _5801_/X VGND VGND VPWR VPWR hold896/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1970 _5691_/X VGND VGND VPWR VPWR hold279/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1981 _7539_/Q VGND VGND VPWR VPWR hold294/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input18_A mask_rev_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1992 _7100_/Q VGND VGND VPWR VPWR hold272/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3767__A1 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3767__B2 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6705__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6705__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3646__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6181__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4192__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _3782_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6469__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4758__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3662__A _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5141__B1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6641__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6930_ _7601_/CLK _6930_/D fanout688/X VGND VGND VPWR VPWR _6930_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6861_ _6861_/A _6873_/B VGND VGND VPWR VPWR _6861_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_6_csclk _7416_/CLK VGND VGND VPWR VPWR _7160_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4643__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2491_A _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5812_ _5866_/B _5956_/B _5956_/C VGND VGND VPWR VPWR _5820_/S sky130_fd_sc_hd__and3_4
X_6792_ _3570_/Y _6792_/A1 _6792_/S VGND VGND VPWR VPWR _7636_/D sky130_fd_sc_hd__mux2_1
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3758__A1 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5743_ _5743_/A0 _5968_/A1 _5748_/S VGND VGND VPWR VPWR _5743_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5674_ _5953_/A1 _5674_/A1 _5676_/S VGND VGND VPWR VPWR _5674_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3556__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7413_ _7478_/CLK _7413_/D fanout715/X VGND VGND VPWR VPWR _7413_/Q sky130_fd_sc_hd__dfrtp_4
X_4625_ _4910_/D _4856_/A _5399_/A VGND VGND VPWR VPWR _4625_/Y sky130_fd_sc_hd__nand3_4
XFILLER_135_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6172__A2 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7344_ _7539_/CLK _7344_/D fanout708/X VGND VGND VPWR VPWR _7344_/Q sky130_fd_sc_hd__dfstp_2
Xhold500 hold500/A VGND VGND VPWR VPWR _7576_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4556_ _5853_/A0 _4556_/A1 _4556_/S VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__mux2_1
Xhold522 _5823_/X VGND VGND VPWR VPWR _7424_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold533 hold533/A VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold544 hold544/A VGND VGND VPWR VPWR _7025_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3507_ _3507_/A hold38/X _4509_/C VGND VGND VPWR VPWR _3507_/X sky130_fd_sc_hd__and3_2
Xhold555 hold555/A VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7275_ _7314_/CLK _7275_/D fanout714/X VGND VGND VPWR VPWR _7275_/Q sky130_fd_sc_hd__dfrtp_1
X_4487_ _5645_/A0 _4487_/A1 _4490_/S VGND VGND VPWR VPWR _4487_/X sky130_fd_sc_hd__mux2_1
Xhold566 _4200_/X VGND VGND VPWR VPWR _6917_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold577 hold577/A VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold588 _5628_/X VGND VGND VPWR VPWR _7254_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6226_ _7300_/Q _6074_/X _6267_/B1 _7396_/Q _6225_/X VGND VGND VPWR VPWR _6226_/X
+ sky130_fd_sc_hd__a221o_1
Xhold599 hold599/A VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3438_ _7338_/Q VGND VGND VPWR VPWR _3438_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6475__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5683__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6152_/X _6157_/B _6157_/C VGND VGND VPWR VPWR _6157_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_131_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout574_A _5635_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1200 hold2905/X VGND VGND VPWR VPWR _5622_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1211 hold2881/X VGND VGND VPWR VPWR _7530_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 hold2872/X VGND VGND VPWR VPWR hold2873/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5108_ _5059_/A _5061_/B _5524_/A3 _5107_/X VGND VGND VPWR VPWR _5111_/B sky130_fd_sc_hd__a31o_1
XANTENNA__6227__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1233 hold2933/X VGND VGND VPWR VPWR _7562_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1244 hold2897/X VGND VGND VPWR VPWR hold2898/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6088_ _7495_/Q _6085_/X _6087_/X _7463_/Q _6083_/X VGND VGND VPWR VPWR _6102_/B
+ sky130_fd_sc_hd__a221o_1
Xhold1255 _4393_/S VGND VGND VPWR VPWR _4391_/S sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1266 hold2947/X VGND VGND VPWR VPWR _7013_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6632__B1 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1277 hold3041/X VGND VGND VPWR VPWR hold3042/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5039_ _5039_/A _5039_/B _5039_/C VGND VGND VPWR VPWR _5041_/A sky130_fd_sc_hd__nor3_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout741_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1288 _5597_/X VGND VGND VPWR VPWR _7229_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1299 hold3261/X VGND VGND VPWR VPWR hold3262/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1689_A _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6699__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6163__A2 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4578__A _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3482__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3237_A _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR _4089_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR _4093_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3180 _7192_/Q VGND VGND VPWR VPWR hold3180/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5901__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR _6809_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3191 _7162_/Q VGND VGND VPWR VPWR hold3191/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR _6814_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR input164/X sky130_fd_sc_hd__buf_6
XANTENNA__4857__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2490 hold713/X VGND VGND VPWR VPWR _5757_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5426__A1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_3_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6387__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3657__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6154__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4410_ _4442_/A0 _5976_/A0 _4422_/S VGND VGND VPWR VPWR _4410_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4165__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5390_ _5390_/A _5518_/C _5473_/C VGND VGND VPWR VPWR _5394_/A sky130_fd_sc_hd__and3_1
X_4341_ _5582_/A0 _4341_/A1 _4345_/S VGND VGND VPWR VPWR _4341_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7060_ _7191_/CLK _7060_/D fanout701/X VGND VGND VPWR VPWR _7060_/Q sky130_fd_sc_hd__dfrtp_2
X_4272_ _4272_/A0 _5876_/A1 _4276_/S VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6011_ _7585_/Q _7584_/Q _6932_/Q _6009_/B VGND VGND VPWR VPWR _6011_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5665__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5811__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2504_A _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3691__A3 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3979__A1 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6913_ _7264_/CLK _6913_/D fanout688/X VGND VGND VPWR VPWR _6913_/Q sky130_fd_sc_hd__dfstp_4
X_6844_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6844_/X sky130_fd_sc_hd__and2_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6775_ _6961_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6775_/X sky130_fd_sc_hd__o21a_1
X_3987_ _7287_/Q _5668_/A _3983_/X _3985_/X _3986_/X VGND VGND VPWR VPWR _3988_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5726_ _5726_/A0 _5726_/A1 _5730_/S VGND VGND VPWR VPWR _5726_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3600__B1 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5657_ _5954_/A1 _5657_/A1 _5657_/S VGND VGND VPWR VPWR _5657_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4156__A1 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4608_ _4879_/D _4747_/B _4887_/B _4945_/A VGND VGND VPWR VPWR _4608_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ _5588_/A0 _5732_/A1 _5589_/S VGND VGND VPWR VPWR _5588_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3903__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7327_ _7327_/CLK _7327_/D fanout703/X VGND VGND VPWR VPWR _7327_/Q sky130_fd_sc_hd__dfstp_2
X_4539_ _5612_/A _5596_/A _4539_/C _5619_/C VGND VGND VPWR VPWR _4544_/S sky130_fd_sc_hd__and4_4
Xhold341 _3466_/X VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3903__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold352 hold352/A VGND VGND VPWR VPWR _7304_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout691_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold363 hold363/A VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7258_ _7578_/CLK hold6/X fanout747/X VGND VGND VPWR VPWR _7258_/Q sky130_fd_sc_hd__dfrtp_4
Xhold396 hold396/A VGND VGND VPWR VPWR _7520_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6209_ _7459_/Q _6080_/X _6092_/X _7531_/Q _6208_/X VGND VGND VPWR VPWR _6209_/X
+ sky130_fd_sc_hd__a221o_1
X_7189_ _7268_/CLK _7189_/D _6869_/A VGND VGND VPWR VPWR _7189_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_58_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 hold3067/X VGND VGND VPWR VPWR hold3068/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1041 hold2830/X VGND VGND VPWR VPWR hold2831/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5408__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1052 _5615_/X VGND VGND VPWR VPWR _7244_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6605__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1063 hold1063/A VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
XTAP_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1074 hold3002/X VGND VGND VPWR VPWR hold1074/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 hold1085/A VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
XFILLER_85_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5022__A _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 hold3010/X VGND VGND VPWR VPWR hold1096/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1973_A _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input85_A spimemio_flash_io0_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6788__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6727__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4855__C1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4247__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7238_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3910_ _7496_/Q hold41/A _3651_/X _7047_/Q _3909_/X VGND VGND VPWR VPWR _3913_/C
+ sky130_fd_sc_hd__a221o_1
X_4890_ _5222_/B _5222_/C _5049_/C _4891_/D VGND VGND VPWR VPWR _5223_/D sky130_fd_sc_hd__nand4_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3841_ _7393_/Q _4473_/A _5785_/B _3665_/X _7124_/Q VGND VGND VPWR VPWR _3841_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4921__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2287_A _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5583__A0 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3772_ _7049_/Q _3651_/X _3767_/X _3769_/X _3771_/X VGND VGND VPWR VPWR _3772_/X
+ sky130_fd_sc_hd__a2111o_1
X_6560_ _7379_/Q _6408_/B _6555_/X _6557_/X _6559_/X VGND VGND VPWR VPWR _6570_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5511_ _4843_/A _4659_/Y _5081_/A _5541_/D _5247_/C VGND VGND VPWR VPWR _5512_/D
+ sky130_fd_sc_hd__o311a_1
X_6491_ _7464_/Q _6434_/X _6460_/X _7384_/Q _6490_/X VGND VGND VPWR VPWR _6494_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5806__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4138__A1 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5442_ _5059_/A _5203_/A _5342_/B _5205_/X VGND VGND VPWR VPWR _5442_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6678__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ _4744_/Y _5509_/A3 _4880_/Y _4846_/Y VGND VGND VPWR VPWR _5373_/X sky130_fd_sc_hd__a31o_1
XFILLER_160_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3897__B1 _3889_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7471_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5107__A _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4324_ hold198/X _4324_/A1 _4327_/S VGND VGND VPWR VPWR _4324_/X sky130_fd_sc_hd__mux2_1
X_7112_ _7186_/CLK _7112_/D fanout725/X VGND VGND VPWR VPWR _7112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7043_ _7201_/CLK _7043_/D _6839_/A VGND VGND VPWR VPWR _7043_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_86_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4255_ _4255_/A0 _5997_/A1 _4258_/S VGND VGND VPWR VPWR _4255_/X sky130_fd_sc_hd__mux2_1
X_4186_ _4186_/A0 _5914_/A1 _4190_/S VGND VGND VPWR VPWR _4186_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7575_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_3_1_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7416_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_103_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4681__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3821__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6827_ _7105_/Q _7105_/D VGND VGND VPWR VPWR _6827_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6366__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4377__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6758_ _7136_/Q _6409_/X _6753_/X _6757_/X _6430_/X VGND VGND VPWR VPWR _6758_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3719__A4 _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5709_ _5952_/A1 _5709_/A1 _5712_/S VGND VGND VPWR VPWR _5709_/X sky130_fd_sc_hd__mux2_1
X_6689_ _7198_/Q _6463_/A _6771_/A3 _6408_/D _7168_/Q VGND VGND VPWR VPWR _6689_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5877__A1 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6120__B _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold171 hold171/A VGND VGND VPWR VPWR _7293_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5629__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5058__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4856__A _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout651 _5404_/D VGND VGND VPWR VPWR _5203_/C sky130_fd_sc_hd__buf_8
Xfanout662 _5068_/B VGND VGND VPWR VPWR _5260_/C sky130_fd_sc_hd__buf_6
XFILLER_144_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout673 wire674/X VGND VGND VPWR VPWR _5134_/A sky130_fd_sc_hd__buf_6
Xfanout684 input99/X VGND VGND VPWR VPWR _4840_/D sky130_fd_sc_hd__buf_6
XANTENNA__4575__B _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout695 _6861_/A VGND VGND VPWR VPWR _6869_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_74_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold3102_A _7479_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6896__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4368__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output289_A _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5868__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3894__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3670__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4040_ _4040_/A _6900_/Q _6901_/Q _4040_/D VGND VGND VPWR VPWR _4042_/A sky130_fd_sc_hd__and4_1
XANTENNA__4485__B _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6045__A1 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6596__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5991_ _5991_/A0 _5991_/A1 _5991_/S VGND VGND VPWR VPWR _5991_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4942_ _4942_/A _5248_/B _4948_/C _4970_/C VGND VGND VPWR VPWR _4944_/B sky130_fd_sc_hd__nand4_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3803__B1 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7661_ _7661_/A VGND VGND VPWR VPWR _7661_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_177_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _4667_/A _4667_/B _4984_/B _4984_/A VGND VGND VPWR VPWR _4873_/X sky130_fd_sc_hd__o22a_4
XFILLER_178_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6612_ _7593_/Q _7581_/Q _6408_/C _6611_/X VGND VGND VPWR VPWR _6612_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4359__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3824_ _7252_/Q _5659_/B _5623_/B _3663_/X _7164_/Q VGND VGND VPWR VPWR _3824_/X
+ sky130_fd_sc_hd__a32o_1
X_7592_ _7610_/CLK _7592_/D fanout693/X VGND VGND VPWR VPWR _7592_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6543_ _7314_/Q _6419_/D _6454_/X _7490_/Q _6542_/X VGND VGND VPWR VPWR _6544_/D
+ sky130_fd_sc_hd__a221o_1
X_3755_ _4168_/D _3552_/X _3652_/X _7150_/Q VGND VGND VPWR VPWR _3755_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold2836_A _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3582__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3686_ _7233_/Q _3617_/X _3681_/X _3683_/X _3685_/X VGND VGND VPWR VPWR _3686_/X
+ sky130_fd_sc_hd__a2111o_4
X_6474_ _7593_/Q _7576_/Q _6408_/C _6058_/X _7528_/Q VGND VGND VPWR VPWR _6474_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3564__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput210 _3438_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
X_5425_ _4888_/C _4997_/B _5199_/C _4758_/X VGND VGND VPWR VPWR _5425_/X sky130_fd_sc_hd__a31o_2
Xoutput221 _7659_/X VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
XANTENNA__6520__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 _7669_/X VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput243 _4152_/X VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__4531__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput254 _4132_/Y VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
X_5356_ _5089_/D _4939_/C _4877_/A VGND VGND VPWR VPWR _5450_/B sky130_fd_sc_hd__o21ai_1
Xoutput265 _7222_/Q VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
Xoutput276 _7235_/Q VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 _6921_/Q VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XANTENNA__3885__A3 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4307_ _4307_/A0 _5625_/A1 _4308_/S VGND VGND VPWR VPWR _4307_/X sky130_fd_sc_hd__mux2_1
Xoutput298 _7247_/Q VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
X_5287_ _5061_/B _5453_/C _4845_/X VGND VGND VPWR VPWR _5294_/B sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout487_A _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5087__A2 _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4238_ _5653_/A1 _5995_/A1 _4248_/S VGND VGND VPWR VPWR _4238_/X sky130_fd_sc_hd__mux2_1
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7026_ _7035_/CLK _7026_/D fanout723/X VGND VGND VPWR VPWR _7026_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_68_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4169_ _4429_/B _4169_/A2 _4168_/Y _4169_/B2 VGND VGND VPWR VPWR _4169_/X sky130_fd_sc_hd__a22o_2
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6587__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5795__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5938__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire348 _3642_/Y VGND VGND VPWR VPWR _3643_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6511__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4522__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3876__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input48_A mgmt_gpio_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3490__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6275__A1 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__B2 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout481 _6404_/Y VGND VGND VPWR VPWR _6561_/A2 sky130_fd_sc_hd__buf_6
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3628__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5483__C1 _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout492 _6056_/X VGND VGND VPWR VPWR _6447_/C sky130_fd_sc_hd__buf_8
XFILLER_120_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4598__A_N _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6290__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6578__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7074__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3649__B _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5250__A2 _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3800__A3 _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3540_ _7438_/Q _3525_/X _3528_/X _3534_/X _3539_/X VGND VGND VPWR VPWR _3568_/A
+ sky130_fd_sc_hd__a2111o_1
Xmax_cap604 _3856_/A VGND VGND VPWR VPWR _3923_/S sky130_fd_sc_hd__clkbuf_4
Xhold907 hold907/A VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold918 hold918/A VGND VGND VPWR VPWR _7027_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold929 hold929/A VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3471_ hold75/X hold38/X VGND VGND VPWR VPWR hold76/A sky130_fd_sc_hd__and2_1
XANTENNA__6502__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap659 _4765_/B VGND VGND VPWR VPWR _4717_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_182_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5210_ _4601_/Y _4716_/Y _4726_/Y _4906_/B VGND VGND VPWR VPWR _5210_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5710__A0 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4513__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6190_ _7282_/Q _6036_/Y _6178_/X _6189_/X _6623_/B1 VGND VGND VPWR VPWR _6190_/X
+ sky130_fd_sc_hd__o221a_1
Xhold3009 _6994_/Q VGND VGND VPWR VPWR _4312_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_170_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5141_ _4706_/Y _4741_/Y _4759_/Y _4761_/Y _5139_/X VGND VGND VPWR VPWR _5143_/B
+ sky130_fd_sc_hd__o221a_1
Xhold2308 _5608_/X VGND VGND VPWR VPWR hold594/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2319 hold747/X VGND VGND VPWR VPWR _5909_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1607 hold129/X VGND VGND VPWR VPWR _7238_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5072_ _5399_/B _5072_/B _5115_/C _5072_/D VGND VGND VPWR VPWR _5072_/Y sky130_fd_sc_hd__nand4_4
Xhold1618 _7293_/Q VGND VGND VPWR VPWR hold170/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1629 _3448_/X VGND VGND VPWR VPWR _3449_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ _4023_/A1 _4007_/B _4022_/X VGND VGND VPWR VPWR _4023_/X sky130_fd_sc_hd__a21o_1
XFILLER_84_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5777__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5974_ _5974_/A _5992_/D VGND VGND VPWR VPWR _5982_/S sky130_fd_sc_hd__nand2_8
XANTENNA__3788__C1 _3787_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4925_ _4925_/A _5444_/C _4925_/C VGND VGND VPWR VPWR _4927_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6650__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7644_ _7646_/CLK _7644_/D fanout753/X VGND VGND VPWR VPWR _7644_/Q sky130_fd_sc_hd__dfrtp_1
X_4856_ _4856_/A _4888_/B _5058_/D VGND VGND VPWR VPWR _4856_/Y sky130_fd_sc_hd__nor3b_2
X_3807_ _6990_/Q _3562_/C _5623_/B _3531_/X _7337_/Q VGND VGND VPWR VPWR _3807_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7575_ _7575_/CLK _7575_/D fanout734/X VGND VGND VPWR VPWR _7575_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6741__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4787_ _4836_/C _4797_/B VGND VGND VPWR VPWR _4787_/Y sky130_fd_sc_hd__nand2_1
X_6526_ _7562_/Q _6419_/C _6466_/X _7506_/Q _6525_/X VGND VGND VPWR VPWR _6526_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4752__B2 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3738_ _7261_/Q _3738_/B _4265_/B VGND VGND VPWR VPWR _3738_/X sky130_fd_sc_hd__and3_1
XFILLER_174_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6457_ _6466_/B _6466_/C _6466_/D _6466_/A VGND VGND VPWR VPWR _6457_/X sky130_fd_sc_hd__and4b_4
XFILLER_173_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3669_ _4515_/B _4509_/C _4352_/A VGND VGND VPWR VPWR _3669_/X sky130_fd_sc_hd__and3_4
X_5408_ _5113_/A _5404_/D _5410_/A VGND VGND VPWR VPWR _5408_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6388_ _7060_/Q _6110_/A _6388_/A3 _6082_/X _7010_/Q VGND VGND VPWR VPWR _6388_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5339_ _5339_/A _5339_/B _5339_/C _5339_/D VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__nand4_2
Xhold2820 _4305_/X VGND VGND VPWR VPWR hold884/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2831 hold2831/A VGND VGND VPWR VPWR _4224_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2842 _6947_/Q VGND VGND VPWR VPWR hold2842/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2853 _6913_/Q VGND VGND VPWR VPWR hold2853/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2864 hold2864/A VGND VGND VPWR VPWR _5606_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2875 hold2875/A VGND VGND VPWR VPWR _5888_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5014__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7009_ _7191_/CLK _7009_/D fanout700/X VGND VGND VPWR VPWR _7009_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2886 _7660_/A VGND VGND VPWR VPWR hold2886/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2897 _7003_/Q VGND VGND VPWR VPWR hold2897/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4853__B _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5030__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4572__C _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input102_A wb_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4440__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5965__A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6193__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6732__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3546__A2 hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5904__S hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5299__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4747__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3651__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5471__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5759__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6036__A _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _5113_/A _5089_/B _5089_/C VGND VGND VPWR VPWR _4803_/A sky130_fd_sc_hd__and3_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A2 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_29_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5690_ _5951_/A1 hold365/X _5694_/S VGND VGND VPWR VPWR _5690_/X sky130_fd_sc_hd__mux2_1
X_4641_ _4641_/A _4641_/B _4730_/C _4768_/B VGND VGND VPWR VPWR _5158_/B sky130_fd_sc_hd__nor4_4
XFILLER_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6723__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5931__A0 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7360_ _7360_/CLK _7360_/D fanout706/X VGND VGND VPWR VPWR _7360_/Q sky130_fd_sc_hd__dfstp_4
X_4572_ _5058_/D _4888_/B _4888_/C VGND VGND VPWR VPWR _4668_/C sky130_fd_sc_hd__and3_4
XFILLER_116_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold704 hold704/A VGND VGND VPWR VPWR _6878_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6311_ _7113_/Q _6317_/C _6074_/X _6968_/Q _6310_/X VGND VGND VPWR VPWR _6311_/X
+ sky130_fd_sc_hd__a221o_1
Xhold715 hold715/A VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3523_ _7374_/Q _5758_/A _3519_/X _7550_/Q _3522_/X VGND VGND VPWR VPWR _3524_/D
+ sky130_fd_sc_hd__a221o_1
Xmax_cap423 _4850_/B VGND VGND VPWR VPWR _5166_/A2 sky130_fd_sc_hd__clkbuf_2
Xhold726 _5844_/X VGND VGND VPWR VPWR _7443_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7291_ _7329_/CLK hold3/X fanout704/X VGND VGND VPWR VPWR _7291_/Q sky130_fd_sc_hd__dfrtp_4
Xhold737 hold737/A VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5814__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold748 hold748/A VGND VGND VPWR VPWR _7501_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap467 _4884_/B VGND VGND VPWR VPWR _4954_/C sky130_fd_sc_hd__buf_4
X_6242_ _7389_/Q _6274_/A3 _6267_/B1 _7397_/Q _6241_/X VGND VGND VPWR VPWR _6242_/X
+ sky130_fd_sc_hd__a221o_1
X_3454_ _4181_/S hold45/X _3453_/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__o21ba_1
Xhold759 hold759/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6173_ _7410_/Q _6144_/C _6089_/C _6144_/B VGND VGND VPWR VPWR _6173_/X sky130_fd_sc_hd__o211a_1
Xhold2105 hold530/X VGND VGND VPWR VPWR _6934_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2116 hold322/X VGND VGND VPWR VPWR _4541_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5115__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2127 _4232_/X VGND VGND VPWR VPWR hold478/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2138 hold399/X VGND VGND VPWR VPWR _4324_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5124_ _5122_/Y _5123_/X _5580_/A2 VGND VGND VPWR VPWR _5124_/X sky130_fd_sc_hd__a21o_1
Xhold1404 hold2958/X VGND VGND VPWR VPWR hold2959/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2149 _7398_/Q VGND VGND VPWR VPWR hold2149/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1415 hold1415/A VGND VGND VPWR VPWR _5635_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1426 _4197_/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1437 _6888_/Q VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5055_ _5295_/A _5113_/A _5055_/C _5295_/D VGND VGND VPWR VPWR _5056_/C sky130_fd_sc_hd__nand4_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1448 _4179_/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1459 hold131/X VGND VGND VPWR VPWR _7492_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4006_ _4006_/A _4006_/B VGND VGND VPWR VPWR _6908_/D sky130_fd_sc_hd__nor2_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4670__B1 _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6411__A1 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5214__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5957_ _5957_/A0 _5993_/A1 _5964_/S VGND VGND VPWR VPWR _5957_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5785__A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__A2 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__A1 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4908_ wire649/X _4877_/A _4907_/X _4906_/Y VGND VGND VPWR VPWR _4913_/A sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout617_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5888_ _5888_/A0 _5978_/A0 hold91/X VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7627_ _7627_/CLK _7627_/D fanout691/X VGND VGND VPWR VPWR _7627_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6175__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4839_ _5011_/B _4839_/B VGND VGND VPWR VPWR _5496_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6714__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__A2 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7558_ _7576_/CLK _7558_/D fanout718/X VGND VGND VPWR VPWR _7558_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_181_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6509_ _7313_/Q _6419_/D _6424_/X _7569_/Q _6508_/X VGND VGND VPWR VPWR _6509_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7489_ _7489_/CLK _7489_/D fanout719/X VGND VGND VPWR VPWR _7489_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5724__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6478__A1 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4489__A0 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3340 _7075_/Q VGND VGND VPWR VPWR _4120_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3351 _6903_/Q VGND VGND VPWR VPWR _4036_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3362 _4064_/X VGND VGND VPWR VPWR _6892_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3373 _6901_/Q VGND VGND VPWR VPWR _4041_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3700__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__buf_6
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__buf_4
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__buf_4
Xhold2650 hold825/X VGND VGND VPWR VPWR _4513_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2661 _4339_/X VGND VGND VPWR VPWR hold730/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_152_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2672 _4375_/X VGND VGND VPWR VPWR hold692/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2683 _7136_/Q VGND VGND VPWR VPWR hold669/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__clkbuf_2
Xhold2694 _7475_/Q VGND VGND VPWR VPWR hold811/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1960 hold146/X VGND VGND VPWR VPWR _5703_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1971 _7148_/Q VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1982 hold294/X VGND VGND VPWR VPWR _5952_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1993 hold272/X VGND VGND VPWR VPWR _4448_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4661__B1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4075__S _4075_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5695__A _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3767__A2 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3927__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6166__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3646__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 _3800_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6469__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4758__B _5012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3662__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4924__D _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6860_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6860_/X sky130_fd_sc_hd__and2_1
X_5811_ _5811_/A0 _5955_/A1 _5811_/S VGND VGND VPWR VPWR _5811_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6791_ _3607_/Y _6791_/A1 _6792_/S VGND VGND VPWR VPWR _7635_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5809__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3758__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5742_ _5742_/A0 _5976_/A0 _5748_/S VGND VGND VPWR VPWR _5742_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4955__B2 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4940__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5673_ _5673_/A0 _7291_/Q _5676_/S VGND VGND VPWR VPWR _5673_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5904__A0 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7412_ _7421_/CLK _7412_/D fanout715/X VGND VGND VPWR VPWR _7412_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3556__C _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4624_ _4910_/D _4856_/A _5399_/A VGND VGND VPWR VPWR _4997_/A sky130_fd_sc_hd__and3_4
X_7343_ _7360_/CLK _7343_/D fanout703/X VGND VGND VPWR VPWR _7343_/Q sky130_fd_sc_hd__dfstp_2
Xhold501 hold501/A VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4555_ _4555_/A0 _4555_/A1 _4556_/S VGND VGND VPWR VPWR _4555_/X sky130_fd_sc_hd__mux2_1
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold523 hold523/A VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold534 hold534/A VGND VGND VPWR VPWR _7077_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3506_ _5740_/A _5938_/A _4509_/C VGND VGND VPWR VPWR _3506_/X sky130_fd_sc_hd__and3_4
Xhold545 hold545/A VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7274_ _7306_/CLK _7274_/D _4079_/A VGND VGND VPWR VPWR _7274_/Q sky130_fd_sc_hd__dfrtp_1
Xhold556 _4264_/X VGND VGND VPWR VPWR _6961_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4486_ _5732_/A1 _4486_/A1 _4490_/S VGND VGND VPWR VPWR _4486_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4668__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold567 hold567/A VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold578 _4208_/X VGND VGND VPWR VPWR _6923_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5132__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold589 hold589/A VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6225_ _7292_/Q _6112_/B _6136_/C _6276_/A3 _7364_/Q VGND VGND VPWR VPWR _6225_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3437_ _7346_/Q VGND VGND VPWR VPWR _3437_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _7369_/Q _6111_/X _6121_/X _7305_/Q _6155_/X VGND VGND VPWR VPWR _6157_/C
+ sky130_fd_sc_hd__a221oi_1
XFILLER_106_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 hold2906/X VGND VGND VPWR VPWR _7249_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1212 hold2926/X VGND VGND VPWR VPWR hold2927/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1223 _4435_/X VGND VGND VPWR VPWR _7088_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5134_/A _5118_/A _5107_/C VGND VGND VPWR VPWR _5107_/X sky130_fd_sc_hd__and3_1
Xhold1234 hold2919/X VGND VGND VPWR VPWR hold2920/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6087_ _6317_/B _6121_/A _6097_/C VGND VGND VPWR VPWR _6087_/X sky130_fd_sc_hd__and3_4
XFILLER_181_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout567_A _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1245 hold2899/X VGND VGND VPWR VPWR _7003_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1256 hold2960/X VGND VGND VPWR VPWR _7058_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1267 hold2948/X VGND VGND VPWR VPWR hold2949/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1278 hold3043/X VGND VGND VPWR VPWR _7450_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5038_ _5038_/A _5038_/B _5038_/C VGND VGND VPWR VPWR _5039_/B sky130_fd_sc_hd__and3_1
Xhold1289 hold3224/X VGND VGND VPWR VPWR hold3225/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5011__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6989_ _6991_/CLK _6989_/D fanout693/X VGND VGND VPWR VPWR _6989_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4850__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5371__A1 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4859__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3482__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6320__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3132_A _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR _4887_/D sky130_fd_sc_hd__buf_4
XFILLER_49_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR input121/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3170 _4468_/X VGND VGND VPWR VPWR hold3170/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR _6800_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input30_A mask_rev_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3181 hold3181/A VGND VGND VPWR VPWR _4546_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR _6803_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3192 hold3192/A VGND VGND VPWR VPWR _4510_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR _6806_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR _6793_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2480 _4405_/X VGND VGND VPWR VPWR hold750/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5426__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2491 _7515_/Q VGND VGND VPWR VPWR hold639/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4634__B1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1790 _7203_/Q VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6387__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_7_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3673__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4340_ _4340_/A _5619_/C VGND VGND VPWR VPWR _4345_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3912__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4271_ _4551_/C _4509_/C _4352_/A _4533_/B VGND VGND VPWR VPWR _4276_/S sky130_fd_sc_hd__and4_2
XANTENNA__6311__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6010_ _7585_/Q _7584_/Q VGND VGND VPWR VPWR _6010_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ _7264_/CLK _6912_/D fanout688/X VGND VGND VPWR VPWR _6912_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_63_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6843_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6843_/X sky130_fd_sc_hd__and2_1
XFILLER_62_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7188__RESET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4443__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2866_A _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6774_ _6758_/X _6774_/B _6774_/C VGND VGND VPWR VPWR _6774_/Y sky130_fd_sc_hd__nand3b_4
X_3986_ _7415_/Q _3544_/X _3565_/X _7463_/Q _3925_/X VGND VGND VPWR VPWR _3986_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6393__A3 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5725_ _5725_/A0 _5995_/A1 _5730_/S VGND VGND VPWR VPWR _5725_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5656_ _5881_/A1 _5656_/A1 _5657_/S VGND VGND VPWR VPWR _5656_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4607_ _4879_/D _4747_/B _4887_/B _4945_/A VGND VGND VPWR VPWR _4645_/D sky130_fd_sc_hd__o211a_4
XANTENNA__6550__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5587_ _5612_/A _5640_/A _5619_/A _5640_/D VGND VGND VPWR VPWR _5589_/S sky130_fd_sc_hd__and4_1
Xhold320 hold320/A VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7326_ _7582_/CLK _7326_/D fanout717/X VGND VGND VPWR VPWR _7326_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 _5826_/X VGND VGND VPWR VPWR _7427_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3903__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4538_ _5826_/A1 _4538_/A1 _4538_/S VGND VGND VPWR VPWR _4538_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold342 _3505_/A VGND VGND VPWR VPWR _3576_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold353 hold353/A VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold364 hold364/A VGND VGND VPWR VPWR _7134_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold375 _7296_/Q VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6302__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7257_ _7580_/CLK _7257_/D fanout735/X VGND VGND VPWR VPWR _7257_/Q sky130_fd_sc_hd__dfrtp_4
Xhold386 hold386/A VGND VGND VPWR VPWR _7536_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4469_ _4553_/A0 _4469_/A1 _4472_/S VGND VGND VPWR VPWR _4469_/X sky130_fd_sc_hd__mux2_1
Xhold397 hold397/A VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6208_ _7427_/Q _6110_/A _6074_/X _6100_/X _7475_/Q VGND VGND VPWR VPWR _6208_/X
+ sky130_fd_sc_hd__a32o_1
X_7188_ _7191_/CLK _7188_/D fanout728/X VGND VGND VPWR VPWR _7188_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _7400_/Q _6091_/X _6119_/D _7312_/Q _6116_/X VGND VGND VPWR VPWR _6139_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 hold3032/X VGND VGND VPWR VPWR hold3033/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1031 _5678_/X VGND VGND VPWR VPWR _7295_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 hold2832/X VGND VGND VPWR VPWR _6936_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5408__A2 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1053 hold2847/X VGND VGND VPWR VPWR hold2848/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1064 hold3092/X VGND VGND VPWR VPWR hold3093/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1075 hold1075/A VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 hold2979/X VGND VGND VPWR VPWR hold1086/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 hold1097/A VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
XANTENNA__5022__B _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6384__A3 _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5592__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3082_A _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input78_A spi_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6541__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_csclk _7416_/CLK VGND VGND VPWR VPWR _7268_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output234_A _4146_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4755__C _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4607__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3668__A _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3840_ _7184_/Q _4533_/A _4497_/A _7154_/Q _3839_/X VGND VGND VPWR VPWR _3840_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_189_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3771_ _7498_/Q hold41/A _5581_/A _7212_/Q _3770_/X VGND VGND VPWR VPWR _3771_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5510_ _5510_/A _5510_/B _5510_/C VGND VGND VPWR VPWR _5548_/A sky130_fd_sc_hd__and3_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6490_ _7496_/Q _6600_/B _6651_/C _6419_/C _7560_/Q VGND VGND VPWR VPWR _6490_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6127__A3 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5441_ _5343_/B _5343_/A _5441_/C _5506_/D VGND VGND VPWR VPWR _5441_/X sky130_fd_sc_hd__and4bb_1
XFILLER_172_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6532__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5372_ _5252_/A _5370_/Y _5371_/X _4854_/X VGND VGND VPWR VPWR _5372_/X sky130_fd_sc_hd__o31a_1
XFILLER_160_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7111_ _7111_/CLK _7111_/D _6780_/B VGND VGND VPWR VPWR _7111_/Q sky130_fd_sc_hd__dfrtp_4
X_4323_ _5732_/A1 _4323_/A1 _4327_/S VGND VGND VPWR VPWR _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5822__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ _7201_/CLK _7042_/D fanout726/X VGND VGND VPWR VPWR _7042_/Q sky130_fd_sc_hd__dfrtp_4
X_4254_ _4254_/A0 _5969_/A1 _4258_/S VGND VGND VPWR VPWR _4254_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4946__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4185_ _4185_/A0 _4185_/A1 _4429_/B VGND VGND VPWR VPWR _4185_/X sky130_fd_sc_hd__mux2_4
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7369__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3821__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3821__B2 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6826_ _7109_/Q _6824_/C _6795_/B _6825_/X VGND VGND VPWR VPWR _6826_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6366__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6757_ _7181_/Q _6058_/X _6755_/X _6756_/X VGND VGND VPWR VPWR _6757_/X sky130_fd_sc_hd__a211o_1
X_3969_ _7026_/Q _4352_/A _4352_/B _3659_/X _7006_/Q VGND VGND VPWR VPWR _3969_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6771__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3585__B1 _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5708_ _5951_/A1 _5708_/A1 _5712_/S VGND VGND VPWR VPWR _5708_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6688_ _7153_/Q _6467_/X _6683_/X _6685_/X _6687_/X VGND VGND VPWR VPWR _6698_/B
+ sky130_fd_sc_hd__a2111oi_4
XFILLER_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5639_ _5975_/A0 _5639_/A1 _5639_/S VGND VGND VPWR VPWR _5639_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3888__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold150 hold150/A VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7309_ _7309_/CLK _7309_/D fanout710/X VGND VGND VPWR VPWR _7309_/Q sky130_fd_sc_hd__dfrtp_4
Xhold161 hold161/A VGND VGND VPWR VPWR _7558_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold172 hold172/A VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold183 hold183/A VGND VGND VPWR VPWR _7301_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold194 hold194/A VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout630 _7084_/Q VGND VGND VPWR VPWR _4429_/B sky130_fd_sc_hd__buf_8
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout652 _4840_/X VGND VGND VPWR VPWR _5404_/D sky130_fd_sc_hd__clkbuf_16
Xfanout663 _5068_/B VGND VGND VPWR VPWR _5387_/C sky130_fd_sc_hd__buf_4
Xfanout685 _6864_/A VGND VGND VPWR VPWR _6873_/A sky130_fd_sc_hd__clkbuf_8
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout696 _6872_/A VGND VGND VPWR VPWR _6861_/A sky130_fd_sc_hd__buf_4
XANTENNA_input132_A wb_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6054__A2 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__A _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3812__B2 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4083__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6762__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5907__S hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3591__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3654__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6817__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6817__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3670__B _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6293__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6045__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5990_ _5990_/A0 _5990_/A1 _5991_/S VGND VGND VPWR VPWR _5990_/X sky130_fd_sc_hd__mux2_1
X_4941_ _4941_/A _4941_/B _4941_/C VGND VGND VPWR VPWR _4944_/A sky130_fd_sc_hd__nor3_1
XANTENNA__4932__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7660_ _7660_/A VGND VGND VPWR VPWR _7660_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4872_ _4840_/D _5399_/A _4910_/D VGND VGND VPWR VPWR _4956_/B sky130_fd_sc_hd__nand3b_4
XFILLER_60_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6348__A3 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6611_ _7437_/Q _6747_/B _6468_/C _6408_/A _7557_/Q VGND VGND VPWR VPWR _6611_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_178_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3823_ _7465_/Q _3565_/X _3651_/X _7048_/Q _3822_/X VGND VGND VPWR VPWR _3828_/C
+ sky130_fd_sc_hd__a221o_1
X_7591_ _7594_/CLK _7591_/D fanout694/X VGND VGND VPWR VPWR _7591_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6753__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5817__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6542_ _7474_/Q _6574_/B _6441_/X _6452_/X _7346_/Q VGND VGND VPWR VPWR _6542_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3754_ _7514_/Q _5920_/A _3673_/X _7200_/Q _3753_/X VGND VGND VPWR VPWR _3759_/B
+ sky130_fd_sc_hd__a221o_1
X_6473_ _6472_/X _6623_/B1 _6067_/B _6573_/S _6473_/B2 VGND VGND VPWR VPWR _6473_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6505__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3685_ _7161_/Q _4539_/C _5632_/B _3684_/X VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__a31o_1
XFILLER_145_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3564__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5424_ _4956_/A _4687_/Y _4726_/Y _4880_/Y VGND VGND VPWR VPWR _5424_/X sky130_fd_sc_hd__o22a_1
Xoutput200 _3413_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 _3437_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 _4155_/X VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput233 _7649_/X VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
XFILLER_160_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput244 _7653_/X VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
XFILLER_114_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5355_ _5355_/A _5355_/B _5355_/C _5355_/D VGND VGND VPWR VPWR _5361_/A sky130_fd_sc_hd__and4_1
Xoutput255 _7232_/Q VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
Xoutput266 _7229_/Q VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_102_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6808__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput277 _7236_/Q VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6808__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4306_ _4306_/A0 _5815_/A1 _4308_/S VGND VGND VPWR VPWR _4306_/X sky130_fd_sc_hd__mux2_1
Xoutput288 _6922_/Q VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput299 _3929_/Y VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
X_5286_ _5222_/A _5059_/A _5203_/A _5285_/X VGND VGND VPWR VPWR _5286_/X sky130_fd_sc_hd__a31o_1
XFILLER_141_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7025_ _7497_/CLK _7025_/D fanout693/X VGND VGND VPWR VPWR _7025_/Q sky130_fd_sc_hd__dfrtp_4
X_4237_ _4237_/A0 _4236_/X _4249_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4295__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6823__A4 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4168_ _4429_/B _7257_/Q _7306_/Q _4168_/D VGND VGND VPWR VPWR _4168_/Y sky130_fd_sc_hd__nor4_2
XFILLER_83_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4692__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4099_ _7584_/Q _7586_/Q _7587_/Q _4099_/D VGND VGND VPWR VPWR _4099_/Y sky130_fd_sc_hd__nor4_1
XFILLER_83_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout647_A _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6809_ _4427_/B _6809_/A2 _6809_/B1 _4426_/Y _6808_/X VGND VGND VPWR VPWR _6809_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6744__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5727__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6412__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire349 _6749_/Y VGND VGND VPWR VPWR wire349/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_70_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3730__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3490__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6275__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 _6106_/X VGND VGND VPWR VPWR _6379_/B1 sky130_fd_sc_hd__buf_8
XANTENNA__4286__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout482 _6402_/Y VGND VGND VPWR VPWR _6468_/C sky130_fd_sc_hd__buf_6
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout493 _6443_/B VGND VGND VPWR VPWR _6467_/A sky130_fd_sc_hd__buf_8
XFILLER_47_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5786__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3649__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7184_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6735__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4210__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3665__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_38_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7580_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold908 hold908/A VGND VGND VPWR VPWR _7193_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold919 hold919/A VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3470_ _3469_/X _3470_/A1 _4181_/S VGND VGND VPWR VPWR _3470_/X sky130_fd_sc_hd__mux2_2
XFILLER_50_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5140_ _4625_/Y _4687_/Y _4761_/Y _4741_/Y _4706_/Y VGND VGND VPWR VPWR _5140_/X
+ sky130_fd_sc_hd__o32a_1
Xhold2309 _7651_/A VGND VGND VPWR VPWR hold573/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_25_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6266__A2 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5071_ _5071_/A _5071_/B _5071_/C _5004_/A1 VGND VGND VPWR VPWR _5071_/Y sky130_fd_sc_hd__nor4b_2
Xhold1608 _7253_/Q VGND VGND VPWR VPWR hold166/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1619 hold170/X VGND VGND VPWR VPWR _5675_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4022_ _4014_/B _4017_/Y _4021_/X _4040_/D VGND VGND VPWR VPWR _4022_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6671__C1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5973_ _5973_/A0 _6000_/A1 _5973_/S VGND VGND VPWR VPWR _5973_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _4997_/B _4924_/B _5053_/C _5342_/B VGND VGND VPWR VPWR _4925_/C sky130_fd_sc_hd__nand4_2
X_7643_ _7646_/CLK _7643_/D fanout753/X VGND VGND VPWR VPWR _7643_/Q sky130_fd_sc_hd__dfrtp_1
X_4855_ _4644_/Y _4646_/Y _5222_/C _5404_/D _4966_/A VGND VGND VPWR VPWR _4855_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_193_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3806_ _7529_/Q _3529_/X _3670_/X _7134_/Q _3805_/X VGND VGND VPWR VPWR _3806_/X
+ sky130_fd_sc_hd__a221o_4
X_7574_ _7574_/CLK _7574_/D fanout745/X VGND VGND VPWR VPWR _7574_/Q sky130_fd_sc_hd__dfrtp_4
X_4786_ _4767_/A _4909_/D _4805_/B _4786_/D VGND VGND VPWR VPWR _4790_/C sky130_fd_sc_hd__and4bb_4
XFILLER_165_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6525_ _7498_/Q _6447_/C _6769_/A3 _6467_/X _7418_/Q VGND VGND VPWR VPWR _6525_/X
+ sky130_fd_sc_hd__a32o_1
X_3737_ _7522_/Q _4431_/A _5938_/C VGND VGND VPWR VPWR _3737_/X sky130_fd_sc_hd__and3_1
XFILLER_109_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6456_ _7487_/Q _6454_/X _6455_/X _7455_/Q _6453_/X VGND VGND VPWR VPWR _6456_/X
+ sky130_fd_sc_hd__a221o_1
X_3668_ _3931_/B _4328_/A _4388_/B VGND VGND VPWR VPWR _4545_/A sky130_fd_sc_hd__and3_4
X_5407_ _5407_/A1 _4844_/B _5399_/B _5404_/D VGND VGND VPWR VPWR _5410_/C sky130_fd_sc_hd__a31o_1
XFILLER_161_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5701__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5162__C1 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6387_ _7146_/Q _6082_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6387_/X sky130_fd_sc_hd__o211a_1
X_3599_ _7317_/Q _5695_/A _5731_/B _3503_/X input32/X VGND VGND VPWR VPWR _3599_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout597_A hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5338_ _5183_/B _5329_/X _5337_/X VGND VGND VPWR VPWR _5340_/B sky130_fd_sc_hd__a21oi_1
Xhold2810 _7140_/Q VGND VGND VPWR VPWR hold995/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2821 _7416_/Q VGND VGND VPWR VPWR hold871/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2832 _4224_/X VGND VGND VPWR VPWR hold2832/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2843 hold2843/A VGND VGND VPWR VPWR _4247_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout764_A _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5269_ _4698_/Y _5255_/X _5561_/A1 _5254_/X _5268_/X VGND VGND VPWR VPWR _5269_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_87_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2854 hold2854/A VGND VGND VPWR VPWR _4194_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2865 _5606_/X VGND VGND VPWR VPWR hold2865/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7008_ _7268_/CLK _7008_/D fanout698/X VGND VGND VPWR VPWR _7008_/Q sky130_fd_sc_hd__dfstp_2
Xhold2876 _5888_/X VGND VGND VPWR VPWR hold2876/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2887 hold2887/A VGND VGND VPWR VPWR _4417_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2898 hold2898/A VGND VGND VPWR VPWR _4325_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6407__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3491__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5768__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3779__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4440__A1 _5650_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5965__B _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6717__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3546__A3 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5940__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input60_A mgmt_gpio_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6496__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6036__B _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5875__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A3 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _4733_/A _4733_/B _4641_/B VGND VGND VPWR VPWR _4778_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__6184__A1 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6184__B2 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4571_ _4887_/B _4945_/A VGND VGND VPWR VPWR _4571_/Y sky130_fd_sc_hd__nand2_8
XFILLER_162_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2262_A _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6310_ _6963_/Q _6144_/A _6144_/B _6379_/B1 _7123_/Q VGND VGND VPWR VPWR _6310_/X
+ sky130_fd_sc_hd__a32o_1
X_3522_ _7446_/Q hold31/A _3872_/A2 _3521_/X _7318_/Q VGND VGND VPWR VPWR _3522_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold705 hold705/A VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7290_ _7334_/CLK _7290_/D fanout710/X VGND VGND VPWR VPWR _7290_/Q sky130_fd_sc_hd__dfrtp_4
Xhold716 hold716/A VGND VGND VPWR VPWR _7414_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold727 hold727/A VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold738 hold738/A VGND VGND VPWR VPWR _7141_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6241_ _7293_/Q _6112_/B _6121_/B _6074_/X _7301_/Q VGND VGND VPWR VPWR _6241_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6487__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3453_ _3452_/X _3453_/A1 _4181_/S VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__mux2_1
Xmax_cap468 _4753_/C VGND VGND VPWR VPWR _4641_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_171_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6172_ _7362_/Q _6276_/A3 _6267_/B1 _7394_/Q _6171_/X VGND VGND VPWR VPWR _6172_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2106 _6935_/Q VGND VGND VPWR VPWR hold507/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2117 _4541_/X VGND VGND VPWR VPWR hold323/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6239__A2 _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5123_ _5495_/C1 _5480_/A1 _4826_/Y _4428_/B VGND VGND VPWR VPWR _5123_/X sky130_fd_sc_hd__o31a_1
Xhold2128 _7502_/Q VGND VGND VPWR VPWR hold2128/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2139 _4324_/X VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1405 _7644_/Q VGND VGND VPWR VPWR _4201_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1416 _5635_/X VGND VGND VPWR VPWR hold1416/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1427 hold16/X VGND VGND VPWR VPWR _4446_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1438 hold9/X VGND VGND VPWR VPWR _4199_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5054_ _5342_/A _5055_/C _5049_/C _5058_/C _5180_/B VGND VGND VPWR VPWR _5056_/B
+ sky130_fd_sc_hd__a32oi_2
XFILLER_85_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5998__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1449 hold25/X VGND VGND VPWR VPWR hold1449/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4005_ _4005_/A _4058_/A _4058_/B _7073_/Q VGND VGND VPWR VPWR _4006_/B sky130_fd_sc_hd__nor4_1
XANTENNA__4446__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5214__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5956_ _5965_/A _5956_/B _5956_/C VGND VGND VPWR VPWR _5964_/S sky130_fd_sc_hd__and3_4
XANTENNA__4422__A1 _4422_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4907_ _4933_/B _4907_/B _5260_/D VGND VGND VPWR VPWR _4907_/X sky130_fd_sc_hd__and3_1
XANTENNA__5785__B _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4973__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5887_ _5887_/A0 _5986_/A1 hold91/X VGND VGND VPWR VPWR _5887_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4181__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7626_ _7627_/CLK _7626_/D fanout690/X VGND VGND VPWR VPWR _7626_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6175__A1 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4838_ _4910_/D _4840_/D _5282_/A _4839_/B VGND VGND VPWR VPWR _4841_/B sky130_fd_sc_hd__and4_1
XANTENNA__6175__B2 _7354_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3528__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7557_ _7581_/CLK _7557_/D fanout716/X VGND VGND VPWR VPWR _7557_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_5_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4769_ _5404_/C _5410_/B VGND VGND VPWR VPWR _4769_/Y sky130_fd_sc_hd__nand2_1
X_6508_ _6429_/C _7577_/Q _6408_/C _6507_/X VGND VGND VPWR VPWR _6508_/X sky130_fd_sc_hd__a31o_1
X_7488_ _7491_/CLK _7488_/D fanout719/X VGND VGND VPWR VPWR _7488_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6478__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6439_ _7399_/Q _6409_/X _6437_/X _6438_/X VGND VGND VPWR VPWR _6439_/X sky130_fd_sc_hd__a211o_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3330 _7620_/Q VGND VGND VPWR VPWR _6599_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3341 _4120_/X VGND VGND VPWR VPWR _7075_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3352 _6896_/Q VGND VGND VPWR VPWR _4051_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__buf_6
Xhold3363 _7585_/Q VGND VGND VPWR VPWR _6012_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3700__A3 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3374 _6908_/Q VGND VGND VPWR VPWR _4005_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__buf_2
Xhold2640 _4454_/X VGND VGND VPWR VPWR hold706/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2651 _7171_/Q VGND VGND VPWR VPWR hold719/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2662 _7279_/Q VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5989__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2673 _7335_/Q VGND VGND VPWR VPWR hold519/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4864__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2684 hold669/X VGND VGND VPWR VPWR _4478_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2695 hold811/X VGND VGND VPWR VPWR _5880_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1950 hold172/X VGND VGND VPWR VPWR _5987_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1961 _5703_/X VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1972 hold463/X VGND VGND VPWR VPWR _4493_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1983 _5952_/X VGND VGND VPWR VPWR hold295/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1994 _4448_/X VGND VGND VPWR VPWR hold273/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6901__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5205__A3 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3927__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6705__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 _3801_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6469__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4758__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3662__C _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4266__S _4270_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6641__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2010_A _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5810_ _5810_/A0 _5999_/A1 _5811_/S VGND VGND VPWR VPWR _5810_/X sky130_fd_sc_hd__mux2_1
X_6790_ _3643_/Y _6790_/A1 _6792_/S VGND VGND VPWR VPWR _7634_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4404__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5741_ _5741_/A0 _5975_/A0 _5748_/S VGND VGND VPWR VPWR _5741_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4955__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5672_ _5951_/A1 _5672_/A1 _5676_/S VGND VGND VPWR VPWR _5672_/X sky130_fd_sc_hd__mux2_1
X_7411_ _7472_/CLK _7411_/D fanout719/X VGND VGND VPWR VPWR _7411_/Q sky130_fd_sc_hd__dfrtp_4
X_4623_ _5127_/A _5222_/A _5059_/A VGND VGND VPWR VPWR _4841_/A sky130_fd_sc_hd__and3_1
XANTENNA__5825__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3915__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7342_ _7579_/CLK _7342_/D fanout731/X VGND VGND VPWR VPWR _7342_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ _5914_/A1 _4554_/A1 _4556_/S VGND VGND VPWR VPWR _4554_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5380__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold502 hold502/A VGND VGND VPWR VPWR _7384_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold513 hold513/A VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold524 _4211_/X VGND VGND VPWR VPWR _6926_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3505_ _3505_/A hold38/X _3505_/C hold88/X VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__nor4_1
X_7273_ _7314_/CLK _7273_/D _4079_/A VGND VGND VPWR VPWR _7273_/Q sky130_fd_sc_hd__dfrtp_1
Xhold535 hold535/A VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4485_ _4485_/A _5640_/D VGND VGND VPWR VPWR _4490_/S sky130_fd_sc_hd__nand2_4
Xhold546 hold546/A VGND VGND VPWR VPWR _6953_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold568 hold568/A VGND VGND VPWR VPWR _7403_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold579 hold579/A VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6224_ _7468_/Q _6087_/X _6220_/X _6221_/X _6223_/X VGND VGND VPWR VPWR _6224_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_89_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3436_ _7354_/Q VGND VGND VPWR VPWR _3436_/Y sky130_fd_sc_hd__inv_2
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _7321_/Q _6119_/D _6081_/X _6075_/X _7425_/Q VGND VGND VPWR VPWR _6155_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 hold2889/X VGND VGND VPWR VPWR hold2890/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3694__A2 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5561_/A1 _4814_/Y _5509_/A3 _5104_/Y VGND VGND VPWR VPWR _5111_/C sky130_fd_sc_hd__o31ai_1
Xhold1213 hold2928/X VGND VGND VPWR VPWR _6990_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _7589_/Q _7588_/Q _6120_/B VGND VGND VPWR VPWR _6086_/X sky130_fd_sc_hd__and3_2
Xhold1224 hold2894/X VGND VGND VPWR VPWR hold2895/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1235 _5870_/X VGND VGND VPWR VPWR _7466_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1246 hold2929/X VGND VGND VPWR VPWR hold2930/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1257 hold2937/X VGND VGND VPWR VPWR hold2938/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5037_ _5037_/A _5037_/B _5037_/C VGND VGND VPWR VPWR _5039_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6632__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1268 _4512_/X VGND VGND VPWR VPWR _7164_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1279 hold3237/X VGND VGND VPWR VPWR hold3238/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6396__A1 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6988_ _7497_/CLK _6988_/D fanout693/X VGND VGND VPWR VPWR _6988_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6396__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5939_ _5939_/A0 _5975_/A0 _5946_/S VGND VGND VPWR VPWR _5939_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4850__D _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7609_ _7610_/CLK _7609_/D fanout693/X VGND VGND VPWR VPWR _7609_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6699__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6420__A _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5371__A2 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input162_A wb_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3482__C _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6320__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5123__A2 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR _4564_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR _5071_/A sky130_fd_sc_hd__buf_2
Xhold3160 hold3160/A VGND VGND VPWR VPWR _4516_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR input122/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3171 _7001_/Q VGND VGND VPWR VPWR hold3171/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3685__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR _6805_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3182 _4546_/X VGND VGND VPWR VPWR hold3182/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR _6812_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3193 _7016_/Q VGND VGND VPWR VPWR hold3193/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR _6817_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR _6825_/A3 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2470 hold873/X VGND VGND VPWR VPWR _4186_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input23_A mask_rev_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2481 _7380_/Q VGND VGND VPWR VPWR hold949/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6623__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2492 hold639/X VGND VGND VPWR VPWR _5925_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4634__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1780 _7446_/Q VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1791 hold37/X VGND VGND VPWR VPWR _3470_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6387__A1 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4398__A0 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6139__A1 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5645__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5898__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3673__B _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4270_ _4270_/A0 _5817_/A1 _4270_/S VGND VGND VPWR VPWR _4270_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3676__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4873__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6614__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6911_ _7263_/CLK _6911_/D fanout688/X VGND VGND VPWR VPWR _6911_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6842_ _6861_/A _6869_/B VGND VGND VPWR VPWR _6842_/X sky130_fd_sc_hd__and2_1
XANTENNA__4389__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6773_ _6773_/A _6773_/B _6773_/C _6773_/D VGND VGND VPWR VPWR _6774_/C sky130_fd_sc_hd__nor4_2
X_3985_ _7648_/A _3933_/A _3598_/B _3984_/X VGND VGND VPWR VPWR _3985_/X sky130_fd_sc_hd__a31o_1
XANTENNA_hold2761_A _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5724_ _5724_/A0 _5949_/A1 _5730_/S VGND VGND VPWR VPWR _5724_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3600__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5655_ _5952_/A1 _5655_/A1 _5657_/S VGND VGND VPWR VPWR _5655_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3864__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4606_ _4879_/D _4747_/B VGND VGND VPWR VPWR _5387_/B sky130_fd_sc_hd__nor2_8
XFILLER_175_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5586_ _5736_/A1 _5586_/A1 _5586_/S VGND VGND VPWR VPWR _5586_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6550__A1 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5353__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7325_ _7582_/CLK _7325_/D fanout716/X VGND VGND VPWR VPWR _7325_/Q sky130_fd_sc_hd__dfrtp_2
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold321 hold321/A VGND VGND VPWR VPWR _7019_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4537_ _4555_/A0 _4537_/A1 _4538_/S VGND VGND VPWR VPWR _4537_/X sky130_fd_sc_hd__mux2_1
Xhold332 hold332/A VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold343 _3576_/X VGND VGND VPWR VPWR _4521_/B sky130_fd_sc_hd__clkbuf_2
Xhold354 hold354/A VGND VGND VPWR VPWR _6965_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7256_ _7266_/CLK _7256_/D fanout694/X VGND VGND VPWR VPWR _7256_/Q sky130_fd_sc_hd__dfrtp_2
Xhold365 _4078_/B VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__buf_6
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4468_ _5912_/A1 _4468_/A1 _4472_/S VGND VGND VPWR VPWR _4468_/X sky130_fd_sc_hd__mux2_1
Xhold387 hold387/A VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6302__B2 _7026_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold398 hold398/A VGND VGND VPWR VPWR _7315_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6207_ _6204_/X _6205_/X _6206_/X _6144_/C VGND VGND VPWR VPWR _6207_/X sky130_fd_sc_hd__o31a_1
X_3419_ _7490_/Q VGND VGND VPWR VPWR _3419_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7187_ _7268_/CLK _7187_/D _6869_/A VGND VGND VPWR VPWR _7187_/Q sky130_fd_sc_hd__dfrtp_4
X_4399_ _5817_/A1 _4399_/A1 _4399_/S VGND VGND VPWR VPWR _4399_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_73_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _7368_/Q _6388_/A3 _6136_/X _6137_/X _6135_/X VGND VGND VPWR VPWR _6138_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1010 _5966_/X VGND VGND VPWR VPWR _7551_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1021 hold3034/X VGND VGND VPWR VPWR _7383_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1032 hold3082/X VGND VGND VPWR VPWR hold3083/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1043 hold3069/X VGND VGND VPWR VPWR hold3070/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6605__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1054 hold2827/X VGND VGND VPWR VPWR hold2828/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6069_ _6751_/S _4117_/B _6067_/X VGND VGND VPWR VPWR _6069_/X sky130_fd_sc_hd__a21o_1
XTAP_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1065 hold3094/X VGND VGND VPWR VPWR _7487_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1076 hold2981/X VGND VGND VPWR VPWR hold1076/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 hold1087/A VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 hold2975/X VGND VGND VPWR VPWR hold1098/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6415__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6369__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6384__A4 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6541__A1 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6541__B2 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__B _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4607__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3830__A2 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6044__B _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3770_ _7029_/Q _4352_/A _4352_/B _3649_/X _7069_/Q VGND VGND VPWR VPWR _3770_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5440_ _5199_/C _5058_/C _5439_/X VGND VGND VPWR VPWR _5506_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__6532__A1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6532__B2 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5371_ _5059_/B _5404_/D _4966_/A _5248_/A VGND VGND VPWR VPWR _5371_/X sky130_fd_sc_hd__o211a_1
X_7110_ _7111_/CLK _7110_/D fanout751/X VGND VGND VPWR VPWR _7110_/Q sky130_fd_sc_hd__dfrtp_4
X_4322_ _4322_/A _5619_/C VGND VGND VPWR VPWR _4327_/S sky130_fd_sc_hd__nand2_4
XFILLER_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold31_A hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7041_ _7201_/CLK _7041_/D _6839_/A VGND VGND VPWR VPWR _7041_/Q sky130_fd_sc_hd__dfrtp_4
X_4253_ _4253_/A0 _5986_/A1 _4258_/S VGND VGND VPWR VPWR _4253_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4184_ _4184_/A0 _4553_/A0 _4190_/S VGND VGND VPWR VPWR _4184_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3821__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_7_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_6825_ _7110_/Q _6824_/C _6825_/A3 _6824_/X VGND VGND VPWR VPWR _6825_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3968_ _7279_/Q _3558_/X _4394_/A _7061_/Q _3967_/X VGND VGND VPWR VPWR _3968_/X
+ sky130_fd_sc_hd__a221o_1
X_6756_ _7065_/Q _6574_/B _6441_/X _6419_/D _7005_/Q VGND VGND VPWR VPWR _6756_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6771__B2 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5707_ _5995_/A1 _5707_/A1 _5712_/S VGND VGND VPWR VPWR _5707_/X sky130_fd_sc_hd__mux2_1
X_6687_ _6968_/Q _6420_/A _6457_/X _7062_/Q _6686_/X VGND VGND VPWR VPWR _6687_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3899_ _7488_/Q _5893_/A _5581_/A _7210_/Q _3898_/X VGND VGND VPWR VPWR _3899_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5638_ _5969_/A1 _5638_/A1 _5639_/S VGND VGND VPWR VPWR _5638_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4534__A0 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5569_ _5569_/A _5569_/B _5569_/C VGND VGND VPWR VPWR _5569_/X sky130_fd_sc_hd__and3_1
XFILLER_191_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3888__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold140 hold140/A VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7308_ _7365_/CLK _7308_/D fanout713/X VGND VGND VPWR VPWR _7308_/Q sky130_fd_sc_hd__dfrtp_4
Xhold151 hold151/A VGND VGND VPWR VPWR _7394_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold173 hold173/A VGND VGND VPWR VPWR _7570_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold195 hold195/A VGND VGND VPWR VPWR _7401_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7239_ _7327_/CLK _7239_/D fanout703/X VGND VGND VPWR VPWR _7239_/Q sky130_fd_sc_hd__dfstp_1
Xfanout620 _7592_/Q VGND VGND VPWR VPWR _6075_/A sky130_fd_sc_hd__buf_6
Xfanout631 _4007_/B VGND VGND VPWR VPWR _4025_/A sky130_fd_sc_hd__buf_6
XFILLER_120_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout664 _4704_/Y VGND VGND VPWR VPWR _5068_/B sky130_fd_sc_hd__buf_4
Xfanout675 _4596_/X VGND VGND VPWR VPWR _5091_/A sky130_fd_sc_hd__buf_12
Xfanout686 _4128_/B VGND VGND VPWR VPWR _6864_/A sky130_fd_sc_hd__buf_4
Xfanout697 fanout750/X VGND VGND VPWR VPWR _6872_/A sky130_fd_sc_hd__buf_6
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input125_A wb_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5262__B2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3488__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7079__RESET_B fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6762__B2 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input90_A spimemio_flash_io2_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6514__A1 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f__1111_ clkbuf_0__1111_/X VGND VGND VPWR VPWR _3734_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6278__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3670__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5253__A1 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4940_ _4954_/A _5453_/A _5260_/D _4940_/D VGND VGND VPWR VPWR _4941_/B sky130_fd_sc_hd__and4_1
XFILLER_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3803__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4871_ _4747_/B _4945_/A _4887_/B _4879_/D VGND VGND VPWR VPWR _4871_/X sky130_fd_sc_hd__and4bb_1
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6610_ _7365_/Q _6462_/X _6607_/X _6609_/X VGND VGND VPWR VPWR _6610_/X sky130_fd_sc_hd__a211o_1
X_3822_ _7159_/Q _4376_/B _4352_/B _3647_/X _7169_/Q VGND VGND VPWR VPWR _3822_/X
+ sky130_fd_sc_hd__a32o_1
X_7590_ _7594_/CLK _7590_/D fanout694/X VGND VGND VPWR VPWR _7590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3567__A1 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6541_ _7394_/Q _6420_/C _6421_/X _7322_/Q _6540_/X VGND VGND VPWR VPWR _6544_/C
+ sky130_fd_sc_hd__a221o_1
X_3753_ input95/X _4431_/A _4265_/B _3526_/X _7506_/Q VGND VGND VPWR VPWR _3753_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_186_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4303__A _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6472_ wire352/X _6471_/Y _7279_/Q _6431_/Y VGND VGND VPWR VPWR _6472_/X sky130_fd_sc_hd__o2bb2a_1
X_3684_ _7283_/Q _3590_/C _4265_/B _5848_/A _7451_/Q VGND VGND VPWR VPWR _3684_/X
+ sky130_fd_sc_hd__a32o_1
X_5423_ _5423_/A _5423_/B VGND VGND VPWR VPWR _5438_/C sky130_fd_sc_hd__and2_1
XFILLER_145_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput201 _3412_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
XANTENNA__5833__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput212 _3436_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
XFILLER_145_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2724_A _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput223 _7660_/X VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput234 _4146_/X VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
X_5354_ _5065_/A _5077_/B _5248_/C _5213_/X _5350_/X VGND VGND VPWR VPWR _5355_/D
+ sky130_fd_sc_hd__a311oi_4
XFILLER_160_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput245 _4151_/X VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
Xoutput256 _7233_/Q VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput267 _7230_/Q VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
XANTENNA__6269__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4305_ _4305_/A0 _5645_/A0 _4308_/S VGND VGND VPWR VPWR _4305_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3861__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput278 _7237_/Q VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
Xoutput289 _6923_/Q VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
X_5285_ _5134_/A _5059_/B _5399_/D _5284_/X VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5134__A _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7024_ _7497_/CLK _7024_/D fanout693/X VGND VGND VPWR VPWR _7024_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4236_ _5652_/A1 _5949_/A1 _4248_/S VGND VGND VPWR VPWR _4236_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4295__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4167_ _7601_/Q _7251_/Q _7255_/Q VGND VGND VPWR VPWR _4167_/X sky130_fd_sc_hd__mux2_8
XFILLER_83_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4098_ _4098_/A1 _4011_/X _4123_/C _4058_/A _4010_/Y VGND VGND VPWR VPWR _7071_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_83_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout542_A _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_csclk _7416_/CLK VGND VGND VPWR VPWR _7179_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ _4427_/D _6808_/A2 _6808_/B1 _4427_/C VGND VGND VPWR VPWR _6808_/X sky130_fd_sc_hd__a22o_1
XFILLER_169_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6744__A1 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6744__B2 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6739_ _7145_/Q _6468_/X _6734_/X _6736_/X _6738_/X VGND VGND VPWR VPWR _6749_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_7_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5743__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3730__B2 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3490__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout450 _5938_/B VGND VGND VPWR VPWR _5722_/B sky130_fd_sc_hd__buf_4
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout461 _6106_/X VGND VGND VPWR VPWR _6267_/B1 sky130_fd_sc_hd__buf_4
Xfanout472 _6433_/X VGND VGND VPWR VPWR _6574_/C sky130_fd_sc_hd__buf_8
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6680__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout483 _6402_/Y VGND VGND VPWR VPWR _6747_/C sky130_fd_sc_hd__buf_6
XANTENNA__4883__A _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout494 _6574_/B VGND VGND VPWR VPWR _6466_/C sky130_fd_sc_hd__buf_8
XFILLER_59_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6432__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4107__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6499__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold909 hold909/A VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5171__B1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3721__A1 input16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4269__S _4270_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5070_ _4810_/C _5115_/C _5260_/D _5134_/A VGND VGND VPWR VPWR _5070_/X sky130_fd_sc_hd__a22o_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 hold166/X VGND VGND VPWR VPWR _5627_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4021_ _6905_/Q _6904_/Q _4025_/B hold44/A VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__a31o_1
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5972_ _5972_/A0 _5972_/A1 _5973_/S VGND VGND VPWR VPWR _5972_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4923_ _5453_/A _4954_/C _4933_/A _4970_/C VGND VGND VPWR VPWR _5444_/C sky130_fd_sc_hd__nand4_1
XANTENNA__5828__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7642_ _7646_/CLK _7642_/D fanout753/X VGND VGND VPWR VPWR _7642_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4854_ _4622_/Y _4654_/Y _4748_/Y _4427_/D VGND VGND VPWR VPWR _4854_/X sky130_fd_sc_hd__o31a_2
XANTENNA__3856__B _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3805_ input97/X _4431_/A _4265_/B _5634_/A _7258_/Q VGND VGND VPWR VPWR _3805_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7573_ _7573_/CLK hold73/X fanout733/X VGND VGND VPWR VPWR _7573_/Q sky130_fd_sc_hd__dfrtp_4
X_4785_ _4700_/Y _4707_/Y _4784_/Y _4781_/Y VGND VGND VPWR VPWR _4791_/B sky130_fd_sc_hd__o211ai_1
XFILLER_193_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3736_ _7218_/Q _3996_/A _3734_/Y _3735_/X VGND VGND VPWR VPWR _7218_/D sky130_fd_sc_hd__a22o_2
X_6524_ _7530_/Q _6058_/X _6409_/X _7402_/Q VGND VGND VPWR VPWR _6524_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3960__A1 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3667_ _5640_/B _5596_/A _4346_/C VGND VGND VPWR VPWR _3667_/X sky130_fd_sc_hd__and3_4
X_6455_ _6463_/A _6455_/B _6466_/D VGND VGND VPWR VPWR _6455_/X sky130_fd_sc_hd__and3_4
XFILLER_109_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5406_ _5282_/A _5011_/B _5113_/A VGND VGND VPWR VPWR _5406_/Y sky130_fd_sc_hd__a21oi_2
X_6386_ _6878_/Q _6112_/X _6121_/X _6992_/Q VGND VGND VPWR VPWR _6386_/X sky130_fd_sc_hd__a22o_1
X_3598_ _5590_/A _3598_/B _5596_/B VGND VGND VPWR VPWR _3598_/X sky130_fd_sc_hd__and3_2
XANTENNA__3712__A1 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5337_ _5034_/B _5053_/C _5328_/X _5336_/X VGND VGND VPWR VPWR _5337_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2800 _4270_/X VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2811 hold995/X VGND VGND VPWR VPWR _4483_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5268_ _5255_/X _4774_/Y _5267_/X _5266_/Y VGND VGND VPWR VPWR _5268_/X sky130_fd_sc_hd__o211a_1
Xhold2822 hold871/X VGND VGND VPWR VPWR _5814_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2833 _7367_/Q VGND VGND VPWR VPWR hold2833/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5465__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2844 _4247_/X VGND VGND VPWR VPWR hold2844/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2855 _7652_/A VGND VGND VPWR VPWR hold2855/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2866 _7289_/Q VGND VGND VPWR VPWR hold2866/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7007_ _7191_/CLK _7007_/D fanout700/X VGND VGND VPWR VPWR _7007_/Q sky130_fd_sc_hd__dfrtp_4
X_4219_ hold261/X _5976_/A0 _4231_/S VGND VGND VPWR VPWR _4219_/X sky130_fd_sc_hd__mux2_1
Xhold2877 _7226_/Q VGND VGND VPWR VPWR hold2877/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5199_ _4888_/C _5342_/A _5199_/C _5342_/C VGND VGND VPWR VPWR _5200_/B sky130_fd_sc_hd__nand4b_2
Xhold2888 _4417_/X VGND VGND VPWR VPWR hold2888/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2899 _4325_/X VGND VGND VPWR VPWR hold2899/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6407__B _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4440__A2 hold365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5965__C hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6423__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6717__B2 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_762 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3951__A1 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3951__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4597__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input53_A mgmt_gpio_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6248__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6653__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7094__RESET_B fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output307_A _4134_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5648__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5875__C _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6184__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4195__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4570_ _4831_/A _4909_/D _4772_/B VGND VGND VPWR VPWR _4570_/Y sky130_fd_sc_hd__nand3_4
X_3521_ _5590_/A _4328_/A _3562_/C VGND VGND VPWR VPWR _3521_/X sky130_fd_sc_hd__and3_4
XANTENNA__3942__A1 input61/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4788__A _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold706 hold706/A VGND VGND VPWR VPWR _7116_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold717 hold717/A VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap425 _4696_/B VGND VGND VPWR VPWR _5138_/C sky130_fd_sc_hd__clkbuf_2
Xhold728 hold728/A VGND VGND VPWR VPWR _7097_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6240_ _7333_/Q _6136_/B _6116_/A _6112_/C VGND VGND VPWR VPWR _6240_/X sky130_fd_sc_hd__a31o_1
XANTENNA_hold2255_A _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3452_ _4028_/A0 _4025_/A hold44/X VGND VGND VPWR VPWR _3452_/X sky130_fd_sc_hd__a21o_1
Xhold739 hold739/A VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6171_ _7298_/Q _6384_/A4 _6270_/C1 _6079_/X _7330_/Q VGND VGND VPWR VPWR _6171_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5122_ _5061_/X _5122_/B _5122_/C VGND VGND VPWR VPWR _5122_/Y sky130_fd_sc_hd__nand3b_1
Xhold2107 hold507/X VGND VGND VPWR VPWR _4222_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2118 _6938_/Q VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2129 hold2129/A VGND VGND VPWR VPWR _5910_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1406 hold1463/X VGND VGND VPWR VPWR hold1464/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6644__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5053_ _5063_/D _5203_/A _5053_/C VGND VGND VPWR VPWR _5058_/C sky130_fd_sc_hd__and3_4
Xhold1417 hold1417/A VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1428 hold1428/A VGND VGND VPWR VPWR _5627_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1439 _4199_/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4004_ _4004_/A _4006_/A VGND VGND VPWR VPWR _6909_/D sky130_fd_sc_hd__xor2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4670__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5955_ _5955_/A0 _5955_/A1 _5955_/S VGND VGND VPWR VPWR _5955_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4970__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _4906_/B _5185_/C _4906_/D VGND VGND VPWR VPWR _4906_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3630__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5886_ _5886_/A0 _5922_/A0 hold91/X VGND VGND VPWR VPWR _5886_/X sky130_fd_sc_hd__mux2_1
X_7625_ _7625_/CLK _7625_/D fanout690/X VGND VGND VPWR VPWR _7625_/Q sky130_fd_sc_hd__dfrtp_1
X_4837_ _4837_/A _4837_/B _4837_/C VGND VGND VPWR VPWR _4841_/C sky130_fd_sc_hd__nand3_1
XFILLER_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6175__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4186__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout505_A _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7556_ _7556_/CLK _7556_/D fanout732/X VGND VGND VPWR VPWR _7556_/Q sky130_fd_sc_hd__dfrtp_4
X_4768_ _4860_/A _4768_/B VGND VGND VPWR VPWR _4768_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_147_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6507_ _7433_/Q _6747_/B _6468_/C _6408_/A _7553_/Q VGND VGND VPWR VPWR _6507_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3719_ _7146_/Q _4364_/A _5938_/B _4515_/B _3718_/X VGND VGND VPWR VPWR _3719_/X
+ sky130_fd_sc_hd__a41o_1
X_7487_ _7576_/CLK _7487_/D fanout718/X VGND VGND VPWR VPWR _7487_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_106_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4699_ _4910_/D _4856_/A _4888_/B VGND VGND VPWR VPWR _5282_/B sky130_fd_sc_hd__nor3_4
XFILLER_146_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6438_ _7391_/Q _6420_/C _6419_/A _7543_/Q VGND VGND VPWR VPWR _6438_/X sky130_fd_sc_hd__a22o_1
XFILLER_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3320 _7614_/Q VGND VGND VPWR VPWR _6401_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6369_ _7004_/Q _6097_/B _6120_/B _6379_/B1 _7125_/Q VGND VGND VPWR VPWR _6369_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3331 _7608_/Q VGND VGND VPWR VPWR _6261_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_22_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7185_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold3342 _7101_/Q VGND VGND VPWR VPWR _4114_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3353 _6931_/Q VGND VGND VPWR VPWR hold3353/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3364 _6893_/Q VGND VGND VPWR VPWR _4057_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2630 _6878_/Q VGND VGND VPWR VPWR hold703/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3375 _6895_/Q VGND VGND VPWR VPWR _4053_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6635__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2641 _7139_/Q VGND VGND VPWR VPWR hold891/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__buf_8
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2652 hold719/X VGND VGND VPWR VPWR _4520_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2663 hold505/X VGND VGND VPWR VPWR _5660_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2674 hold519/X VGND VGND VPWR VPWR _5723_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1940 _7582_/Q VGND VGND VPWR VPWR hold184/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2685 _4478_/X VGND VGND VPWR VPWR hold670/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4110__A1 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1951 _5987_/X VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__clkbuf_2
Xhold2696 _7184_/Q VGND VGND VPWR VPWR hold983/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1962 _7282_/Q VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1973 _7283_/Q VGND VGND VPWR VPWR hold300/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_37_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7578_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1984 _6875_/Q VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1995 _7313_/Q VGND VGND VPWR VPWR hold427/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1989_A _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5610__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clkbuf_0_mgmt_gpio_in[4]/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5695__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6166__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5992__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6600__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_8 _3859_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6469__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5216__B _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output257_A _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5931__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_532 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5429__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6626__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6047__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5601__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5740_ _5740_/A _5956_/B _5992_/D VGND VGND VPWR VPWR _5748_/S sky130_fd_sc_hd__and3_4
XANTENNA__3612__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4955__A3 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5671_ _5815_/A1 _5671_/A1 _5676_/S VGND VGND VPWR VPWR _5671_/X sky130_fd_sc_hd__mux2_1
X_7410_ _7421_/CLK _7410_/D fanout715/X VGND VGND VPWR VPWR _7410_/Q sky130_fd_sc_hd__dfrtp_4
X_4622_ _4870_/A _4657_/A VGND VGND VPWR VPWR _4622_/Y sky130_fd_sc_hd__nand2_8
XFILLER_175_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7341_ _7478_/CLK _7341_/D fanout714/X VGND VGND VPWR VPWR _7341_/Q sky130_fd_sc_hd__dfrtp_4
X_4553_ _4553_/A0 _4553_/A1 _4556_/S VGND VGND VPWR VPWR _4553_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5380__A3 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold503 hold503/A VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold514 _5895_/X VGND VGND VPWR VPWR _7488_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold525 hold525/A VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3504_ _3504_/A _3504_/B VGND VGND VPWR VPWR _3504_/Y sky130_fd_sc_hd__nor2_1
X_4484_ _4484_/A0 _5853_/A0 _4484_/S VGND VGND VPWR VPWR _4484_/X sky130_fd_sc_hd__mux2_1
X_7272_ _7314_/CLK _7272_/D _4079_/A VGND VGND VPWR VPWR _7272_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6314__C1 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold536 hold536/A VGND VGND VPWR VPWR _7547_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold547 hold547/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4668__D _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold558 hold558/A VGND VGND VPWR VPWR _7387_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold569 hold569/A VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6223_ _7532_/Q _6092_/X _6112_/X _7484_/Q _6222_/X VGND VGND VPWR VPWR _6223_/X
+ sky130_fd_sc_hd__a221o_1
X_3435_ _7362_/Q VGND VGND VPWR VPWR _3435_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _7353_/Q _6099_/X _6110_/X _7433_/Q _6153_/X VGND VGND VPWR VPWR _6157_/B
+ sky130_fd_sc_hd__a221oi_2
XFILLER_98_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3694__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 _5626_/X VGND VGND VPWR VPWR _7252_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5105_ _5107_/C _5399_/C _5453_/C VGND VGND VPWR VPWR _5105_/X sky130_fd_sc_hd__and3_1
Xhold1214 hold2869/X VGND VGND VPWR VPWR hold2870/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _7590_/Q _6121_/A _6110_/A _6099_/D VGND VGND VPWR VPWR _6085_/X sky130_fd_sc_hd__and4b_4
Xhold1225 hold2896/X VGND VGND VPWR VPWR _7458_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 hold2940/X VGND VGND VPWR VPWR hold2941/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1247 _4506_/X VGND VGND VPWR VPWR _7159_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5036_ _4821_/Y _4862_/X _4865_/Y _4992_/Y _5035_/Y VGND VGND VPWR VPWR _5037_/A
+ sky130_fd_sc_hd__o311a_1
Xhold1258 hold2939/X VGND VGND VPWR VPWR _7018_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1269 hold2961/X VGND VGND VPWR VPWR hold2962/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5840__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout455_A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ _7630_/CLK _6987_/D VGND VGND VPWR VPWR _6987_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6396__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout622_A _7591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3603__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5938_ _5938_/A _5938_/B _5938_/C _5956_/C VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__and4_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5869_ _5869_/A0 _5986_/A1 _5874_/S VGND VGND VPWR VPWR _5869_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7608_ _7621_/CLK _7608_/D fanout711/X VGND VGND VPWR VPWR _7608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3906__A1 input15/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7539_ _7539_/CLK _7539_/D fanout708/X VGND VGND VPWR VPWR _7539_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3906__B2 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6420__B _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6320__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input155_A wb_dat_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4875__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR _4564_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3150 _7503_/Q VGND VGND VPWR VPWR hold3150/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR _5004_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__6608__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3161 _4516_/X VGND VGND VPWR VPWR hold3161/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR input123/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3172 hold3172/A VGND VGND VPWR VPWR _4323_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3685__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR _6808_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3183 _7142_/Q VGND VGND VPWR VPWR hold3183/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR _6814_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3194 hold3194/A VGND VGND VPWR VPWR _4341_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2460 hold915/X VGND VGND VPWR VPWR _4511_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR _6820_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR _6795_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2471 _4186_/X VGND VGND VPWR VPWR hold874/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2482 hold949/X VGND VGND VPWR VPWR _5773_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2493 _5925_/X VGND VGND VPWR VPWR hold640/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1770 _5727_/X VGND VGND VPWR VPWR hold119/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5292__C1 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5831__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4634__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input16_A mask_rev_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1781 hold101/X VGND VGND VPWR VPWR _5847_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6899__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1792 _3470_/X VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6387__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6139__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4131__A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6311__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4428__A_N _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3676__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold2218_A _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6614__A3 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5822__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6910_ _7075_/CLK _6910_/D _6860_/X VGND VGND VPWR VPWR _6910_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3833__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6841_ _6861_/A _6869_/B VGND VGND VPWR VPWR _6841_/X sky130_fd_sc_hd__and2_1
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5586__A0 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6772_ _6971_/Q _6420_/A _6422_/X _6966_/Q _6771_/X VGND VGND VPWR VPWR _6773_/D
+ sky130_fd_sc_hd__a221o_1
X_3984_ input4/X _3503_/X _3675_/X _7187_/Q VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__a22o_1
X_5723_ _5723_/A0 hold487/X _5730_/S VGND VGND VPWR VPWR _5723_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5836__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5654_ _5951_/A1 _5654_/A1 _5657_/S VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5889__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3864__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4605_ _5260_/A _5260_/B VGND VGND VPWR VPWR _4605_/Y sky130_fd_sc_hd__nand2_8
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5585_ _5585_/A0 _5585_/A1 _5586_/S VGND VGND VPWR VPWR _5585_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6550__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5353__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold300 hold300/A VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7324_ _7478_/CLK _7324_/D fanout715/X VGND VGND VPWR VPWR _7324_/Q sky130_fd_sc_hd__dfrtp_4
Xhold311 hold311/A VGND VGND VPWR VPWR _7508_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4536_ _5914_/A1 _4536_/A1 _4538_/S VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__mux2_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold333 _5751_/X VGND VGND VPWR VPWR _7360_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold344 _4524_/X VGND VGND VPWR VPWR _7174_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold355 hold355/A VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold366 hold366/A VGND VGND VPWR VPWR _7306_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7255_ _7255_/CLK _7255_/D fanout689/X VGND VGND VPWR VPWR _7255_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6302__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4467_ _4467_/A _4551_/D VGND VGND VPWR VPWR _4472_/S sky130_fd_sc_hd__nand2_4
Xhold377 hold377/A VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold388 hold388/A VGND VGND VPWR VPWR _7280_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6206_ _7299_/Q _6384_/A4 _6270_/C1 _6274_/A3 _7387_/Q VGND VGND VPWR VPWR _6206_/X
+ sky130_fd_sc_hd__a32o_1
X_3418_ _7498_/Q VGND VGND VPWR VPWR _3418_/Y sky130_fd_sc_hd__inv_2
X_4398_ _5625_/A1 _4398_/A1 _4399_/S VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__mux2_1
X_7186_ _7186_/CLK _7186_/D fanout725/X VGND VGND VPWR VPWR _7186_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input8_A mask_rev_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ _7288_/Q _6112_/B _6136_/C _6079_/X _7328_/Q VGND VGND VPWR VPWR _6137_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1000 hold3050/X VGND VGND VPWR VPWR _7262_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout572_A _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 hold3075/X VGND VGND VPWR VPWR hold3076/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1022 hold3051/X VGND VGND VPWR VPWR hold3052/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1033 hold3084/X VGND VGND VPWR VPWR _7527_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1044 hold3071/X VGND VGND VPWR VPWR _7056_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6605__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6649_/S _4117_/B _6067_/X VGND VGND VPWR VPWR _6068_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1055 hold2829/X VGND VGND VPWR VPWR _6943_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 hold2989/X VGND VGND VPWR VPWR hold1066/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5813__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1077 hold1077/A VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_100_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1088 hold2994/X VGND VGND VPWR VPWR hold1088/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5019_ _5024_/A1 _4669_/X _4974_/B _5180_/A _5158_/A VGND VGND VPWR VPWR _5021_/C
+ sky130_fd_sc_hd__o2111ai_2
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 hold1099/A VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6415__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6369__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5746__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1854_A _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6541__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3493__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4886__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4304__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3235_A _6941_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4607__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5804__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2290 _7278_/Q VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5280__A2 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3830__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4126__A _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3594__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6532__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4543__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5370_ _4659_/Y _5509_/A3 _5457_/B _5512_/A _5367_/Y VGND VGND VPWR VPWR _5370_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_160_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4321_ _3570_/Y _4321_/A1 _4321_/S VGND VGND VPWR VPWR _7000_/D sky130_fd_sc_hd__mux2_1
XFILLER_99_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5099__A2 _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7040_ _7179_/CLK _7040_/D fanout698/X VGND VGND VPWR VPWR _7040_/Q sky130_fd_sc_hd__dfrtp_4
X_4252_ hold261/X _5985_/A1 _4258_/S VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4183_ _4183_/A0 _7638_/Q _4429_/B VGND VGND VPWR VPWR _4183_/X sky130_fd_sc_hd__mux2_4
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6599__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3859__B _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3821__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6824_ _7111_/Q _6824_/B _6824_/C VGND VGND VPWR VPWR _6824_/X sky130_fd_sc_hd__and3_1
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6220__A1 _7348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6755_ _7166_/Q _6463_/X _6466_/X _7213_/Q _6754_/X VGND VGND VPWR VPWR _6755_/X
+ sky130_fd_sc_hd__a221o_1
X_3967_ _7051_/Q _3931_/B _5619_/B _3966_/X VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6771__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5706_ _5949_/A1 _5706_/A1 _5712_/S VGND VGND VPWR VPWR _5706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3585__A2 _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6686_ _7173_/Q _6747_/B _6747_/C _6425_/X _7017_/Q VGND VGND VPWR VPWR _6686_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout418_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3898_ _7173_/Q _4551_/B _4364_/B _3647_/X _7168_/Q VGND VGND VPWR VPWR _3898_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5637_ _5985_/A1 _5637_/A1 _5639_/S VGND VGND VPWR VPWR _5637_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5568_ _5568_/A _5568_/B _5568_/C VGND VGND VPWR VPWR _5569_/C sky130_fd_sc_hd__and3_1
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7307_ _7539_/CLK _7307_/D fanout708/X VGND VGND VPWR VPWR _7307_/Q sky130_fd_sc_hd__dfrtp_4
Xhold141 hold141/A VGND VGND VPWR VPWR _6954_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4519_ _4519_/A0 _5625_/A1 _4520_/S VGND VGND VPWR VPWR _4519_/X sky130_fd_sc_hd__mux2_1
Xhold152 hold152/A VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5499_ _5499_/A _5499_/B _5433_/C VGND VGND VPWR VPWR _5572_/A sky130_fd_sc_hd__nor3b_1
Xhold163 hold163/A VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold174 hold174/A VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6287__B2 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold185 hold185/A VGND VGND VPWR VPWR _7582_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7238_ _7238_/CLK _7238_/D fanout690/X VGND VGND VPWR VPWR _7238_/Q sky130_fd_sc_hd__dfstp_2
Xhold196 hold196/A VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout610 _3408_/Y VGND VGND VPWR VPWR _6623_/B1 sky130_fd_sc_hd__buf_4
Xfanout621 _7592_/Q VGND VGND VPWR VPWR _6080_/A sky130_fd_sc_hd__clkbuf_4
Xfanout632 _4058_/B VGND VGND VPWR VPWR _4007_/B sky130_fd_sc_hd__buf_4
XFILLER_132_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout643 _4888_/Y VGND VGND VPWR VPWR _5528_/A3 sky130_fd_sc_hd__clkbuf_16
X_7169_ _7181_/CLK _7169_/D fanout721/X VGND VGND VPWR VPWR _7169_/Q sky130_fd_sc_hd__dfstp_2
Xfanout676 _4583_/B VGND VGND VPWR VPWR _5494_/B2 sky130_fd_sc_hd__buf_12
Xfanout687 fanout750/X VGND VGND VPWR VPWR _4128_/B sky130_fd_sc_hd__buf_6
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold365_A _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout698 fanout702/X VGND VGND VPWR VPWR fanout698/X sky130_fd_sc_hd__buf_8
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5798__A0 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input118_A wb_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4470__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3488__C _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6762__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input83_A spimemio_flash_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6514__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3352_A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4525__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4289__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6450__A1 _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3803__A3 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4870_ _4870_/A _5065_/A _4907_/B VGND VGND VPWR VPWR _4877_/A sky130_fd_sc_hd__and3_4
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3821_ _7028_/Q _4346_/C _5632_/B _5848_/A _7449_/Q VGND VGND VPWR VPWR _3828_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6753__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__A2 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6540_ _7378_/Q _6408_/B _6460_/X _7386_/Q VGND VGND VPWR VPWR _6540_/X sky130_fd_sc_hd__a22o_1
X_3752_ _7530_/Q _3529_/X _3535_/X _7482_/Q _3751_/X VGND VGND VPWR VPWR _3759_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7472__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6471_ _6471_/A _6471_/B _6471_/C _6471_/D VGND VGND VPWR VPWR _6471_/Y sky130_fd_sc_hd__nor4_2
XFILLER_158_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4303__B _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3683_ _7228_/Q _3848_/A2 _5640_/C _5630_/S _7250_/Q VGND VGND VPWR VPWR _3683_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__6505__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5422_ _5422_/A _5422_/B _5496_/A _5422_/D VGND VGND VPWR VPWR _5422_/X sky130_fd_sc_hd__and4_1
Xoutput202 _3411_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 _4156_/X VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
XFILLER_145_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput224 _7661_/X VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
Xoutput235 _4147_/X VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
X_5353_ _4622_/Y _4726_/Y _4946_/Y _4898_/Y _5352_/Y VGND VGND VPWR VPWR _5355_/C
+ sky130_fd_sc_hd__o311a_1
Xoutput246 _4128_/Y VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
Xoutput257 _7234_/Q VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
X_4304_ _4304_/A0 _5948_/A1 _4308_/S VGND VGND VPWR VPWR _4304_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3861__C _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput268 _7231_/Q VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
XANTENNA__6269__B2 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput279 _7238_/Q VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5284_ _5399_/B _5081_/A _5115_/X _5281_/X VGND VGND VPWR VPWR _5284_/X sky130_fd_sc_hd__a31o_1
XFILLER_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7023_ _7497_/CLK _7023_/D fanout707/X VGND VGND VPWR VPWR _7023_/Q sky130_fd_sc_hd__dfstp_4
X_4235_ _4235_/A0 _4234_/X _4249_/S VGND VGND VPWR VPWR _4235_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4166_ _7599_/Q _7252_/Q _7255_/Q VGND VGND VPWR VPWR _4166_/X sky130_fd_sc_hd__mux2_4
XFILLER_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4097_ _4171_/B _4084_/X _4096_/X _4114_/B VGND VGND VPWR VPWR _7107_/D sky130_fd_sc_hd__a22o_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4692__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6807_ _6806_/X _6807_/A1 _6822_/S VGND VGND VPWR VPWR _7639_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4999_ _5339_/A _5183_/B _5018_/B VGND VGND VPWR VPWR _5026_/A sky130_fd_sc_hd__and3_1
XANTENNA__6744__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout702_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6738_ _7019_/Q _6425_/X _6457_/X _7064_/Q _6737_/X VGND VGND VPWR VPWR _6738_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6412__C _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6669_ _7122_/Q _6420_/C _6467_/X _7152_/Q _6668_/X VGND VGND VPWR VPWR _6669_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7141__RESET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4507__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5028__C _5028_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3730__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout440 _3502_/X VGND VGND VPWR VPWR _4455_/C sky130_fd_sc_hd__buf_6
Xfanout451 hold105/X VGND VGND VPWR VPWR _5938_/B sky130_fd_sc_hd__buf_12
Xfanout462 _6073_/X VGND VGND VPWR VPWR _6317_/C sky130_fd_sc_hd__buf_8
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout473 _6433_/X VGND VGND VPWR VPWR _6771_/A3 sky130_fd_sc_hd__clkbuf_8
Xfanout484 _6093_/X VGND VGND VPWR VPWR _6332_/C sky130_fd_sc_hd__buf_8
XFILLER_171_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout495 _6447_/B VGND VGND VPWR VPWR _6574_/B sky130_fd_sc_hd__buf_12
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3100_A _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6432__A1 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5934__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5171__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3721__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4020_ _4019_/X _4018_/X _4040_/A _3450_/B VGND VGND VPWR VPWR _6907_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5971_ _5971_/A0 _5998_/A1 _5973_/S VGND VGND VPWR VPWR _5971_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4922_ _4922_/A _4922_/B _4922_/C VGND VGND VPWR VPWR _4925_/A sky130_fd_sc_hd__nor3_1
X_7641_ _7641_/CLK _7641_/D fanout753/X VGND VGND VPWR VPWR _7641_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6187__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4853_ _5248_/A _5089_/D VGND VGND VPWR VPWR _4853_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5934__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3804_ _7521_/Q hold77/A _5776_/A _7385_/Q _3803_/X VGND VGND VPWR VPWR _3804_/X
+ sky130_fd_sc_hd__a221o_1
X_7572_ _7572_/CLK _7572_/D fanout736/X VGND VGND VPWR VPWR _7572_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4784_ _4811_/D _4784_/B VGND VGND VPWR VPWR _4784_/Y sky130_fd_sc_hd__nand2_1
X_6523_ _6522_/X _6523_/A1 _6573_/S VGND VGND VPWR VPWR _7617_/D sky130_fd_sc_hd__mux2_1
X_3735_ _3797_/A1 _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__o211a_1
X_6454_ _6466_/B _6463_/A _6466_/D _6466_/A VGND VGND VPWR VPWR _6454_/X sky130_fd_sc_hd__and4b_4
Xmgmt_gpio_31_buff_inst _4163_/X VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__clkbuf_8
X_3666_ _5612_/A _5596_/A _4346_/C VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__and3_4
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5405_ _4756_/X _5134_/X _5405_/C _5405_/D VGND VGND VPWR VPWR _5538_/B sky130_fd_sc_hd__and4bb_1
XFILLER_133_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5162__A1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6385_ _7065_/Q _6032_/Y _6081_/X _7196_/Q _6384_/X VGND VGND VPWR VPWR _6385_/X
+ sky130_fd_sc_hd__a221o_2
X_3597_ _7509_/Q _3872_/A2 _4527_/A _3535_/X _7485_/Q VGND VGND VPWR VPWR _3597_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_115_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5336_ _4996_/A _5034_/B _5328_/X _5335_/X VGND VGND VPWR VPWR _5336_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3712__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2801 _7180_/Q VGND VGND VPWR VPWR hold959/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2812 _4483_/X VGND VGND VPWR VPWR hold996/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5267_ _4803_/A _4775_/C _5516_/A3 _4717_/Y VGND VGND VPWR VPWR _5267_/X sky130_fd_sc_hd__o2bb2a_1
Xhold2823 _5814_/X VGND VGND VPWR VPWR hold872/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2834 hold2834/A VGND VGND VPWR VPWR _5759_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2845 _6959_/Q VGND VGND VPWR VPWR hold2845/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7006_ _7160_/CLK _7006_/D fanout700/X VGND VGND VPWR VPWR _7006_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6662__A1 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2856 hold2856/A VGND VGND VPWR VPWR _4245_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4218_ _4218_/A0 _4217_/X _4232_/S VGND VGND VPWR VPWR _4218_/X sky130_fd_sc_hd__mux2_1
Xhold2867 hold2867/A VGND VGND VPWR VPWR _5671_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2878 hold2878/A VGND VGND VPWR VPWR _5593_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5198_ _4672_/X _4893_/Y _4873_/X _5423_/A _5196_/X VGND VGND VPWR VPWR _5200_/A
+ sky130_fd_sc_hd__o311a_1
Xhold2889 _7252_/Q VGND VGND VPWR VPWR hold2889/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4149_ _6935_/Q _4076_/B _6899_/Q VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5217__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5622__C1 _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4976__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4440__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6717__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5925__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6193__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7214__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1934_A _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3951__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6350__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5055__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3703__A2 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4900__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input46_A mgmt_gpio_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4894__A _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_64_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3467__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6317__C _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3449__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire660 _4715_/Y VGND VGND VPWR VPWR _4765_/B sky130_fd_sc_hd__clkbuf_2
X_3520_ _5590_/A hold32/A _4328_/A VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__and3_4
Xhold707 hold707/A VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold718 hold718/A VGND VGND VPWR VPWR _7321_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold729 hold729/A VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5144__A1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3451_ hold44/X _4007_/B _3451_/B1 VGND VGND VPWR VPWR _3451_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_171_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2248_A _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6170_ _6170_/A1 _4116_/X _6067_/X _6169_/X VGND VGND VPWR VPWR _7604_/D sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_3_csclk _7416_/CLK VGND VGND VPWR VPWR _7164_/CLK sky130_fd_sc_hd__clkbuf_16
X_5121_ _4722_/Y _4880_/Y _4826_/Y _5495_/C1 VGND VGND VPWR VPWR _5122_/C sky130_fd_sc_hd__a211o_1
Xhold2108 _4222_/X VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2119 hold493/X VGND VGND VPWR VPWR _4228_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5447__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1407 hold1871/X VGND VGND VPWR VPWR hold1872/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1418 _6886_/Q VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5052_ _5052_/A _5052_/B _5052_/C VGND VGND VPWR VPWR _5056_/A sky130_fd_sc_hd__nor3_1
Xhold1429 _5602_/X VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3458__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4003_ _4003_/A _4003_/B VGND VGND VPWR VPWR _6910_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5954_ _5954_/A0 _5954_/A1 _5955_/S VGND VGND VPWR VPWR _5954_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4970__C _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4905_ _5065_/A _4954_/C _4907_/B _5260_/D VGND VGND VPWR VPWR _4906_/B sky130_fd_sc_hd__nand4_2
X_5885_ _5885_/A0 _5975_/A0 hold91/X VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7624_ _7625_/CLK _7624_/D fanout706/X VGND VGND VPWR VPWR _7624_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5907__A0 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4836_ _4836_/A _5260_/B _4836_/C _5089_/D VGND VGND VPWR VPWR _4837_/C sky130_fd_sc_hd__nand4_1
XFILLER_21_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3918__C1 _3917_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7555_ _7579_/CLK _7555_/D fanout731/X VGND VGND VPWR VPWR _7555_/Q sky130_fd_sc_hd__dfrtp_4
X_4767_ _4767_/A _4767_/B VGND VGND VPWR VPWR _5410_/B sky130_fd_sc_hd__nor2_8
XANTENNA__6580__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6506_ _7329_/Q _6423_/X _6503_/X _6505_/X VGND VGND VPWR VPWR _6506_/X sky130_fd_sc_hd__a211o_1
X_3718_ _7030_/Q _4352_/A _4352_/B _3520_/X _7443_/Q VGND VGND VPWR VPWR _3718_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout400_A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7486_ _7525_/CLK hold96/X fanout746/X VGND VGND VPWR VPWR _7486_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4698__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4698_ _4772_/A _4797_/B _4814_/C VGND VGND VPWR VPWR _4698_/Y sky130_fd_sc_hd__nand3_4
XFILLER_107_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6437_ _7551_/Q _6408_/A _6434_/X _7463_/Q _6436_/X VGND VGND VPWR VPWR _6437_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5135__B2 _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3649_ _4515_/B _4527_/A _5596_/B VGND VGND VPWR VPWR _3649_/X sky130_fd_sc_hd__and3_2
XFILLER_134_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6368_ _6970_/Q _6384_/A4 _6144_/B _6032_/Y _7024_/Q VGND VGND VPWR VPWR _6368_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3310 _7622_/Q VGND VGND VPWR VPWR _6650_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3321 _6401_/X VGND VGND VPWR VPWR _7614_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3332 _7207_/Q VGND VGND VPWR VPWR _5566_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3343 _7105_/Q VGND VGND VPWR VPWR _4424_/B sky130_fd_sc_hd__clkdlybuf4s50_2
X_5319_ _5319_/A _5531_/B _5491_/C VGND VGND VPWR VPWR _5319_/X sky130_fd_sc_hd__and3_1
Xhold3354 _7598_/Q VGND VGND VPWR VPWR _6060_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6299_ _7056_/Q _6332_/B _6388_/A3 _6097_/X _7182_/Q VGND VGND VPWR VPWR _6299_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3365 hold24/A VGND VGND VPWR VPWR _6828_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5603__A _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2620 hold933/X VGND VGND VPWR VPWR _4494_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3376 _6910_/Q VGND VGND VPWR VPWR _4000_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2631 hold703/X VGND VGND VPWR VPWR _4190_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2642 hold891/X VGND VGND VPWR VPWR _4482_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2653 _4520_/X VGND VGND VPWR VPWR hold720/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6418__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2664 _5660_/X VGND VGND VPWR VPWR hold506/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2675 _5723_/X VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1930 _4379_/X VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2686 _7489_/Q VGND VGND VPWR VPWR hold985/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1941 hold184/X VGND VGND VPWR VPWR _6000_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1952 _7174_/Q VGND VGND VPWR VPWR hold1952/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2697 hold983/X VGND VGND VPWR VPWR _4536_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1963 hold359/X VGND VGND VPWR VPWR _5663_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_17_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1974 hold300/X VGND VGND VPWR VPWR _5664_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4661__A3 _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1985 hold453/X VGND VGND VPWR VPWR _4184_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6399__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1996 hold427/X VGND VGND VPWR VPWR _5698_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input100_A wb_adr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__B2 _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_566 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5992__B hold40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5374__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6600__C _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_9 _3866_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5429__A2 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6626__B2 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4790__C _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__A1 _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B2 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5670_ _5949_/A1 _5670_/A1 _5676_/S VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__mux2_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5365__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4621_ _4947_/C _4954_/A VGND VGND VPWR VPWR _4966_/A sky130_fd_sc_hd__and2_4
XANTENNA__6562__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7340_ _7576_/CLK _7340_/D fanout718/X VGND VGND VPWR VPWR _7340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ _5912_/A1 _4552_/A1 _4556_/S VGND VGND VPWR VPWR _4552_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3915__A2 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 _5967_/X VGND VGND VPWR VPWR _7552_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3503_ _4328_/A _3598_/B _4388_/B VGND VGND VPWR VPWR _3503_/X sky130_fd_sc_hd__and3_4
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7271_ _7330_/CLK _7271_/D _4079_/A VGND VGND VPWR VPWR _7271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold526 _4202_/X VGND VGND VPWR VPWR _6918_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4483_ _4483_/A0 _4555_/A0 _4484_/S VGND VGND VPWR VPWR _4483_/X sky130_fd_sc_hd__mux2_1
Xhold537 hold537/A VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold548 _5988_/X VGND VGND VPWR VPWR _7571_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold559 hold559/A VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6222_ _7428_/Q _6075_/A _6074_/X _6094_/X _7508_/Q VGND VGND VPWR VPWR _6222_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_89_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3434_ _7370_/Q VGND VGND VPWR VPWR _3434_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _7457_/Q _6112_/C _6079_/X _6119_/X _7401_/Q VGND VGND VPWR VPWR _6153_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__A1 _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5104_ _5407_/A1 _5091_/A _4817_/X _5103_/Y VGND VGND VPWR VPWR _5104_/Y sky130_fd_sc_hd__a31oi_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__B2 _7509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1204 hold2860/X VGND VGND VPWR VPWR hold2861/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ _6081_/C _6099_/D _7588_/Q _7589_/Q VGND VGND VPWR VPWR _6084_/X sky130_fd_sc_hd__and4b_4
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1215 hold2871/X VGND VGND VPWR VPWR _7514_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1226 hold2914/X VGND VGND VPWR VPWR hold2915/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 _4397_/X VGND VGND VPWR VPWR _7063_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1248 hold2916/X VGND VGND VPWR VPWR hold2917/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5035_ _5035_/A _5035_/B _5035_/C _5035_/D VGND VGND VPWR VPWR _5035_/Y sky130_fd_sc_hd__nor4_1
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1259 hold2923/X VGND VGND VPWR VPWR hold2924/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4981__B _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3851__B2 _4174_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6986_ _7000_/CLK _6986_/D VGND VGND VPWR VPWR _6986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5937_ hold20/X _5937_/A1 _5937_/S VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__mux2_1
XANTENNA__3603__A1 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3603__B2 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_12_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout615_A _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5868_ hold383/X _5985_/A1 _5871_/S VGND VGND VPWR VPWR _5868_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6148__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7607_ _7621_/CLK _7607_/D fanout705/X VGND VGND VPWR VPWR _7607_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4819_ _4888_/B _4856_/A _5058_/D VGND VGND VPWR VPWR _5011_/B sky130_fd_sc_hd__and3b_4
XANTENNA__5356__A1 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5799_ _5997_/A1 _5799_/A1 _5802_/S VGND VGND VPWR VPWR _5799_/X sky130_fd_sc_hd__mux2_1
X_7538_ _7542_/CLK _7538_/D fanout713/X VGND VGND VPWR VPWR _7538_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3906__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6420__C _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6305__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7469_ _7525_/CLK _7469_/D fanout745/X VGND VGND VPWR VPWR _7469_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold1632_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6320__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3140 _7137_/Q VGND VGND VPWR VPWR hold3140/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR _4563_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3151 hold3151/A VGND VGND VPWR VPWR _5912_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR _5071_/C sky130_fd_sc_hd__buf_6
XFILLER_49_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3162 _7415_/Q VGND VGND VPWR VPWR hold3162/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6608__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR input124/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3173 _4323_/X VGND VGND VPWR VPWR hold3173/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input148_A wb_dat_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR _6811_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3184 hold3184/A VGND VGND VPWR VPWR _4486_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR _6818_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2450 hold879/X VGND VGND VPWR VPWR _5702_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3195 _4341_/X VGND VGND VPWR VPWR hold3195/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR _6809_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2461 _7364_/Q VGND VGND VPWR VPWR hold897/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR _6824_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2472 _7178_/Q VGND VGND VPWR VPWR hold881/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2483 _7168_/Q VGND VGND VPWR VPWR hold885/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2494 _7032_/Q VGND VGND VPWR VPWR hold919/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1760 _5951_/X VGND VGND VPWR VPWR hold275/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1771 hold119/X VGND VGND VPWR VPWR _7339_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4634__A3 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1782 _5847_/X VGND VGND VPWR VPWR hold102/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1793 hold38/X VGND VGND VPWR VPWR _3576_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3842__A1 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4383__S _4387_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5595__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6792__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4131__B _4131_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5243__A _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7425__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4293__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6840_ _6861_/A _6869_/B VGND VGND VPWR VPWR _6840_/X sky130_fd_sc_hd__and2_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6783__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6771_ _7055_/Q _6434_/B _6771_/A3 _6419_/C _7141_/Q VGND VGND VPWR VPWR _6771_/X
+ sky130_fd_sc_hd__a32o_1
X_3983_ _7343_/Q _3545_/X _3980_/X _3981_/X _3982_/X VGND VGND VPWR VPWR _3983_/X
+ sky130_fd_sc_hd__a2111o_1
X_5722_ hold40/X _5722_/B _5731_/B _5893_/B VGND VGND VPWR VPWR _5730_/S sky130_fd_sc_hd__and4_4
XANTENNA__3597__B1 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7395_/CLK sky130_fd_sc_hd__clkbuf_16
X_5653_ _5995_/A1 _5653_/A1 _5658_/S VGND VGND VPWR VPWR _5653_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4604_ _4831_/A _4860_/A _4772_/A _4805_/B VGND VGND VPWR VPWR _4604_/Y sky130_fd_sc_hd__nor4_1
XFILLER_176_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3864__C _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5584_ _5950_/A1 _5584_/A1 _5586_/S VGND VGND VPWR VPWR _5584_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7095_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_163_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7323_ _7539_/CLK _7323_/D fanout708/X VGND VGND VPWR VPWR _7323_/Q sky130_fd_sc_hd__dfrtp_4
Xhold301 hold301/A VGND VGND VPWR VPWR _7283_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ _4553_/A0 _4535_/A1 _4538_/S VGND VGND VPWR VPWR _4535_/X sky130_fd_sc_hd__mux2_1
Xhold312 hold312/A VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5852__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold323 hold323/A VGND VGND VPWR VPWR _7188_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2914_A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7254_ _7263_/CLK _7254_/D fanout689/X VGND VGND VPWR VPWR _7254_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold345 hold345/A VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold356 hold356/A VGND VGND VPWR VPWR _7094_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4466_ _4466_/A0 _5853_/A0 _4466_/S VGND VGND VPWR VPWR _4466_/X sky130_fd_sc_hd__mux2_1
Xhold367 hold367/A VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold378 hold378/A VGND VGND VPWR VPWR _7274_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6205_ _7291_/Q _6144_/A _6270_/C1 _6032_/Y _7347_/Q VGND VGND VPWR VPWR _6205_/X
+ sky130_fd_sc_hd__a32o_1
Xhold389 hold389/A VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3417_ _7506_/Q VGND VGND VPWR VPWR _3417_/Y sky130_fd_sc_hd__inv_2
X_7185_ _7185_/CLK _7185_/D fanout725/X VGND VGND VPWR VPWR _7185_/Q sky130_fd_sc_hd__dfrtp_4
X_4397_ _5815_/A1 _4397_/A1 _4399_/S VGND VGND VPWR VPWR _4397_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout398_A _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _7296_/Q _6136_/B _6136_/C VGND VGND VPWR VPWR _6136_/X sky130_fd_sc_hd__and3_1
XFILLER_86_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1001 hold2990/X VGND VGND VPWR VPWR hold2991/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1012 _4432_/X VGND VGND VPWR VPWR _7085_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 _4441_/X VGND VGND VPWR VPWR _7093_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1034 hold2836/X VGND VGND VPWR VPWR hold2837/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6067_ _6067_/A _6067_/B VGND VGND VPWR VPWR _6067_/X sky130_fd_sc_hd__and2_4
XANTENNA__4992__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout565_A _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1045 hold3100/X VGND VGND VPWR VPWR hold3101/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1056 hold2886/X VGND VGND VPWR VPWR hold2887/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1067 hold1067/A VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
X_5018_ _5034_/C _5018_/B VGND VGND VPWR VPWR _5021_/B sky130_fd_sc_hd__nand2_1
Xhold1078 hold3012/X VGND VGND VPWR VPWR hold1078/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 hold1089/A VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6369__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _7176_/CLK _6969_/D fanout722/X VGND VGND VPWR VPWR _6969_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6526__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5762__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold890 hold890/A VGND VGND VPWR VPWR _7049_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold3130_A _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5213__D _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2280 hold801/X VGND VGND VPWR VPWR _5665_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4068__B2 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2291 hold607/X VGND VGND VPWR VPWR _5658_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3815__A1 _6913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1590 hold83/X VGND VGND VPWR VPWR _5981_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6765__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5937__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3579__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4240__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6517__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3594__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4142__A _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4320_ _3607_/Y _4320_/A1 _4321_/S VGND VGND VPWR VPWR _6999_/D sky130_fd_sc_hd__mux2_1
XFILLER_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4796__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6296__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4288__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4251_ _4251_/A0 _5993_/A1 _4258_/S VGND VGND VPWR VPWR _4251_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2230_A _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4182_ _4182_/A0 _5876_/A1 _4190_/S VGND VGND VPWR VPWR _4182_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6048__A2 _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7432__SET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3806__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3806__B2 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4317__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3859__C _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6823_ _4114_/B _7105_/D _6823_/A3 _4428_/Y _4430_/B VGND VGND VPWR VPWR _7645_/D
+ sky130_fd_sc_hd__o41ai_2
XANTENNA__6756__B1 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6220__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6754_ _7176_/Q _6747_/B _6747_/C _6443_/X _7196_/Q VGND VGND VPWR VPWR _6754_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3966_ _6911_/Q _5612_/B _5947_/A _5713_/A _7327_/Q VGND VGND VPWR VPWR _3966_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4231__A1 _4422_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5705_ _5894_/A0 _5705_/A1 _5712_/S VGND VGND VPWR VPWR _5705_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3585__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6685_ _7042_/Q _6408_/B _6462_/X _7032_/Q _6684_/X VGND VGND VPWR VPWR _6685_/X
+ sky130_fd_sc_hd__a221o_1
X_3897_ _7002_/Q _4322_/A _3889_/X _3892_/X _3896_/X VGND VGND VPWR VPWR _3897_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3990__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5636_ _5979_/A0 _5636_/A1 _5639_/S VGND VGND VPWR VPWR _5636_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5567_ _4778_/A _5410_/X _5308_/C _5148_/C _5308_/A VGND VGND VPWR VPWR _5568_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_105_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7306_ _7306_/CLK _7306_/D _4079_/A VGND VGND VPWR VPWR _7306_/Q sky130_fd_sc_hd__dfrtp_4
Xhold120 _6922_/Q VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3742__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4518_ _4518_/A0 _5788_/A1 _4520_/S VGND VGND VPWR VPWR _4518_/X sky130_fd_sc_hd__mux2_1
Xhold131 hold131/A VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold142 _6916_/Q VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold153 hold153/A VGND VGND VPWR VPWR _6914_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5498_ _5053_/C _4876_/Y _5328_/X _5497_/X VGND VGND VPWR VPWR _5499_/B sky130_fd_sc_hd__a31o_1
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold175 hold175/A VGND VGND VPWR VPWR _7251_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7237_ _7238_/CLK _7237_/D fanout690/X VGND VGND VPWR VPWR _7237_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6287__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold186 hold186/A VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout682_A _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4449_ _4473_/A _4455_/A _4455_/C _4533_/B VGND VGND VPWR VPWR _4454_/S sky130_fd_sc_hd__and4_4
Xhold197 hold197/A VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__buf_12
Xfanout600 hold1449/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__buf_6
Xfanout611 _7596_/Q VGND VGND VPWR VPWR _6441_/D sky130_fd_sc_hd__clkbuf_8
Xfanout622 _7591_/Q VGND VGND VPWR VPWR _6099_/D sky130_fd_sc_hd__buf_6
XFILLER_120_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1428_A hold1428/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout633 hold3326/X VGND VGND VPWR VPWR _4058_/B sky130_fd_sc_hd__buf_4
Xfanout644 _4887_/X VGND VGND VPWR VPWR _5049_/C sky130_fd_sc_hd__clkbuf_16
X_7168_ _7181_/CLK _7168_/D fanout721/X VGND VGND VPWR VPWR _7168_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6119_/A _6119_/B _6121_/A _6119_/D VGND VGND VPWR VPWR _6119_/X sky130_fd_sc_hd__and4_4
XFILLER_86_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout677 _4581_/X VGND VGND VPWR VPWR _5038_/A sky130_fd_sc_hd__buf_8
Xfanout688 fanout691/X VGND VGND VPWR VPWR fanout688/X sky130_fd_sc_hd__buf_8
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ _7197_/CLK hold11/X fanout742/X VGND VGND VPWR VPWR _7099_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout699 fanout702/X VGND VGND VPWR VPWR fanout699/X sky130_fd_sc_hd__clkbuf_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5970__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3981__B1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input76_A qspi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3345_A _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5789__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6450__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6738__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6202__A2 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3820_ _6876_/Q _3931_/B _5632_/B _3564_/X _7361_/Q VGND VGND VPWR VPWR _3828_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4213__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3751_ _6877_/Q _4551_/B _4352_/B _4497_/A _7155_/Q VGND VGND VPWR VPWR _3751_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5961__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6470_ _7503_/Q _6466_/X _6467_/X _7415_/Q _6469_/X VGND VGND VPWR VPWR _6471_/D
+ sky130_fd_sc_hd__a221o_1
X_3682_ _3682_/A _4491_/C _5640_/C VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__and3_2
XFILLER_173_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5421_ _4595_/Y _5495_/C1 _4956_/A _4834_/Y _5494_/B2 VGND VGND VPWR VPWR _5422_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6498__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput203 wire378/X VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XANTENNA__3724__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput214 _4149_/X VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ _4907_/B _4940_/D _5346_/X _5217_/X _5065_/A VGND VGND VPWR VPWR _5352_/Y
+ sky130_fd_sc_hd__a32oi_4
Xoutput225 _7662_/X VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
XFILLER_99_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput236 _7670_/X VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput247 _4125_/X VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
X_4303_ _4346_/C _5623_/B _5619_/C VGND VGND VPWR VPWR _4303_/X sky130_fd_sc_hd__and3_1
Xoutput258 _7243_/Q VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
Xoutput269 _6919_/Q VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
X_5283_ _5059_/B _5115_/X _5282_/X VGND VGND VPWR VPWR _5481_/A sky130_fd_sc_hd__a21oi_1
X_7022_ _7497_/CLK _7022_/D fanout707/X VGND VGND VPWR VPWR _7022_/Q sky130_fd_sc_hd__dfrtp_4
X_4234_ _5651_/A1 _5894_/A0 _4248_/S VGND VGND VPWR VPWR _4234_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4165_ _6938_/Q input93/X _7262_/Q VGND VGND VPWR VPWR _4165_/X sky130_fd_sc_hd__mux2_2
XFILLER_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4096_ input123/X input122/X _4096_/C _4096_/D VGND VGND VPWR VPWR _4096_/X sky130_fd_sc_hd__and4bb_2
XFILLER_71_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4452__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6729__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6806_ _4427_/B _6806_/A2 _6806_/B1 _4426_/Y _6805_/X VGND VGND VPWR VPWR _6806_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4204__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ _5024_/A1 _4669_/X _5038_/A _4974_/B VGND VGND VPWR VPWR _5018_/B sky130_fd_sc_hd__o211a_2
XANTENNA__5952__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3949_ _7016_/Q _4346_/C _5619_/B _3948_/X VGND VGND VPWR VPWR _3949_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3465__A_N _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6737_ _6991_/Q _6420_/B _6462_/X _7034_/Q VGND VGND VPWR VPWR _6737_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6668_ _7056_/Q _6466_/D _6651_/C _6452_/X _7021_/Q VGND VGND VPWR VPWR _6668_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5619_ _5619_/A _5619_/B _5619_/C VGND VGND VPWR VPWR _5620_/S sky130_fd_sc_hd__and3_1
X_6599_ _6599_/A1 _4116_/X _6067_/X _6598_/X VGND VGND VPWR VPWR _7620_/D sky130_fd_sc_hd__o31a_1
XFILLER_191_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3715__B1 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1545_A _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout441 _5612_/C VGND VGND VPWR VPWR _5596_/A sky130_fd_sc_hd__buf_8
Xfanout452 hold40/X VGND VGND VPWR VPWR _5640_/A sky130_fd_sc_hd__buf_6
Xfanout463 _6073_/X VGND VGND VPWR VPWR _6274_/A3 sky130_fd_sc_hd__buf_6
XFILLER_93_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6680__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout474 _6429_/X VGND VGND VPWR VPWR _6651_/C sky130_fd_sc_hd__buf_8
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout485 _6093_/X VGND VGND VPWR VPWR _6276_/A3 sky130_fd_sc_hd__buf_6
XANTENNA__4883__C _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout496 _6042_/X VGND VGND VPWR VPWR _6434_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA_input130_A wb_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6904__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6432__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4443__A1 _5635_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__A1 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__B2 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5943__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6499__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3706__B1 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6671__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3470__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2026_A _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5970_ _5970_/A0 _5997_/A1 _5973_/S VGND VGND VPWR VPWR _5970_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4434__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4921_ _5213_/A _4997_/B _4933_/A _5260_/D VGND VGND VPWR VPWR _4922_/B sky130_fd_sc_hd__and4_1
XFILLER_80_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7640_ _7641_/CLK _7640_/D fanout753/X VGND VGND VPWR VPWR _7640_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6082__A _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6187__A1 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4852_ _5494_/B2 _4595_/Y _4695_/Y _4427_/C VGND VGND VPWR VPWR _5294_/A sky130_fd_sc_hd__o31a_2
XANTENNA__6187__B2 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3803_ _7353_/Q _5803_/A hold90/A _5758_/A _7369_/Q VGND VGND VPWR VPWR _3803_/X
+ sky130_fd_sc_hd__a32o_1
X_7571_ _7573_/CLK _7571_/D fanout733/X VGND VGND VPWR VPWR _7571_/Q sky130_fd_sc_hd__dfrtp_4
X_4783_ _4772_/A _4801_/B _5404_/A _5410_/B VGND VGND VPWR VPWR _4783_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6522_ _6521_/X _6522_/A1 _6751_/S VGND VGND VPWR VPWR _6522_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3734_ _3923_/S _3734_/B VGND VGND VPWR VPWR _3734_/Y sky130_fd_sc_hd__nand2_2
XFILLER_174_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6453_ _7479_/Q _6447_/C _6459_/C _6452_/X _7343_/Q VGND VGND VPWR VPWR _6453_/X
+ sky130_fd_sc_hd__a32o_1
X_3665_ _4473_/A _4551_/A _4551_/C VGND VGND VPWR VPWR _3665_/X sky130_fd_sc_hd__and3_2
X_5404_ _5404_/A _5404_/B _5404_/C _5404_/D VGND VGND VPWR VPWR _5405_/C sky130_fd_sc_hd__nand4_1
X_6384_ _7191_/Q _6099_/D _7590_/Q _6384_/A4 _6082_/C VGND VGND VPWR VPWR _6384_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_133_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3596_ _7293_/Q _5668_/A _3592_/X _3593_/X _3595_/X VGND VGND VPWR VPWR _3606_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_127_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5335_ _5034_/B _5030_/C _5339_/B _5334_/X VGND VGND VPWR VPWR _5335_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5860__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2802 hold959/X VGND VGND VPWR VPWR _4531_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5266_ _5266_/A _5266_/B _5256_/X VGND VGND VPWR VPWR _5266_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2813 _7143_/Q VGND VGND VPWR VPWR hold939/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2824 _7655_/A VGND VGND VPWR VPWR hold997/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7005_ _7210_/CLK _7005_/D fanout702/X VGND VGND VPWR VPWR _7005_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2835 _5759_/X VGND VGND VPWR VPWR _7367_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5465__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2846 hold2846/A VGND VGND VPWR VPWR _4262_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6662__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4217_ _4251_/A0 _5993_/A1 _4231_/S VGND VGND VPWR VPWR _4217_/X sky130_fd_sc_hd__mux2_1
Xhold2857 _4245_/X VGND VGND VPWR VPWR hold2857/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5197_ _4858_/Y _5528_/A3 _4873_/X _4672_/X _5046_/A VGND VGND VPWR VPWR _5423_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold2868 _5671_/X VGND VGND VPWR VPWR hold2868/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout478_A _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2879 _7530_/Q VGND VGND VPWR VPWR hold2879/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4148_ _7268_/Q input81/X _4174_/B VGND VGND VPWR VPWR _4148_/X sky130_fd_sc_hd__mux2_8
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4079_ _4079_/A _6839_/B VGND VGND VPWR VPWR _4079_/X sky130_fd_sc_hd__and2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4976__A2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1495_A _4422_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5689__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3951__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4878__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6350__A1 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6350__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5055__B _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5770__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6653__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4386__S _4387_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input39_A mgmt_gpio_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5208__A3 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4416__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6708__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5916__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7399__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire650 _4856_/Y VGND VGND VPWR VPWR _5199_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_171_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold708 _5683_/X VGND VGND VPWR VPWR _7300_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold719 hold719/A VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3450_ _4007_/B _3450_/B VGND VGND VPWR VPWR _3450_/X sky130_fd_sc_hd__and2b_1
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_672 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5120_ _4845_/X _5180_/B _5119_/X VGND VGND VPWR VPWR _5122_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2109 _6939_/Q VGND VGND VPWR VPWR hold489/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _5051_/A _5051_/B _5051_/C VGND VGND VPWR VPWR _5052_/C sky130_fd_sc_hd__nand3_1
XANTENNA__6644__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1408 _6884_/Q VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1419 hold1/X VGND VGND VPWR VPWR _4189_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4655__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4002_ _6910_/Q _6909_/Q _4006_/A VGND VGND VPWR VPWR _4003_/B sky130_fd_sc_hd__and3_1
XFILLER_93_751 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4407__A1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7220__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5953_ _5953_/A0 _5953_/A1 _5955_/S VGND VGND VPWR VPWR _5953_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5080__B2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4904_ _4904_/A _4904_/B VGND VGND VPWR VPWR _4906_/A sky130_fd_sc_hd__nor2_1
X_5884_ _5938_/C _5956_/B _5992_/D VGND VGND VPWR VPWR hold91/A sky130_fd_sc_hd__and3_1
XANTENNA__3630__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7623_ _7625_/CLK _7623_/D fanout706/X VGND VGND VPWR VPWR _7623_/Q sky130_fd_sc_hd__dfrtp_1
X_4835_ _5494_/B2 _4595_/Y _4832_/Y _4834_/Y _4956_/A VGND VGND VPWR VPWR _4837_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5855__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4766_ _4766_/A _4766_/B VGND VGND VPWR VPWR _4766_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6580__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7554_ _7575_/CLK _7554_/D fanout734/X VGND VGND VPWR VPWR _7554_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6505_ _7297_/Q _6420_/A _6421_/X _7321_/Q _6504_/X VGND VGND VPWR VPWR _6505_/X
+ sky130_fd_sc_hd__a221o_1
X_3717_ _7459_/Q _5857_/A _3713_/X _3714_/X _3716_/X VGND VGND VPWR VPWR _3717_/X
+ sky130_fd_sc_hd__a2111o_1
X_7485_ _7565_/CLK hold92/X fanout746/X VGND VGND VPWR VPWR _7485_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4697_ _4909_/D _4797_/B _4814_/C VGND VGND VPWR VPWR _5091_/C sky130_fd_sc_hd__and3_4
XFILLER_119_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4698__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3648_ _4364_/A _4388_/B _5596_/B VGND VGND VPWR VPWR _3648_/X sky130_fd_sc_hd__and3_2
X_6436_ _7319_/Q _6421_/X _6435_/X _7511_/Q VGND VGND VPWR VPWR _6436_/X sky130_fd_sc_hd__a22o_1
XFILLER_161_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6367_ _7115_/Q _6317_/C _6332_/C _7034_/Q _6366_/X VGND VGND VPWR VPWR _6367_/X
+ sky130_fd_sc_hd__a221o_1
X_3579_ _5659_/B _5623_/B _3578_/X _4248_/S input69/X VGND VGND VPWR VPWR _3579_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3300 _7621_/Q VGND VGND VPWR VPWR _6649_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3311 _7619_/Q VGND VGND VPWR VPWR _6598_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout595_A hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3322 _7603_/Q VGND VGND VPWR VPWR _6169_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5318_ _5494_/B2 _4821_/Y _4802_/Y _4595_/Y VGND VGND VPWR VPWR _5531_/B sky130_fd_sc_hd__a211o_1
Xhold3333 _7601_/Q VGND VGND VPWR VPWR _6066_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3344 _7597_/Q VGND VGND VPWR VPWR _6055_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6298_ _7172_/Q _6110_/X _6112_/X _6874_/Q _6297_/X VGND VGND VPWR VPWR _6303_/B
+ sky130_fd_sc_hd__a221o_1
Xhold2610 _5783_/X VGND VGND VPWR VPWR hold900/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3355 _7628_/Q VGND VGND VPWR VPWR _6779_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3366 _6829_/X VGND VGND VPWR VPWR _7646_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2621 _7276_/Q VGND VGND VPWR VPWR hold989/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5603__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6635__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__buf_8
Xhold2632 _4190_/X VGND VGND VPWR VPWR hold704/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3377 _7587_/Q VGND VGND VPWR VPWR _4100_/A3 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5249_ _4659_/Y _5516_/A3 _5247_/X VGND VGND VPWR VPWR _5249_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout762_A _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2643 _7022_/Q VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2654 _7151_/Q VGND VGND VPWR VPWR hold791/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2665 _7443_/Q VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1920 _7039_/Q VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6418__C _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2676 hold520/X VGND VGND VPWR VPWR _7335_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1931 _7558_/Q VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1942 _6000_/X VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2687 hold985/X VGND VGND VPWR VPWR _5896_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2698 _7429_/Q VGND VGND VPWR VPWR hold943/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1953 hold1953/A VGND VGND VPWR VPWR _4524_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1964 _5663_/X VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1975 _5664_/X VGND VGND VPWR VPWR hold301/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1986 _4184_/X VGND VGND VPWR VPWR hold454/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6399__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1997 _5698_/X VGND VGND VPWR VPWR hold428/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6434__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3621__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6020__A0 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5765__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3909__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6571__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4689__B1_N _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3688__A2 _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6626__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5429__A3 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4129__B _4129_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4627__B1_N _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3612__A2 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4616_/Y _4617_/Y _4618_/Y _4615_/Y VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__a22oi_4
XANTENNA__6562__A1 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4551_ _4551_/A _4551_/B _4551_/C _4551_/D VGND VGND VPWR VPWR _4556_/S sky130_fd_sc_hd__nand4_4
XANTENNA__3915__A3 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3502_ _3576_/C _3576_/B VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__and2_4
X_7270_ _7522_/CLK _7270_/D fanout744/X VGND VGND VPWR VPWR _7270_/Q sky130_fd_sc_hd__dfrtp_1
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4482_ _4482_/A0 _5914_/A1 _4484_/S VGND VGND VPWR VPWR _4482_/X sky130_fd_sc_hd__mux2_1
Xhold516 _5760_/X VGND VGND VPWR VPWR _7368_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold527 hold527/A VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold538 hold538/A VGND VGND VPWR VPWR _6992_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6221_ _7324_/Q _6119_/D _6081_/X _6090_/X _7380_/Q VGND VGND VPWR VPWR _6221_/X
+ sky130_fd_sc_hd__a32o_1
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold47_A hold47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3433_ _7378_/Q VGND VGND VPWR VPWR _3433_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3679__A2 _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5704__A _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _7481_/Q _6112_/X _6151_/X _6150_/X _6149_/X VGND VGND VPWR VPWR _6152_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5561_/A1 _4806_/Y _5509_/A3 _5102_/Y _5101_/Y VGND VGND VPWR VPWR _5103_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6617__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _7455_/Q _6075_/A _6079_/X _6082_/X _7319_/Q VGND VGND VPWR VPWR _6083_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1205 hold2862/X VGND VGND VPWR VPWR _7506_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1216 hold2891/X VGND VGND VPWR VPWR hold2892/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1227 _5933_/X VGND VGND VPWR VPWR _7522_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5038_/A _5034_/B _5034_/C VGND VGND VPWR VPWR _5035_/C sky130_fd_sc_hd__and3_1
Xhold1238 hold2953/X VGND VGND VPWR VPWR hold2954/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1249 hold2918/X VGND VGND VPWR VPWR _7008_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2894_A _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6985_ _7000_/CLK _6985_/D VGND VGND VPWR VPWR _6985_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6250__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5936_ _5990_/A1 _5936_/A1 _5937_/S VGND VGND VPWR VPWR _5936_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ _5867_/A0 _5975_/A0 _5871_/S VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7606_ _7621_/CLK _7606_/D fanout708/X VGND VGND VPWR VPWR _7606_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout510_A _4857_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4818_ _4818_/A _4818_/B _4818_/C VGND VGND VPWR VPWR _4824_/A sky130_fd_sc_hd__nor3_1
XANTENNA_fanout608_A _3444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5798_ _5969_/A1 _5798_/A1 _5802_/S VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__mux2_1
X_7537_ _7537_/CLK _7537_/D fanout707/X VGND VGND VPWR VPWR _7537_/Q sky130_fd_sc_hd__dfrtp_4
X_4749_ _4814_/C _4899_/A2 _4657_/C VGND VGND VPWR VPWR _4884_/B sky130_fd_sc_hd__a21oi_2
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5108__A2 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7468_ _7565_/CLK _7468_/D fanout748/X VGND VGND VPWR VPWR _7468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6419_ _6419_/A _6419_/B _6419_/C _6419_/D VGND VGND VPWR VPWR _6419_/Y sky130_fd_sc_hd__nor4_1
X_7399_ _7399_/CLK _7399_/D fanout719/X VGND VGND VPWR VPWR _7399_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5614__A _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3130 _7439_/Q VGND VGND VPWR VPWR hold3130/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3141 hold3141/A VGND VGND VPWR VPWR _4480_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR _4563_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3152 _7265_/Q VGND VGND VPWR VPWR hold3152/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6608__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR _5071_/B sky130_fd_sc_hd__buf_6
Xhold3163 hold3163/A VGND VGND VPWR VPWR _5813_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR input125/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3174 _7209_/Q VGND VGND VPWR VPWR hold3174/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR _6815_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4619__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3185 _7248_/Q VGND VGND VPWR VPWR hold3185/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2440 _7259_/Q VGND VGND VPWR VPWR hold581/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2451 _5702_/X VGND VGND VPWR VPWR hold880/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR _6821_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3196 _7061_/Q VGND VGND VPWR VPWR hold3196/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR _6812_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2462 hold897/X VGND VGND VPWR VPWR _5755_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput169 wb_stb_i VGND VGND VPWR VPWR _4093_/B sky130_fd_sc_hd__buf_4
Xhold2473 hold881/X VGND VGND VPWR VPWR _4529_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2484 hold885/X VGND VGND VPWR VPWR _4517_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2495 hold919/X VGND VGND VPWR VPWR _4360_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1750 hold150/X VGND VGND VPWR VPWR _5789_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1761 _7091_/Q VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1772 _7432_/Q VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1783 hold102/X VGND VGND VPWR VPWR _7446_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4891__C _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1794 _4203_/X VGND VGND VPWR VPWR _4207_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3842__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6241__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk _7416_/CLK VGND VGND VPWR VPWR _7266_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6529__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3375_A _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output262_A _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6058__C _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5283__A1 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6480__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3833__A2 _3492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6074__B _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3982_ _7244_/Q _3590_/C _5614_/B _5893_/A _7487_/Q VGND VGND VPWR VPWR _3982_/X
+ sky130_fd_sc_hd__a32o_1
X_6770_ _7126_/Q _6420_/C _6455_/X _7201_/Q _6769_/X VGND VGND VPWR VPWR _6773_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3597__A1 _7509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5721_ _5955_/A1 _5721_/A1 _5721_/S VGND VGND VPWR VPWR _5721_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3597__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _5949_/A1 _5652_/A1 _5658_/S VGND VGND VPWR VPWR _5652_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6535__A1 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4603__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4603_ _4831_/A _4860_/A VGND VGND VPWR VPWR _5260_/B sky130_fd_sc_hd__nor2_8
X_5583_ hold198/X _5583_/A1 _5586_/S VGND VGND VPWR VPWR _5583_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7322_ _7581_/CLK _7322_/D fanout716/X VGND VGND VPWR VPWR _7322_/Q sky130_fd_sc_hd__dfrtp_4
X_4534_ _5876_/A1 _4534_/A1 _4538_/S VGND VGND VPWR VPWR _4534_/X sky130_fd_sc_hd__mux2_1
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold313 hold313/A VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6299__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold324 hold324/A VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4465_ _4465_/A0 _5585_/A0 _4466_/S VGND VGND VPWR VPWR _4465_/X sky130_fd_sc_hd__mux2_1
X_7253_ _7263_/CLK _7253_/D fanout689/X VGND VGND VPWR VPWR _7253_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold346 hold346/A VGND VGND VPWR VPWR _6969_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold357 hold357/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold368 hold368/A VGND VGND VPWR VPWR _7346_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3416_ _7514_/Q VGND VGND VPWR VPWR _3416_/Y sky130_fd_sc_hd__inv_2
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6204_ _7363_/Q _6332_/C _6379_/B1 _7395_/Q _6203_/X VGND VGND VPWR VPWR _6204_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7184_ _7184_/CLK _7184_/D fanout725/X VGND VGND VPWR VPWR _7184_/Q sky130_fd_sc_hd__dfstp_4
X_4396_ hold198/X _4396_/A1 _4399_/S VGND VGND VPWR VPWR _4396_/X sky130_fd_sc_hd__mux2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _7344_/Q _6032_/Y _6274_/A3 _7384_/Q _6134_/X VGND VGND VPWR VPWR _6135_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 hold2992/X VGND VGND VPWR VPWR _6949_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1013 _4078_/A VGND VGND VPWR VPWR _5650_/A1 sky130_fd_sc_hd__buf_6
X_6066_ _4099_/D _7584_/Q _6065_/Y _6062_/X _6066_/B2 VGND VGND VPWR VPWR _6066_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1024 hold3055/X VGND VGND VPWR VPWR hold3056/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1035 hold3060/X VGND VGND VPWR VPWR hold3061/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__C1 _3806_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1046 _5867_/X VGND VGND VPWR VPWR _7463_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1057 hold2888/X VGND VGND VPWR VPWR _7080_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5006_/Y _5008_/X _5016_/Y VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__a21oi_1
Xhold1068 hold3000/X VGND VGND VPWR VPWR hold1068/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1079 hold1079/A VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
XANTENNA_fanout558_A _5673_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3824__A2 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6968_ _7176_/CLK _6968_/D fanout722/X VGND VGND VPWR VPWR _6968_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5919_ _5919_/A0 _5991_/A1 _5919_/S VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__mux2_1
X_6899_ _7075_/CLK _6899_/D _6849_/X VGND VGND VPWR VPWR _6899_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5329__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6526__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6526__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5328__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1742_A _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3760__A1 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3760__B2 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input160_A wb_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold880 hold880/A VGND VGND VPWR VPWR _7317_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold891 hold891/A VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2270 _5960_/X VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input21_A mask_rev_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2281 _5665_/X VGND VGND VPWR VPWR hold802/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2292 _5658_/X VGND VGND VPWR VPWR hold608/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1580 _5908_/X VGND VGND VPWR VPWR hold223/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1591 _5981_/X VGND VGND VPWR VPWR hold84/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_189_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6765__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3579__A1 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4142__B _4142_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7528__SET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4250_ _4250_/A1 hold365/X _4168_/D _4231_/S _5956_/C VGND VGND VPWR VPWR _4258_/S
+ sky130_fd_sc_hd__o311a_4
X_4181_ _4076_/B _4181_/A1 _4181_/S VGND VGND VPWR VPWR _4181_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5404__D _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5256__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3806__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6205__B1 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6822_ _6821_/X _6822_/A1 _6822_/S VGND VGND VPWR VPWR _7644_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6753_ _7131_/Q _6424_/X _6427_/X _7121_/Q VGND VGND VPWR VPWR _6753_/X sky130_fd_sc_hd__a22o_1
X_3965_ _7455_/Q _4431_/A _5866_/B _3964_/X VGND VGND VPWR VPWR _3965_/X sky130_fd_sc_hd__a31o_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5704_ _5704_/A _5947_/C VGND VGND VPWR VPWR _5712_/S sky130_fd_sc_hd__nand2_8
XANTENNA__6508__A1 _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3896_ _7424_/Q _3537_/X _3862_/X _3893_/X _3895_/X VGND VGND VPWR VPWR _3896_/X
+ sky130_fd_sc_hd__a2111o_1
X_6684_ _7027_/Q _6459_/B _6459_/C _6460_/X _7113_/Q VGND VGND VPWR VPWR _6684_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3990__B2 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5635_ _5635_/A0 _5635_/A1 _5639_/S VGND VGND VPWR VPWR _5635_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5863__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5566_ _5566_/A1 _5580_/A2 _5565_/X _5557_/X VGND VGND VPWR VPWR _7207_/D sky130_fd_sc_hd__a211o_1
XFILLER_3_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold110 hold110/A VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7305_ _7329_/CLK _7305_/D fanout704/X VGND VGND VPWR VPWR _7305_/Q sky130_fd_sc_hd__dfrtp_4
Xhold121 hold121/A VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3742__A1 _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold132 hold132/A VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4517_ _4517_/A0 _4547_/A0 _4520_/S VGND VGND VPWR VPWR _4517_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5497_ _5183_/B _4876_/Y _5425_/X _5172_/X VGND VGND VPWR VPWR _5497_/X sky130_fd_sc_hd__a31o_1
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold154 hold154/A VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold165 hold165/A VGND VGND VPWR VPWR _7422_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7236_ _7238_/CLK _7236_/D fanout690/X VGND VGND VPWR VPWR _7236_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6287__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4448_ _4448_/A0 _5991_/A1 _4448_/S VGND VGND VPWR VPWR _4448_/X sky130_fd_sc_hd__mux2_1
Xfanout601 _4101_/X VGND VGND VPWR VPWR _6463_/A sky130_fd_sc_hd__buf_8
Xhold187 hold187/A VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout612 _7596_/Q VGND VGND VPWR VPWR _6466_/A sky130_fd_sc_hd__buf_6
Xhold198 hold198/A VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__buf_8
XANTENNA__5495__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6692__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout623 _7591_/Q VGND VGND VPWR VPWR _6119_/A sky130_fd_sc_hd__buf_6
Xfanout634 _7071_/Q VGND VGND VPWR VPWR _4058_/A sky130_fd_sc_hd__buf_8
X_7167_ _7213_/CLK _7167_/D fanout700/X VGND VGND VPWR VPWR _7167_/Q sky130_fd_sc_hd__dfrtp_2
X_4379_ _4379_/A0 _5788_/A1 _4381_/S VGND VGND VPWR VPWR _4379_/X sky130_fd_sc_hd__mux2_1
Xfanout645 _4887_/X VGND VGND VPWR VPWR _5260_/D sky130_fd_sc_hd__buf_6
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6110_/A _6115_/X _6117_/X _6114_/X _6108_/X VGND VGND VPWR VPWR _6118_/Y
+ sky130_fd_sc_hd__a2111oi_1
X_7098_ _7197_/CLK hold17/X fanout742/X VGND VGND VPWR VPWR _7098_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout678 _4581_/X VGND VGND VPWR VPWR _4823_/D sky130_fd_sc_hd__buf_6
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 fanout691/X VGND VGND VPWR VPWR fanout689/X sky130_fd_sc_hd__clkbuf_8
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6444__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6047_/Y _6048_/X _6019_/A _6019_/Y _6433_/D VGND VGND VPWR VPWR _7595_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_86_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3412__A _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6426__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3981__B2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5773__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input69_A mgmt_gpio_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__A _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3338_A _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6278__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7561_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5238__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_35_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7267_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3750_ _7378_/Q _3498_/X _3745_/X _3747_/X _3749_/X VGND VGND VPWR VPWR _3750_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_13_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6071__C _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3681_ _7065_/Q _4394_/A _3676_/X _3677_/X _3680_/X VGND VGND VPWR VPWR _3681_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5174__B1 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5420_ _4595_/Y _4956_/A _4730_/Y _5529_/A _5419_/X VGND VGND VPWR VPWR _5422_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3724__A1 _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput204 _4143_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
X_5351_ _4601_/Y _4956_/B _4726_/Y _4622_/Y VGND VGND VPWR VPWR _5355_/B sky130_fd_sc_hd__a211o_1
XANTENNA__3724__B2 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput215 _7654_/X VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_154_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput226 _7663_/X VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
Xoutput237 _4148_/X VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput248 _4126_/Y VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_4302_ _3570_/Y _4302_/A1 _4302_/S VGND VGND VPWR VPWR _6987_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6123__C1 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput259 _7223_/Q VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
XANTENNA__6269__A3 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5282_ _5282_/A _5282_/B _5282_/C _5282_/D VGND VGND VPWR VPWR _5282_/X sky130_fd_sc_hd__and4_1
XANTENNA__5477__A1 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7021_ _7497_/CLK _7021_/D fanout707/X VGND VGND VPWR VPWR _7021_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6674__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4233_ _6839_/B _3541_/Y _4248_/S _4215_/X _5956_/C VGND VGND VPWR VPWR _4249_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ _7091_/Q _4164_/A1 _7259_/Q VGND VGND VPWR VPWR _4164_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5229__A1 _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4095_ _5115_/A _4095_/B _4095_/C _4095_/D VGND VGND VPWR VPWR _4096_/D sky130_fd_sc_hd__and4_1
XANTENNA__4328__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5858__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6729__B2 _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6805_ _4427_/D _6805_/A2 _6805_/B1 _4427_/C VGND VGND VPWR VPWR _6805_/X sky130_fd_sc_hd__a22o_1
X_4997_ _4997_/A _4997_/B _5404_/C _5410_/B VGND VGND VPWR VPWR _5028_/C sky130_fd_sc_hd__nand4_4
X_6736_ _7044_/Q _6408_/B _6460_/X _7115_/Q _6735_/X VGND VGND VPWR VPWR _6736_/X
+ sky130_fd_sc_hd__a221o_1
X_3948_ _5619_/A _5623_/B _3864_/X _7222_/Q _3947_/X VGND VGND VPWR VPWR _3948_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3963__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6667_ _7197_/Q _6463_/A _6574_/C _6463_/X _7162_/Q VGND VGND VPWR VPWR _6667_/X
+ sky130_fd_sc_hd__a32o_1
X_3879_ _3879_/A _3879_/B _3879_/C _3879_/D VGND VGND VPWR VPWR _3922_/A sky130_fd_sc_hd__nor4_2
XFILLER_191_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5618_ hold288/X _5951_/A1 _5618_/S VGND VGND VPWR VPWR _5618_/X sky130_fd_sc_hd__mux2_1
X_6598_ _6649_/S _6598_/A2 _6573_/S _6597_/X VGND VGND VPWR VPWR _6598_/X sky130_fd_sc_hd__a211o_1
XFILLER_152_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5549_ _5203_/A _5089_/D _5549_/A3 _5343_/A _5343_/B VGND VGND VPWR VPWR _5550_/D
+ sky130_fd_sc_hd__a311oi_4
XFILLER_151_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1538_A _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5468__A1 _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5468__B2 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6665__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7219_ _4150_/A1 _7219_/D _6871_/X VGND VGND VPWR VPWR _7219_/Q sky130_fd_sc_hd__dfrtn_1
Xfanout420 _5213_/C VGND VGND VPWR VPWR _4907_/B sky130_fd_sc_hd__buf_8
XANTENNA__3479__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout431 _5063_/D VGND VGND VPWR VPWR _5339_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA_hold1705_A _7496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout442 _3489_/Y VGND VGND VPWR VPWR _5612_/C sky130_fd_sc_hd__buf_8
Xfanout453 hold40/X VGND VGND VPWR VPWR _5938_/A sky130_fd_sc_hd__buf_6
Xfanout464 _4876_/Y VGND VGND VPWR VPWR _5216_/A sky130_fd_sc_hd__buf_6
Xfanout475 _6429_/X VGND VGND VPWR VPWR _6769_/A3 sky130_fd_sc_hd__buf_8
Xfanout486 _6084_/X VGND VGND VPWR VPWR _6388_/A3 sky130_fd_sc_hd__clkbuf_16
XFILLER_171_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout497 _6136_/C VGND VGND VPWR VPWR _6121_/B sky130_fd_sc_hd__buf_8
XFILLER_100_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input123_A wb_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5768__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6196__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3954__A1 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3954__B2 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6353__C1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6499__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output175_A _4160_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5171__A3 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_6_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__5459__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6656__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3890__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4920_ _5213_/A _5065_/A _5183_/C _4924_/B VGND VGND VPWR VPWR _4922_/A sky130_fd_sc_hd__and4_1
XFILLER_178_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6082__B _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4851_ _4851_/A _4851_/B _5294_/C VGND VGND VPWR VPWR _4851_/Y sky130_fd_sc_hd__nand3_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3802_ input5/X _3486_/X _3490_/X input13/X _3801_/X VGND VGND VPWR VPWR _3802_/X
+ sky130_fd_sc_hd__a221o_2
X_7570_ _7580_/CLK _7570_/D fanout745/X VGND VGND VPWR VPWR _7570_/Q sky130_fd_sc_hd__dfrtp_4
X_4782_ _4772_/A _4801_/B _5410_/A _5410_/B VGND VGND VPWR VPWR _4784_/B sky130_fd_sc_hd__and4b_1
XFILLER_119_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6521_ _6501_/X _6511_/X _6520_/X _6431_/Y _7281_/Q VGND VGND VPWR VPWR _6521_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3733_ _3686_/X _3689_/X _3733_/C _3733_/D VGND VGND VPWR VPWR _3733_/X sky130_fd_sc_hd__and4bb_2
XANTENNA_hold77_A hold77/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6452_ _7595_/Q _6466_/C _6462_/C _6466_/A VGND VGND VPWR VPWR _6452_/X sky130_fd_sc_hd__and4b_4
X_3664_ _4364_/A _5640_/B _5596_/A VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__and3_4
XFILLER_134_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5698__A1 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5403_ _5402_/X _5345_/Y _5322_/Y hold87/A _4428_/Y VGND VGND VPWR VPWR _7204_/D
+ sky130_fd_sc_hd__o32a_1
X_3595_ _7453_/Q _5848_/A _3529_/X _7533_/Q _3594_/X VGND VGND VPWR VPWR _3595_/X
+ sky130_fd_sc_hd__a221o_1
X_6383_ _6971_/Q _6074_/X _6317_/B _6382_/X _6380_/X VGND VGND VPWR VPWR _6383_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_133_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5334_ _5183_/B _5216_/A _5328_/X _5333_/X VGND VGND VPWR VPWR _5334_/X sky130_fd_sc_hd__a31o_1
XFILLER_142_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5265_ _5265_/A _5265_/B _5564_/A _5265_/D VGND VGND VPWR VPWR _5266_/B sky130_fd_sc_hd__nand4_1
Xhold2803 _4531_/X VGND VGND VPWR VPWR hold960/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2814 hold939/X VGND VGND VPWR VPWR _4487_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4984__C _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2825 hold997/X VGND VGND VPWR VPWR _4226_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_7004_ _7213_/CLK _7004_/D fanout700/X VGND VGND VPWR VPWR _7004_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2836 _7319_/Q VGND VGND VPWR VPWR hold2836/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4216_ _6839_/B _3481_/Y _4231_/S _4215_/X _5956_/C VGND VGND VPWR VPWR _4232_/S
+ sky130_fd_sc_hd__o221a_4
Xhold2847 _7303_/Q VGND VGND VPWR VPWR hold2847/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6662__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5196_ _4672_/X _4858_/Y _4980_/X _5044_/C _5195_/X VGND VGND VPWR VPWR _5196_/X
+ sky130_fd_sc_hd__o311a_1
Xhold2858 _7474_/Q VGND VGND VPWR VPWR hold2858/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2869 _7514_/Q VGND VGND VPWR VPWR hold2869/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4147_ _7266_/Q input78/X _4174_/B VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__mux2_8
XFILLER_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4078_ _4078_/A _4078_/B _4168_/D VGND VGND VPWR VPWR _4078_/Y sky130_fd_sc_hd__nor3_2
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout540_A hold1494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1488_A _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6719_ _7048_/Q _6435_/X _6446_/X _7189_/Q _6718_/X VGND VGND VPWR VPWR _6719_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3936__B2 _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4521__A _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4361__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4900__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6638__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4894__C _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4664__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5613__A1 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3624__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output292_A _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4431__A _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold709 hold709/A VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__7419__RESET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5144__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6629__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5050_ _5113_/A _5399_/C _5282_/C VGND VGND VPWR VPWR _5052_/B sky130_fd_sc_hd__and3_1
Xhold1409 hold4/X VGND VGND VPWR VPWR _4185_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5447__A4 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6644__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4655__A2 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4001_ _6910_/Q _6909_/Q VGND VGND VPWR VPWR _4001_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__6792__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4700__A_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5604__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4606__A _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5952_ _5952_/A0 _5952_/A1 _5955_/S VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3615__B1 _3549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4903_ _5065_/A _4907_/B _5049_/C _4940_/D VGND VGND VPWR VPWR _4903_/Y sky130_fd_sc_hd__nand4_1
X_5883_ _5883_/A0 _5955_/A1 _5883_/S VGND VGND VPWR VPWR _5883_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3630__A3 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7622_ _7625_/CLK _7622_/D fanout706/X VGND VGND VPWR VPWR _7622_/Q sky130_fd_sc_hd__dfrtp_1
X_4834_ _5127_/A _4834_/B VGND VGND VPWR VPWR _4834_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3918__A1 input96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7553_ _7581_/CLK _7553_/D fanout716/X VGND VGND VPWR VPWR _7553_/Q sky130_fd_sc_hd__dfrtp_2
X_4765_ _5260_/C _4765_/B _5059_/B VGND VGND VPWR VPWR _4766_/A sky130_fd_sc_hd__and3_1
XANTENNA__6580__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4979__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6504_ _7385_/Q _6413_/C _6426_/X _6451_/X _7481_/Q VGND VGND VPWR VPWR _6504_/X
+ sky130_fd_sc_hd__a32o_1
X_3716_ _7411_/Q _3493_/X hold41/A _7499_/Q _3715_/X VGND VGND VPWR VPWR _3716_/X
+ sky130_fd_sc_hd__a221o_2
X_7484_ _7574_/CLK _7484_/D fanout745/X VGND VGND VPWR VPWR _7484_/Q sky130_fd_sc_hd__dfrtp_4
X_4696_ _5297_/A _4696_/B VGND VGND VPWR VPWR _5531_/C sky130_fd_sc_hd__nand2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ _6441_/D _6466_/B _6467_/A _6466_/D VGND VGND VPWR VPWR _6435_/X sky130_fd_sc_hd__and4_4
X_3647_ _3647_/A _4515_/B _4539_/C VGND VGND VPWR VPWR _3647_/X sky130_fd_sc_hd__and3_4
XFILLER_134_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6366_ _6965_/Q _6144_/A _6144_/B _6079_/X _7014_/Q VGND VGND VPWR VPWR _6366_/X
+ sky130_fd_sc_hd__a32o_1
X_3578_ _7627_/Q _7254_/Q _7255_/Q VGND VGND VPWR VPWR _3578_/X sky130_fd_sc_hd__mux2_8
Xhold3301 _6625_/X VGND VGND VPWR VPWR _7621_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3312 _7072_/Q VGND VGND VPWR VPWR _4113_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3697__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3323 _7642_/Q VGND VGND VPWR VPWR _6816_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5317_ _5317_/A _5317_/B _5317_/C _5531_/A VGND VGND VPWR VPWR _5319_/A sky130_fd_sc_hd__nor4b_1
Xhold3334 _6066_/X VGND VGND VPWR VPWR _7601_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout490_A _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6297_ _7066_/Q _6110_/A _6332_/C _6119_/X _7132_/Q VGND VGND VPWR VPWR _6297_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout588_A hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3345 _6898_/Q VGND VGND VPWR VPWR _4048_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2600 _6963_/Q VGND VGND VPWR VPWR hold973/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6096__B2 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2611 _7065_/Q VGND VGND VPWR VPWR hold709/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3356 _6779_/X VGND VGND VPWR VPWR _7628_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3367 _6932_/Q VGND VGND VPWR VPWR _4112_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2622 hold989/X VGND VGND VPWR VPWR _5656_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5603__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2633 _7166_/Q VGND VGND VPWR VPWR hold751/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5248_ _5248_/A _5248_/B _5248_/C VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__and3_1
Xhold3378 _7257_/Q VGND VGND VPWR VPWR _4250_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2644 hold699/X VGND VGND VPWR VPWR _4348_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1910 hold174/X VGND VGND VPWR VPWR _5625_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__buf_6
Xhold2655 hold791/X VGND VGND VPWR VPWR _4496_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2666 hold725/X VGND VGND VPWR VPWR _5844_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1921 hold308/X VGND VGND VPWR VPWR _4368_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2677 _7097_/Q VGND VGND VPWR VPWR hold727/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1932 hold160/X VGND VGND VPWR VPWR _5973_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_188_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5179_ _5177_/Y _4986_/Y _5173_/X _5176_/X VGND VGND VPWR VPWR _5179_/Y sky130_fd_sc_hd__o211ai_2
Xhold1943 _7169_/Q VGND VGND VPWR VPWR hold403/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2688 _7014_/Q VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1954 _7306_/Q VGND VGND VPWR VPWR _4078_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1403_A _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2699 hold943/X VGND VGND VPWR VPWR _5828_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1965 _7028_/Q VGND VGND VPWR VPWR hold431/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1976 _7553_/Q VGND VGND VPWR VPWR hold449/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6399__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1987 _7033_/Q VGND VGND VPWR VPWR hold423/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1998 _7353_/Q VGND VGND VPWR VPWR hold417/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3420__A _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6434__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3909__B2 _7400_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6571__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5066__B _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6323__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5781__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input51_A mgmt_gpio_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3688__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5834__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3845__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4426__A _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output305_A _4166_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3612__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6562__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4550_ _5817_/A1 _4550_/A1 _4550_/S VGND VGND VPWR VPWR _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3501_ _5992_/A _5938_/A _3637_/C VGND VGND VPWR VPWR _3501_/X sky130_fd_sc_hd__and3_4
Xwire470 _4657_/A VGND VGND VPWR VPWR _4954_/A sky130_fd_sc_hd__clkbuf_8
Xhold506 hold506/A VGND VGND VPWR VPWR _7279_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4481_ _4481_/A0 _4553_/A0 _4484_/S VGND VGND VPWR VPWR _4481_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6314__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5117__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold517 hold517/A VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold528 hold528/A VGND VGND VPWR VPWR _6944_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6220_ _7348_/Q _6070_/X _6218_/X _6219_/X _6217_/X VGND VGND VPWR VPWR _6220_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold539 hold539/A VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3432_ _7386_/Q VGND VGND VPWR VPWR _3432_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5704__B _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3679__A3 _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _7409_/Q _6119_/D _6116_/C _6121_/B VGND VGND VPWR VPWR _6151_/X sky130_fd_sc_hd__o211a_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5453_/B _5102_/B VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__nand2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6112_/B _6120_/B _6082_/C VGND VGND VPWR VPWR _6082_/X sky130_fd_sc_hd__and3_4
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5825__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1206 hold2858/X VGND VGND VPWR VPWR hold2859/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1217 hold2893/X VGND VGND VPWR VPWR _7498_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5033_/A _5033_/B _5033_/C _5033_/D VGND VGND VPWR VPWR _5035_/D sky130_fd_sc_hd__nand4_1
Xhold1228 hold3177/X VGND VGND VPWR VPWR hold3178/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1239 _4488_/X VGND VGND VPWR VPWR _7144_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3836__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3851__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6984_ _7633_/CLK _6984_/D VGND VGND VPWR VPWR _6984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6250__B2 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5935_ _5998_/A1 _5935_/A1 _5937_/S VGND VGND VPWR VPWR _5935_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5866_ _5938_/A _5866_/B _5938_/B _5956_/C VGND VGND VPWR VPWR _5874_/S sky130_fd_sc_hd__and4_4
X_7605_ _7621_/CLK _7605_/D fanout705/X VGND VGND VPWR VPWR _7605_/Q sky130_fd_sc_hd__dfrtp_1
X_4817_ _5399_/C _5089_/B _5089_/C VGND VGND VPWR VPWR _4817_/X sky130_fd_sc_hd__and3_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5797_ _5968_/A1 _5797_/A1 _5802_/S VGND VGND VPWR VPWR _5797_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6553__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7536_ _7542_/CLK _7536_/D fanout708/X VGND VGND VPWR VPWR _7536_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5761__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4748_ _4748_/A _4844_/B _5091_/A VGND VGND VPWR VPWR _4748_/Y sky130_fd_sc_hd__nand3_4
XFILLER_135_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7467_ _7563_/CLK _7467_/D fanout739/X VGND VGND VPWR VPWR _7467_/Q sky130_fd_sc_hd__dfrtp_4
X_4679_ _4679_/A _4788_/C _4679_/C VGND VGND VPWR VPWR _4679_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6305__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4316__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6418_ _6455_/B _6574_/B _6459_/B VGND VGND VPWR VPWR _6419_/D sky130_fd_sc_hd__and3_4
X_7398_ _7579_/CLK hold49/X fanout731/X VGND VGND VPWR VPWR _7398_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5614__B _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6349_ _7023_/Q _6070_/X _6090_/X _7043_/Q _6348_/X VGND VGND VPWR VPWR _6349_/X
+ sky130_fd_sc_hd__a221o_1
Xhold3120 hold3120/A VGND VGND VPWR VPWR _4552_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3415__A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3131 hold3131/A VGND VGND VPWR VPWR _5840_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3142 _4480_/X VGND VGND VPWR VPWR hold3142/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6429__C _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR _4563_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3153 hold3153/A VGND VGND VPWR VPWR _5644_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR _4091_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3164 _5813_/X VGND VGND VPWR VPWR hold3164/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR input126/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2430 hold799/X VGND VGND VPWR VPWR _5756_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3175 hold3175/A VGND VGND VPWR VPWR _5582_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5816__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR _6817_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3186 hold3186/A VGND VGND VPWR VPWR _5620_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2441 hold581/X VGND VGND VPWR VPWR _5636_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR _6799_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3197 hold3197/A VGND VGND VPWR VPWR _4395_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2452 _7340_/Q VGND VGND VPWR VPWR hold957/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR _6815_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2463 _7435_/Q VGND VGND VPWR VPWR hold591/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2474 _4529_/X VGND VGND VPWR VPWR hold882/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1740 _4332_/X VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2485 _4517_/X VGND VGND VPWR VPWR hold886/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2496 _7010_/Q VGND VGND VPWR VPWR hold735/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1751 _5789_/X VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1762 hold148/X VGND VGND VPWR VPWR _4438_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1773 hold373/X VGND VGND VPWR VPWR _5832_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1784 _7560_/Q VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1795 _4207_/X VGND VGND VPWR VPWR hold121/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3842__A3 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1987_A _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input99_A wb_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3763__C1 _3762_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4307__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5807__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3833__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6232__A1 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6232__B2 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3981_ _7056_/Q _5947_/B _5623_/B _7447_/Q _5848_/A VGND VGND VPWR VPWR _3981_/X
+ sky130_fd_sc_hd__a32o_1
X_5720_ _5954_/A1 _5720_/A1 _5721_/S VGND VGND VPWR VPWR _5720_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5651_ _5894_/A0 _5651_/A1 _5658_/S VGND VGND VPWR VPWR _5651_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4603__B _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_51_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6535__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2370_A _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4602_ _4772_/A _4772_/B VGND VGND VPWR VPWR _5260_/A sky130_fd_sc_hd__nor2_8
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5582_ _5582_/A0 _5582_/A1 _5586_/S VGND VGND VPWR VPWR _5582_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7321_ _7539_/CLK _7321_/D fanout708/X VGND VGND VPWR VPWR _7321_/Q sky130_fd_sc_hd__dfrtp_4
X_4533_ _4533_/A _4533_/B VGND VGND VPWR VPWR _4538_/S sky130_fd_sc_hd__nand2_4
Xhold303 hold303/A VGND VGND VPWR VPWR _7323_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold314 hold314/A VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6299__B2 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold325 hold325/A VGND VGND VPWR VPWR _7560_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7252_ _7263_/CLK _7252_/D fanout689/X VGND VGND VPWR VPWR _7252_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_171_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ _4464_/A0 _5914_/A1 _4466_/S VGND VGND VPWR VPWR _4464_/X sky130_fd_sc_hd__mux2_1
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3793__A_N _3764_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold347 hold347/A VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold358 hold358/A VGND VGND VPWR VPWR _7352_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6203_ _7331_/Q _6384_/A4 _6097_/C _6388_/A3 _7371_/Q VGND VGND VPWR VPWR _6203_/X
+ sky130_fd_sc_hd__a32o_1
X_3415_ _7522_/Q VGND VGND VPWR VPWR _3415_/Y sky130_fd_sc_hd__inv_2
X_7183_ _7185_/CLK _7183_/D fanout737/X VGND VGND VPWR VPWR _7183_/Q sky130_fd_sc_hd__dfrtp_4
X_4395_ _5582_/A0 _4395_/A1 _4399_/S VGND VGND VPWR VPWR _4395_/X sky130_fd_sc_hd__mux2_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ _7360_/Q _6276_/A3 _6267_/B1 _7392_/Q VGND VGND VPWR VPWR _6134_/X sky130_fd_sc_hd__a22o_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1003 hold3037/X VGND VGND VPWR VPWR hold3038/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _7586_/Q _7587_/Q _6065_/C VGND VGND VPWR VPWR _6065_/Y sky130_fd_sc_hd__nor3_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 hold3005/X VGND VGND VPWR VPWR _7257_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1025 hold3057/X VGND VGND VPWR VPWR _7431_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1036 hold3062/X VGND VGND VPWR VPWR _7243_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1047 hold3072/X VGND VGND VPWR VPWR hold3073/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5016_ _4956_/A _5012_/Y _5014_/Y _5011_/Y VGND VGND VPWR VPWR _5016_/Y sky130_fd_sc_hd__o211ai_1
Xhold1058 hold3105/X VGND VGND VPWR VPWR hold3106/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1069 hold1069/A VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3824__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout453_A hold40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6223__A1 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _7212_/CLK _6967_/D fanout724/X VGND VGND VPWR VPWR _6967_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5918_ _5918_/A0 _5990_/A1 _5919_/S VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3588__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5982__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6898_ _7075_/CLK _6898_/D _6848_/X VGND VGND VPWR VPWR _6898_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout718_A fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5849_ _5912_/A1 _5849_/A1 _5856_/S VGND VGND VPWR VPWR _5849_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5329__A3 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6526__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold1568_A _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7519_ _7519_/CLK _7519_/D fanout741/X VGND VGND VPWR VPWR _7519_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_163_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3760__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold870 hold870/A VGND VGND VPWR VPWR _7014_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold881 hold881/A VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold892 _4482_/X VGND VGND VPWR VPWR _7139_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5063__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input153_A wb_dat_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2260 hold613/X VGND VGND VPWR VPWR _5744_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2271 _7426_/Q VGND VGND VPWR VPWR hold665/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2282 _7542_/Q VGND VGND VPWR VPWR hold575/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2293 _7404_/Q VGND VGND VPWR VPWR hold789/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1570 hold262/X VGND VGND VPWR VPWR _6950_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input14_A mask_rev_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1581 _7204_/Q VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1592 _7510_/Q VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_60_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6765__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3579__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3751__A2 _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6150__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4180_ _4551_/B _5938_/B _4388_/B _4533_/B VGND VGND VPWR VPWR _4190_/S sky130_fd_sc_hd__and4_2
XFILLER_121_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6453__A1 _7479_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6453__B2 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6085__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6205__A1 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6205__B2 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6821_ _7109_/Q _6821_/A2 _6821_/B1 wire536/A _6820_/X VGND VGND VPWR VPWR _6821_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4216__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6756__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6752_ _6751_/X _6776_/A2 _6777_/S VGND VGND VPWR VPWR _7626_/D sky130_fd_sc_hd__mux2_1
X_3964_ _7431_/Q _3525_/X _3537_/X _7423_/Q _3963_/X VGND VGND VPWR VPWR _3964_/X
+ sky130_fd_sc_hd__a221o_1
X_5703_ _5703_/A0 _6000_/A1 _5703_/S VGND VGND VPWR VPWR _5703_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6683_ _7057_/Q _6447_/C _6769_/A3 _6447_/X _7183_/Q VGND VGND VPWR VPWR _6683_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3895_ _7472_/Q _3494_/X _5857_/A _7456_/Q _3894_/X VGND VGND VPWR VPWR _3895_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5716__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4519__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5634_ _5634_/A _5956_/C VGND VGND VPWR VPWR _5639_/S sky130_fd_sc_hd__nand2_4
XANTENNA__3990__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5565_ _5562_/Y _5564_/Y _5560_/X VGND VGND VPWR VPWR _5565_/X sky130_fd_sc_hd__o21a_1
XFILLER_145_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4987__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold100 hold100/A VGND VGND VPWR VPWR _7574_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7304_ _7542_/CLK _7304_/D fanout708/X VGND VGND VPWR VPWR _7304_/Q sky130_fd_sc_hd__dfrtp_4
X_4516_ _4516_/A0 _5582_/A0 _4520_/S VGND VGND VPWR VPWR _4516_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3742__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold111 hold111/A VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold122 _7207_/Q VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5496_ _5496_/A _5496_/B _5496_/C VGND VGND VPWR VPWR _5529_/C sky130_fd_sc_hd__and3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold144 hold144/A VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7235_ _7238_/CLK _7235_/D fanout690/X VGND VGND VPWR VPWR _7235_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_105_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold155 hold155/A VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4447_ _4447_/A0 _4447_/A1 _4448_/S VGND VGND VPWR VPWR _4447_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold166 hold166/A VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6141__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold188 hold188/A VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold199 hold199/A VGND VGND VPWR VPWR _7408_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5495__A2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout613 _6433_/D VGND VGND VPWR VPWR _6466_/B sky130_fd_sc_hd__buf_6
XFILLER_59_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout624 _7590_/Q VGND VGND VPWR VPWR _6081_/C sky130_fd_sc_hd__buf_6
XANTENNA__6692__B2 _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7166_ _7212_/CLK _7166_/D fanout724/X VGND VGND VPWR VPWR _7166_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout635 _6067_/B VGND VGND VPWR VPWR _6019_/A sky130_fd_sc_hd__buf_8
X_4378_ _4378_/A0 _4547_/A0 _4381_/S VGND VGND VPWR VPWR _4378_/X sky130_fd_sc_hd__mux2_1
Xfanout646 _4918_/D VGND VGND VPWR VPWR _5342_/B sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_1_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7250_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout657 _5094_/A VGND VGND VPWR VPWR _5089_/D sky130_fd_sc_hd__buf_12
XANTENNA_input6_A mask_rev_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6117_ _6144_/C _6116_/C _6144_/B _6116_/X _7311_/Q VGND VGND VPWR VPWR _6117_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout570_A _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7097_ _7197_/CLK _7097_/D fanout742/X VGND VGND VPWR VPWR _7097_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5180__A _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6444__A1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6444__B2 _7327_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _7594_/Q _6429_/C _6433_/D VGND VGND VPWR VPWR _6048_/X sky130_fd_sc_hd__a21o_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5707__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3981__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6132__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold3233_A _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6683__B2 _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2090 _7062_/Q VGND VGND VPWR VPWR hold314/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_799 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6738__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4749__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3972__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3680_ _7363_/Q _3564_/X _3648_/X _7040_/Q _3679_/X VGND VGND VPWR VPWR _3680_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_185_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5174__A1 _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5350_ _5089_/D _4939_/C _4891_/D _5065_/A VGND VGND VPWR VPWR _5350_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3724__A2 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput205 _4141_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput216 _7655_/X VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
Xoutput227 _7664_/X VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_142_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput238 _4139_/X VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
X_4301_ _3607_/Y _4301_/A1 _4302_/S VGND VGND VPWR VPWR _6986_/D sky130_fd_sc_hd__mux2_1
XFILLER_142_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput249 _4133_/X VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
X_5281_ _4836_/A _5282_/D _5134_/C _5280_/X VGND VGND VPWR VPWR _5281_/X sky130_fd_sc_hd__a31o_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7020_ _7213_/CLK _7020_/D fanout702/X VGND VGND VPWR VPWR _7020_/Q sky130_fd_sc_hd__dfrtp_4
X_4232_ _4232_/A0 _4231_/X _4232_/S VGND VGND VPWR VPWR _4232_/X sky130_fd_sc_hd__mux2_1
X_4163_ _7092_/Q _4163_/A1 _7261_/Q VGND VGND VPWR VPWR _4163_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4094_ _4825_/A _4674_/A _4564_/A _4564_/B VGND VGND VPWR VPWR _4095_/D sky130_fd_sc_hd__a211oi_1
XANTENNA__4328__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6729__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6804_ _6803_/X _6804_/A1 _6822_/S VGND VGND VPWR VPWR _7638_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5937__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4996_ _4996_/A _5339_/A _5203_/C _5034_/B VGND VGND VPWR VPWR _5033_/D sky130_fd_sc_hd__nand4_1
XANTENNA__5401__A2 _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6735_ _7029_/Q _6459_/B _6459_/C _6451_/X _6877_/Q VGND VGND VPWR VPWR _6735_/X
+ sky130_fd_sc_hd__a32o_1
X_3947_ _7235_/Q _5619_/A _5632_/B _3542_/X _6919_/Q VGND VGND VPWR VPWR _3947_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6666_ _7167_/Q _6408_/D _6657_/X _6662_/X _6665_/X VGND VGND VPWR VPWR _6666_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3963__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3878_ _7037_/Q _3648_/X _3659_/X _7007_/Q _3877_/X VGND VGND VPWR VPWR _3879_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout416_A hold47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5617_ _5617_/A0 _5995_/A1 _5618_/S VGND VGND VPWR VPWR _5617_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5165__B2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6597_ _6595_/X _6430_/X _6587_/X _6596_/X VGND VGND VPWR VPWR _6597_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3715__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5548_ _5548_/A _5548_/B _5575_/B VGND VGND VPWR VPWR _5548_/Y sky130_fd_sc_hd__nand3_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6114__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5479_ _4679_/Y _4814_/Y _4971_/X _5478_/Y VGND VGND VPWR VPWR _5482_/B sky130_fd_sc_hd__o31a_1
XANTENNA__6665__A1 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7218_ _4150_/A1 _7218_/D _6870_/X VGND VGND VPWR VPWR _7218_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_48_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout410 _5695_/A VGND VGND VPWR VPWR _3872_/A2 sky130_fd_sc_hd__buf_4
Xfanout421 _4924_/B VGND VGND VPWR VPWR _4933_/A sky130_fd_sc_hd__clkbuf_8
Xfanout443 _3860_/D VGND VGND VPWR VPWR _4515_/B sky130_fd_sc_hd__buf_8
Xfanout454 hold39/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__buf_6
X_7149_ _7395_/CLK _7149_/D fanout738/X VGND VGND VPWR VPWR _7149_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_101_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3423__A _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout465 _5038_/B VGND VGND VPWR VPWR _5034_/B sky130_fd_sc_hd__buf_4
XFILLER_171_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout476 _6428_/X VGND VGND VPWR VPWR _6459_/C sky130_fd_sc_hd__buf_8
XFILLER_86_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout487 _6116_/A VGND VGND VPWR VPWR _6120_/B sky130_fd_sc_hd__buf_6
Xfanout498 _6136_/C VGND VGND VPWR VPWR _6144_/B sky130_fd_sc_hd__buf_8
XFILLER_171_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input116_A wb_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__A0 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5069__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5784__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3954__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input81_A spi_sdo VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4701__B _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold3350_A _7221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5459__A2 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4850_ _5295_/D _4850_/B _5029_/A _5295_/A VGND VGND VPWR VPWR _5294_/C sky130_fd_sc_hd__nand4_4
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6082__C _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6187__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ _3485_/X _5612_/C _4491_/C _3501_/X _7577_/Q VGND VGND VPWR VPWR _3801_/X
+ sky130_fd_sc_hd__a32o_2
X_4781_ _4781_/A _4781_/B VGND VGND VPWR VPWR _4781_/Y sky130_fd_sc_hd__nor2_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6520_ _7409_/Q _6468_/X _6430_/X _6519_/X _6516_/X VGND VGND VPWR VPWR _6520_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3945__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3732_ _3732_/A _3732_/B _3732_/C _3732_/D VGND VGND VPWR VPWR _3733_/D sky130_fd_sc_hd__nor4_2
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6451_ _6466_/B _6467_/A _6600_/B _6466_/A VGND VGND VPWR VPWR _6451_/X sky130_fd_sc_hd__and4b_4
XFILLER_174_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6344__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3663_ _4551_/B _4515_/B _4509_/C VGND VGND VPWR VPWR _3663_/X sky130_fd_sc_hd__and3_4
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3508__A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5402_ _5374_/X _5401_/X _5402_/B1 _5372_/X VGND VGND VPWR VPWR _5402_/X sky130_fd_sc_hd__a211o_1
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6382_ _7116_/Q _6317_/C _6089_/X _7045_/Q _6381_/X VGND VGND VPWR VPWR _6382_/X
+ sky130_fd_sc_hd__a221o_1
X_3594_ _7397_/Q _5803_/A _3933_/A _3519_/X _7549_/Q VGND VGND VPWR VPWR _3594_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5333_ _5053_/C _5216_/A _5328_/X _5332_/X VGND VGND VPWR VPWR _5333_/X sky130_fd_sc_hd__a31o_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5264_ _4772_/B _5079_/B _5102_/B _5263_/X VGND VGND VPWR VPWR _5265_/D sky130_fd_sc_hd__a31oi_2
Xhold2804 _6912_/Q VGND VGND VPWR VPWR hold773/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_7003_ _7164_/CLK _7003_/D fanout698/X VGND VGND VPWR VPWR _7003_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_87_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2815 _7130_/Q VGND VGND VPWR VPWR hold991/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4215_ _4078_/A _4078_/B _4168_/D _5785_/B _5992_/C VGND VGND VPWR VPWR _4215_/X
+ sky130_fd_sc_hd__o311a_2
Xhold2826 _4226_/X VGND VGND VPWR VPWR hold998/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2837 hold2837/A VGND VGND VPWR VPWR _5705_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2848 hold2848/A VGND VGND VPWR VPWR _5687_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5195_ _4672_/X _5174_/Y _4986_/Y _5169_/X _5194_/Y VGND VGND VPWR VPWR _5195_/X
+ sky130_fd_sc_hd__o311a_1
Xhold2859 hold2859/A VGND VGND VPWR VPWR _5879_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4146_ _7265_/Q input80/X _4174_/B VGND VGND VPWR VPWR _4146_/X sky130_fd_sc_hd__mux2_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4077_ _3400_/Y _4076_/C _4076_/X VGND VGND VPWR VPWR _6882_/D sky130_fd_sc_hd__o21bai_1
XANTENNA__5083__B1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A hold31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5622__A2 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3633__B2 _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5386__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4979_ _4996_/A _5328_/A _5328_/B VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__and3_2
XANTENNA__6583__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6718_ _7184_/Q _6466_/C _6574_/C _6443_/X _7194_/Q VGND VGND VPWR VPWR _6718_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_50_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6649_ _6648_/X _6649_/A1 _6649_/S VGND VGND VPWR VPWR _6649_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6335__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3418__A _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6350__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7525_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_180_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5310__A1 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_csclk _7399_/CLK VGND VGND VPWR VPWR _7582_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_93_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5779__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6326__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire674 _4604_/Y VGND VGND VPWR VPWR wire674/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3560__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6629__A1 _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6629__B2 hold52/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5301__A1 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4159__A input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4000_ _6909_/Q _4006_/A _4000_/B1 VGND VGND VPWR VPWR _4003_/A sky130_fd_sc_hd__a21oi_1
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5951_ _5951_/A0 _5951_/A1 _5955_/S VGND VGND VPWR VPWR _5951_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3615__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4606__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3615__B2 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5080__A3 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4902_ _4902_/A _4902_/B _5448_/D _5223_/D VGND VGND VPWR VPWR _4904_/B sky130_fd_sc_hd__nand4_1
X_5882_ _5882_/A0 _5999_/A1 _5883_/S VGND VGND VPWR VPWR _5882_/X sky130_fd_sc_hd__mux2_1
X_7621_ _7621_/CLK _7621_/D fanout711/X VGND VGND VPWR VPWR _7621_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4833_ _4833_/A _4834_/B _5295_/A VGND VGND VPWR VPWR _4839_/B sky130_fd_sc_hd__and3_1
XANTENNA__6565__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2665_A _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7552_ _7582_/CLK _7552_/D fanout717/X VGND VGND VPWR VPWR _7552_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3918__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4764_ _4700_/Y _4727_/Y _4718_/Y _4763_/Y VGND VGND VPWR VPWR _4766_/B sky130_fd_sc_hd__o211ai_1
XFILLER_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6503_ _7353_/Q _6413_/C _6459_/C _6408_/B _7377_/Q VGND VGND VPWR VPWR _6503_/X
+ sky130_fd_sc_hd__a32o_1
X_3715_ _6915_/Q _5612_/B _5947_/A _3515_/X _7239_/Q VGND VGND VPWR VPWR _3715_/X
+ sky130_fd_sc_hd__a32o_2
X_7483_ _7563_/CLK _7483_/D fanout740/X VGND VGND VPWR VPWR _7483_/Q sky130_fd_sc_hd__dfrtp_4
X_4695_ _4802_/A _4794_/A VGND VGND VPWR VPWR _4695_/Y sky130_fd_sc_hd__nand2_2
X_6434_ _6455_/B _6434_/B _6600_/B VGND VGND VPWR VPWR _6434_/X sky130_fd_sc_hd__and3_4
XFILLER_174_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3646_ _4328_/A _5596_/A _4346_/C VGND VGND VPWR VPWR _4322_/A sky130_fd_sc_hd__and3_4
X_6365_ _7195_/Q _6144_/A _6097_/C _6364_/X VGND VGND VPWR VPWR _6365_/X sky130_fd_sc_hd__a31o_1
X_3577_ _4388_/B _5596_/B _5640_/C VGND VGND VPWR VPWR _5630_/S sky130_fd_sc_hd__and3_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4995__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3302 _7616_/Q VGND VGND VPWR VPWR _6522_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3551__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5316_ _4605_/Y _4625_/Y _4731_/Y _4755_/Y _4814_/Y VGND VGND VPWR VPWR _5531_/A
+ sky130_fd_sc_hd__o32a_1
Xhold3313 _4113_/X VGND VGND VPWR VPWR _7072_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3324 _7627_/Q VGND VGND VPWR VPWR _6777_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6296_ _7177_/Q _6092_/X _6295_/X _6294_/X _6293_/X VGND VGND VPWR VPWR _6303_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold3335 _7205_/Q VGND VGND VPWR VPWR _5484_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3346 _4048_/X VGND VGND VPWR VPWR _6898_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2601 hold973/X VGND VGND VPWR VPWR _4267_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2612 hold709/X VGND VGND VPWR VPWR _4399_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3357 _6904_/Q VGND VGND VPWR VPWR _4033_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ _5419_/A _5247_/B _5247_/C VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__and3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3368 _4112_/X VGND VGND VPWR VPWR _6929_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2623 _5656_/X VGND VGND VPWR VPWR hold990/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3379 _7205_/Q VGND VGND VPWR VPWR hold103/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2634 hold751/X VGND VGND VPWR VPWR _4514_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__buf_12
Xhold2645 _4348_/X VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1900 _6965_/Q VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1911 _5625_/X VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2656 _7493_/Q VGND VGND VPWR VPWR hold893/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1922 _4368_/X VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_46_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__buf_6
Xhold2667 _7126_/Q VGND VGND VPWR VPWR hold739/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1933 _5973_/X VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5178_ _5203_/C _5183_/C _5216_/A VGND VGND VPWR VPWR _5178_/X sky130_fd_sc_hd__o21a_1
Xhold2678 hold727/X VGND VGND VPWR VPWR _4445_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1944 hold403/X VGND VGND VPWR VPWR _4518_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2689 hold869/X VGND VGND VPWR VPWR _4338_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1955 _5690_/X VGND VGND VPWR VPWR hold366/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4129_ _6897_/Q _4129_/B VGND VGND VPWR VPWR _4130_/A sky130_fd_sc_hd__nand2b_2
Xhold1966 hold431/X VGND VGND VPWR VPWR _4355_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1977 hold449/X VGND VGND VPWR VPWR _5968_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout748_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1988 hold423/X VGND VGND VPWR VPWR _4361_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1999 hold417/X VGND VGND VPWR VPWR _5743_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1598_A _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6556__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3909__A2 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6308__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6323__A3 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A mgmt_gpio_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5598__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4426__B _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4270__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3410__1_A _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6547__B1 _6545_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5770__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5972__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3500_ _3511_/A _3500_/B _3511_/C VGND VGND VPWR VPWR _3500_/X sky130_fd_sc_hd__and3_4
XFILLER_116_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4480_ _4480_/A0 _5912_/A1 _4484_/S VGND VGND VPWR VPWR _4480_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold518 _5877_/X VGND VGND VPWR VPWR _7472_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3431_ _7394_/Q VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3533__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3679__A4 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6150_ _7513_/Q _6080_/A _6317_/C _6087_/X _7465_/Q VGND VGND VPWR VPWR _6150_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5407_/A1 _5091_/A _5100_/X _5099_/Y VGND VGND VPWR VPWR _5101_/Y sky130_fd_sc_hd__a31oi_2
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _7589_/Q _6099_/D _6081_/C _7588_/Q VGND VGND VPWR VPWR _6081_/X sky130_fd_sc_hd__and4bb_4
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1207 _5879_/X VGND VGND VPWR VPWR _7474_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4984_/B _4984_/A _4660_/Y _4862_/X _4759_/Y VGND VGND VPWR VPWR _5033_/B
+ sky130_fd_sc_hd__a2111o_1
Xhold1218 hold2874/X VGND VGND VPWR VPWR hold2875/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1229 hold3179/X VGND VGND VPWR VPWR _6933_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3521__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5589__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6983_ _7000_/CLK _6983_/D VGND VGND VPWR VPWR _6983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5934_ _5979_/A0 _5934_/A1 _5937_/S VGND VGND VPWR VPWR _5934_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4261__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5865_ hold20/X _5865_/A1 _5865_/S VGND VGND VPWR VPWR _5865_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7604_ _7625_/CLK _7604_/D fanout705/X VGND VGND VPWR VPWR _7604_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4352__A _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4816_ _5410_/A _5061_/B _5399_/C VGND VGND VPWR VPWR _4818_/B sky130_fd_sc_hd__and3_1
XFILLER_167_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5796_ _5949_/A1 _5796_/A1 _5802_/S VGND VGND VPWR VPWR _5796_/X sky130_fd_sc_hd__mux2_1
X_4747_ _4879_/D _4747_/B _4887_/B _4945_/A VGND VGND VPWR VPWR _5094_/A sky130_fd_sc_hd__and4b_4
X_7535_ _7537_/CLK _7535_/D fanout707/X VGND VGND VPWR VPWR _7535_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5882__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7466_ _7522_/CLK _7466_/D fanout743/X VGND VGND VPWR VPWR _7466_/Q sky130_fd_sc_hd__dfrtp_4
X_4678_ _4679_/A _4788_/C _4679_/C VGND VGND VPWR VPWR _5342_/A sky130_fd_sc_hd__and3_4
X_6417_ _6427_/A _6434_/B _6468_/C VGND VGND VPWR VPWR _6419_/C sky130_fd_sc_hd__and3_4
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3629_ _7412_/Q _3493_/X _5686_/A _7308_/Q _3628_/X VGND VGND VPWR VPWR _3632_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4316__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6710__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7397_ _7582_/CLK _7397_/D fanout718/X VGND VGND VPWR VPWR _7397_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5614__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6348_ _7211_/Q _6332_/B _6089_/X _6100_/X _7063_/Q VGND VGND VPWR VPWR _6348_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_143_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3110 _4450_/X VGND VGND VPWR VPWR hold3110/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3121 _4552_/X VGND VGND VPWR VPWR hold3121/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3132 _7117_/Q VGND VGND VPWR VPWR hold3132/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6069__A2 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3143 _7041_/Q VGND VGND VPWR VPWR hold3143/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR _4563_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_6279_ _7350_/Q _6070_/X _6082_/X _7326_/Q _6278_/X VGND VGND VPWR VPWR _6280_/D
+ sky130_fd_sc_hd__a221o_1
Xhold3154 _7182_/Q VGND VGND VPWR VPWR hold3154/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR input116/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2420 _7285_/Q VGND VGND VPWR VPWR hold771/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3165 _7559_/Q VGND VGND VPWR VPWR hold3165/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR input127/X sky130_fd_sc_hd__clkbuf_2
Xhold2431 _7348_/Q VGND VGND VPWR VPWR hold901/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3176 _5582_/X VGND VGND VPWR VPWR hold3176/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5911__A _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR _6820_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3187 _5620_/X VGND VGND VPWR VPWR hold3187/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2442 _5636_/X VGND VGND VPWR VPWR hold582/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR _6802_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3198 _6962_/Q VGND VGND VPWR VPWR hold3198/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2453 hold957/X VGND VGND VPWR VPWR _5728_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2464 hold591/X VGND VGND VPWR VPWR _5835_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1730 hold421/X VGND VGND VPWR VPWR _4433_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2475 _7388_/Q VGND VGND VPWR VPWR hold925/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1741 hold233/X VGND VGND VPWR VPWR _7009_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2486 _7193_/Q VGND VGND VPWR VPWR hold907/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1752 _7298_/Q VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4527__A _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2497 hold735/X VGND VGND VPWR VPWR _4333_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1763 _4438_/X VGND VGND VPWR VPWR hold149/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1774 _5832_/X VGND VGND VPWR VPWR hold374/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3431__A _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1785 hold324/X VGND VGND VPWR VPWR _5976_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1796 hold121/X VGND VGND VPWR VPWR _6922_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6241__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4252__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5752__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5792__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6480__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6768__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5967__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6232__A2 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3980_ _7036_/Q _3648_/X _4545_/A _7192_/Q _3927_/X VGND VGND VPWR VPWR _3980_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3597__A3 _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5991__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5650_ _5650_/A1 hold365/X _4168_/D _4248_/S _5947_/C VGND VGND VPWR VPWR _5658_/S
+ sky130_fd_sc_hd__o311ai_4
XFILLER_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6090__C _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4601_ _5091_/A _5399_/A VGND VGND VPWR VPWR _4601_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__5743__A1 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5581_ _5581_/A _5619_/C VGND VGND VPWR VPWR _5586_/S sky130_fd_sc_hd__nand2_4
XFILLER_157_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7320_ _7542_/CLK _7320_/D fanout708/X VGND VGND VPWR VPWR _7320_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A0 _5817_/A1 _4532_/S VGND VGND VPWR VPWR _4532_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold52_A hold52/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7251_ _7263_/CLK _7251_/D fanout692/X VGND VGND VPWR VPWR _7251_/Q sky130_fd_sc_hd__dfrtp_4
Xhold315 _4396_/X VGND VGND VPWR VPWR _7062_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4463_ _4463_/A0 _4553_/A0 _4466_/S VGND VGND VPWR VPWR _4463_/X sky130_fd_sc_hd__mux2_1
Xhold337 hold337/A VGND VGND VPWR VPWR _7330_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold348 hold348/A VGND VGND VPWR VPWR _7528_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6202_ _7523_/Q _6379_/B1 _6200_/X _6201_/X VGND VGND VPWR VPWR _6202_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3516__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3414_ _7530_/Q VGND VGND VPWR VPWR _3414_/Y sky130_fd_sc_hd__inv_2
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7182_ _7184_/CLK _7182_/D fanout725/X VGND VGND VPWR VPWR _7182_/Q sky130_fd_sc_hd__dfrtp_4
X_4394_ _4394_/A _5619_/C VGND VGND VPWR VPWR _4399_/S sky130_fd_sc_hd__nand2_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _6075_/A _6130_/X _6132_/X _6126_/X _6128_/X VGND VGND VPWR VPWR _6133_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_124_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5731__A _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6064_ _6064_/A1 _6062_/X _6063_/X VGND VGND VPWR VPWR _7600_/D sky130_fd_sc_hd__a21bo_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1004 hold3039/X VGND VGND VPWR VPWR hold3040/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 hold2833/X VGND VGND VPWR VPWR hold2834/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1026 hold3065/X VGND VGND VPWR VPWR hold3066/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5038_/A _5216_/A _5030_/C _5013_/X VGND VGND VPWR VPWR _5015_/X sky130_fd_sc_hd__a31o_1
Xhold1037 hold3102/X VGND VGND VPWR VPWR hold3103/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1048 hold3074/X VGND VGND VPWR VPWR _7011_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1059 hold3107/X VGND VGND VPWR VPWR _7132_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4482__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6759__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5877__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6223__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4234__A1 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6966_ _7180_/CLK _6966_/D fanout721/X VGND VGND VPWR VPWR _6966_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_fanout446_A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5431__B1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5917_ _5917_/A0 _5980_/A0 _5919_/S VGND VGND VPWR VPWR _5917_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3588__A3 _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6897_ _7075_/CLK _6897_/D _6847_/X VGND VGND VPWR VPWR _6897_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3993__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5848_ _5848_/A _5956_/C VGND VGND VPWR VPWR _5856_/S sky130_fd_sc_hd__nand2_8
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5734__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5779_ _5968_/A1 _5779_/A1 _5784_/S VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold1463_A _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7518_ _7565_/CLK _7518_/D fanout748/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfrtp_4
XFILLER_107_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7449_ _7519_/CLK _7449_/D fanout742/X VGND VGND VPWR VPWR _7449_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3760__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold860 _5898_/X VGND VGND VPWR VPWR _7491_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold871 hold871/A VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold882 hold882/A VGND VGND VPWR VPWR _7178_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold893 hold893/A VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input146_A wb_dat_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2250 _7233_/Q VGND VGND VPWR VPWR hold571/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6907__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2261 _5744_/X VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2272 hold665/X VGND VGND VPWR VPWR _5825_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2283 hold575/X VGND VGND VPWR VPWR _5955_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2294 hold789/X VGND VGND VPWR VPWR _5800_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1560 _7444_/Q VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5670__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1571 _7509_/Q VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1582 hold87/X VGND VGND VPWR VPWR _3463_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1593 hold97/X VGND VGND VPWR VPWR _5919_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5787__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4225__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3579__A3 _3578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5973__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3984__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6517__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5725__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3751__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6150__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6150__B2 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6453__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4464__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5697__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6205__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A3 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6820_ _4427_/D _6820_/A2 _6820_/B1 _4427_/C VGND VGND VPWR VPWR _6820_/X sky130_fd_sc_hd__a22o_1
XFILLER_51_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4216__A1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6756__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6751_ _6750_/X _6751_/A1 _6751_/S VGND VGND VPWR VPWR _6751_/X sky130_fd_sc_hd__mux2_1
X_3963_ _7257_/Q _5965_/A _4352_/B _3669_/X _6967_/Q VGND VGND VPWR VPWR _3963_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5964__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5702_ _5702_/A0 _5954_/A1 _5703_/S VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__mux2_1
X_6682_ _7128_/Q _6424_/X _6677_/X _6681_/X _6430_/X VGND VGND VPWR VPWR _6682_/X
+ sky130_fd_sc_hd__a2111o_1
X_3894_ _7057_/Q _4376_/B _4364_/B _3663_/X _7163_/Q VGND VGND VPWR VPWR _3894_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_176_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6508__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5633_ _5633_/A0 _5993_/A1 _5633_/S VGND VGND VPWR VPWR _5633_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5564_ _5564_/A _5564_/B _5564_/C VGND VGND VPWR VPWR _5564_/Y sky130_fd_sc_hd__nand3_2
XFILLER_191_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7303_ _7309_/CLK _7303_/D fanout704/X VGND VGND VPWR VPWR _7303_/Q sky130_fd_sc_hd__dfstp_4
X_4515_ _5938_/B _4515_/B _4527_/A _4551_/D VGND VGND VPWR VPWR _4520_/S sky130_fd_sc_hd__and4_4
Xhold101 hold101/A VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold123 _3459_/A VGND VGND VPWR VPWR _3511_/C sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3742__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5495_ _4956_/A _4956_/B _4595_/Y _5495_/C1 VGND VGND VPWR VPWR _5529_/B sky130_fd_sc_hd__a211o_1
XANTENNA_hold2912_A _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold134 hold134/A VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold145 hold145/A VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4446_ _4446_/A0 _4446_/A1 _4448_/S VGND VGND VPWR VPWR _4446_/X sky130_fd_sc_hd__mux2_1
Xhold156 hold156/A VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7234_ _7255_/CLK _7234_/D fanout688/X VGND VGND VPWR VPWR _7234_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6141__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold167 hold167/A VGND VGND VPWR VPWR _7253_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4152__A0 _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold178 hold178/A VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold189 hold189/A VGND VGND VPWR VPWR _6951_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7165_ _7181_/CLK _7165_/D fanout721/X VGND VGND VPWR VPWR _7165_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__6692__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout614 _7595_/Q VGND VGND VPWR VPWR _6433_/D sky130_fd_sc_hd__clkbuf_8
X_4377_ _4377_/A0 _5876_/A1 _4381_/S VGND VGND VPWR VPWR _4377_/X sky130_fd_sc_hd__mux2_1
Xfanout625 _7590_/Q VGND VGND VPWR VPWR _6119_/B sky130_fd_sc_hd__buf_6
XANTENNA_fanout396_A _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout636 hold3353/X VGND VGND VPWR VPWR _6067_/B sky130_fd_sc_hd__clkbuf_8
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6116_/A _6119_/D _6116_/C VGND VGND VPWR VPWR _6116_/X sky130_fd_sc_hd__and3_4
Xfanout647 _4970_/C VGND VGND VPWR VPWR _5180_/B sky130_fd_sc_hd__buf_8
X_7096_ _7267_/CLK _7096_/D fanout749/X VGND VGND VPWR VPWR _7096_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5180__B _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6047_ _6433_/D _6434_/B VGND VGND VPWR VPWR _6047_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6444__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout563_A _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout730_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4207__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5955__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6949_ _7575_/CLK _6949_/D fanout735/X VGND VGND VPWR VPWR _6949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3966__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3981__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6132__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6683__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold690 hold690/A VGND VGND VPWR VPWR _7161_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6467__A _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4446__A1 _4446_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2080 _7424_/Q VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2091 hold314/X VGND VGND VPWR VPWR _4396_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1390 hold1414/X VGND VGND VPWR VPWR hold1415/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5946__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7066__RESET_B _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3972__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6371__A1 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6371__B2 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput206 _3405_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
XFILLER_114_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput217 _4165_/X VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ _3643_/Y _4300_/A1 _4302_/S VGND VGND VPWR VPWR _6985_/D sky130_fd_sc_hd__mux2_1
Xoutput228 _7665_/X VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput239 _4138_/X VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
XANTENNA__6123__A1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5280_ _4836_/A _5061_/B _5399_/C _5279_/Y VGND VGND VPWR VPWR _5280_/X sky130_fd_sc_hd__a31o_1
XFILLER_153_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4231_ _4258_/A0 _4422_/A1 _4231_/S VGND VGND VPWR VPWR _4231_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6674__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ _6939_/Q _4164_/A1 _7258_/Q VGND VGND VPWR VPWR _4162_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4093_ _4093_/A _4093_/B _4093_/C _4093_/D VGND VGND VPWR VPWR _4096_/C sky130_fd_sc_hd__and4_1
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4328__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6729__A3 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6803_ _4427_/C _6803_/A2 _6803_/B1 _4426_/Y _6802_/X VGND VGND VPWR VPWR _6803_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4995_ _4996_/A _5339_/A _5029_/A _5034_/B VGND VGND VPWR VPWR _5033_/C sky130_fd_sc_hd__nand4_1
XANTENNA__5401__A3 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6734_ _7054_/Q _6434_/B _6771_/A3 _6420_/C _7125_/Q VGND VGND VPWR VPWR _6734_/X
+ sky130_fd_sc_hd__a32o_1
X_3946_ _7295_/Q _5965_/B _3562_/C _3666_/X _7011_/Q VGND VGND VPWR VPWR _3946_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3877_ _7027_/Q _4352_/A _3514_/X _5668_/A _7288_/Q VGND VGND VPWR VPWR _3877_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3963__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6665_ _7001_/Q _6419_/D _6424_/X _7127_/Q _6664_/X VGND VGND VPWR VPWR _6665_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5616_ _5616_/A0 _5949_/A1 _5618_/S VGND VGND VPWR VPWR _5616_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5165__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6596_ _7284_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6596_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4373__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3715__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5547_ _4741_/Y _5065_/Y _5352_/Y _5448_/B _5546_/X VGND VGND VPWR VPWR _5575_/B
+ sky130_fd_sc_hd__o2111a_2
XFILLER_191_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7671__A _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5478_ _5478_/A _5478_/B _5559_/B VGND VGND VPWR VPWR _5478_/Y sky130_fd_sc_hd__nor3_1
XFILLER_172_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4125__A0 input84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7217_ _4150_/A1 _7217_/D _6869_/X VGND VGND VPWR VPWR _7217_/Q sky130_fd_sc_hd__dfrtn_1
XANTENNA__6665__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4429_ _4114_/B _4429_/B VGND VGND VPWR VPWR _4430_/D sky130_fd_sc_hd__nand2b_1
Xfanout400 _5965_/A VGND VGND VPWR VPWR _5992_/C sky130_fd_sc_hd__buf_4
XANTENNA__3479__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout411 _3484_/X VGND VGND VPWR VPWR _5695_/A sky130_fd_sc_hd__buf_8
Xfanout422 _4860_/Y VGND VGND VPWR VPWR _4924_/B sky130_fd_sc_hd__buf_6
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout444 _3860_/D VGND VGND VPWR VPWR _4551_/C sky130_fd_sc_hd__buf_4
X_7148_ _7561_/CLK _7148_/D fanout738/X VGND VGND VPWR VPWR _7148_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout455 _3682_/A VGND VGND VPWR VPWR _5590_/A sky130_fd_sc_hd__clkbuf_16
Xfanout466 _4861_/X VGND VGND VPWR VPWR _5038_/B sky130_fd_sc_hd__buf_4
Xfanout477 _6651_/B VGND VGND VPWR VPWR _6462_/C sky130_fd_sc_hd__clkbuf_8
X_7079_ _7095_/CLK _7079_/D fanout749/X VGND VGND VPWR VPWR _7659_/A sky130_fd_sc_hd__dfrtp_1
Xfanout488 _6116_/A VGND VGND VPWR VPWR _6097_/C sky130_fd_sc_hd__clkbuf_4
Xfanout499 _6136_/C VGND VGND VPWR VPWR _6270_/C1 sky130_fd_sc_hd__buf_4
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A wb_adr_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input74_A pad_flash_io1_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6105__A1 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6656__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3890__A2 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5919__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3800_ _7139_/Q _4479_/A _3576_/X _3798_/X VGND VGND VPWR VPWR _3800_/X sky130_fd_sc_hd__a31o_4
X_4780_ _5091_/C _5260_/C _5059_/B VGND VGND VPWR VPWR _4781_/A sky130_fd_sc_hd__and3_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A1 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _4177_/B _4231_/S _3727_/X _3729_/X _3730_/X VGND VGND VPWR VPWR _3732_/D
+ sky130_fd_sc_hd__a2111o_2
Xclkbuf_leaf_0_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7232_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2276_A _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4180__A _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3662_ _3931_/B _5640_/B _5596_/A VGND VGND VPWR VPWR _4394_/A sky130_fd_sc_hd__and3_4
X_6450_ _7559_/Q _6419_/C _6442_/X _6445_/X _6449_/X VGND VGND VPWR VPWR _6471_/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5147__A2 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6344__B2 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5001__D1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5401_ _4836_/A _5399_/A _5134_/A _5400_/Y VGND VGND VPWR VPWR _5401_/X sky130_fd_sc_hd__a31o_1
X_6381_ _6966_/Q _6144_/A _6144_/B _6332_/C _7035_/Q VGND VGND VPWR VPWR _6381_/X
+ sky130_fd_sc_hd__a32o_1
X_3593_ _7413_/Q _5803_/A _5731_/A _5713_/A _7333_/Q VGND VGND VPWR VPWR _3593_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2443_A _7414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5332_ _5183_/A _5011_/A _5339_/B _5331_/Y VGND VGND VPWR VPWR _5332_/X sky130_fd_sc_hd__a31o_1
XFILLER_126_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5263_ _5222_/A _5068_/B _5387_/D _4756_/X VGND VGND VPWR VPWR _5263_/X sky130_fd_sc_hd__a31o_1
XFILLER_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5855__A0 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2805 hold773/X VGND VGND VPWR VPWR _4193_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4214_ _4214_/A0 _5645_/A0 _4214_/S VGND VGND VPWR VPWR _4214_/X sky130_fd_sc_hd__mux2_1
X_7002_ _7210_/CLK _7002_/D fanout700/X VGND VGND VPWR VPWR _7002_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2816 hold991/X VGND VGND VPWR VPWR _4471_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2827 _7649_/A VGND VGND VPWR VPWR hold2827/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5194_ _5339_/A _5188_/X _5183_/B _5170_/X _5193_/X VGND VGND VPWR VPWR _5194_/Y
+ sky130_fd_sc_hd__a311oi_2
Xhold2838 _5705_/X VGND VGND VPWR VPWR _7319_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2849 _5687_/X VGND VGND VPWR VPWR _7303_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4145_ _7562_/Q _4174_/B _4144_/Y VGND VGND VPWR VPWR _4145_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3881__A2 _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ _6909_/Q _4076_/B _4076_/C _6910_/Q VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__and4b_1
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout359_A _3552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3633__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5386__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6583__A1 _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4978_ _5410_/A _5029_/A VGND VGND VPWR VPWR _4978_/Y sky130_fd_sc_hd__nand2_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6583__B2 _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6717_ _7159_/Q _6419_/A _6419_/C _7139_/Q _6716_/X VGND VGND VPWR VPWR _6717_/X
+ sky130_fd_sc_hd__a221o_1
X_3929_ _3929_/A VGND VGND VPWR VPWR _3929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3936__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_42_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6648_ wire351/X _6647_/Y _7286_/Q _6431_/Y VGND VGND VPWR VPWR _6648_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_166_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6335__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__C _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6579_ _7372_/Q _6413_/C _6651_/C _6058_/X _7532_/Q VGND VGND VPWR VPWR _6579_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6638__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3434__A _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6271__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4265__A _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3624__A2 _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5795__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5129__A2 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire642 _5071_/Y VGND VGND VPWR VPWR _5072_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_171_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap419 _6411_/Y VGND VGND VPWR VPWR _6431_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_136_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6629__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2024_A _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6262__B1 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4175__A _4175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5950_ _5950_/A0 _5950_/A1 _5955_/S VGND VGND VPWR VPWR _5950_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3615__A2 _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4901_ _4726_/Y _4899_/Y _4898_/Y _4894_/Y _4891_/Y VGND VGND VPWR VPWR _4902_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5881_ _5881_/A0 _5881_/A1 _5883_/S VGND VGND VPWR VPWR _5881_/X sky130_fd_sc_hd__mux2_1
X_7620_ _7625_/CLK _7620_/D fanout711/X VGND VGND VPWR VPWR _7620_/Q sky130_fd_sc_hd__dfrtp_1
X_4832_ _5260_/B _4836_/C VGND VGND VPWR VPWR _4832_/Y sky130_fd_sc_hd__nand2_8
XFILLER_33_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6565__A1 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6565__B2 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7551_ _7551_/CLK _7551_/D fanout734/X VGND VGND VPWR VPWR _7551_/Q sky130_fd_sc_hd__dfstp_1
X_4763_ _4763_/A _4763_/B _4763_/C VGND VGND VPWR VPWR _4763_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3918__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3519__A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6502_ _7401_/Q _6409_/X _6420_/B _7305_/Q _6499_/X VGND VGND VPWR VPWR _6502_/X
+ sky130_fd_sc_hd__a221o_1
X_3714_ _6966_/Q _4352_/B _4265_/B _3663_/X _7166_/Q VGND VGND VPWR VPWR _3714_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7482_ _7565_/CLK _7482_/D fanout743/X VGND VGND VPWR VPWR _7482_/Q sky130_fd_sc_hd__dfrtp_4
X_4694_ _4768_/B _4753_/C _4730_/C _4801_/C VGND VGND VPWR VPWR _4696_/B sky130_fd_sc_hd__nor4_4
XFILLER_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6433_ _6441_/D _7598_/Q _7597_/Q _6433_/D VGND VGND VPWR VPWR _6433_/X sky130_fd_sc_hd__and4bb_4
X_3645_ _3644_/X _3645_/A1 _3996_/A VGND VGND VPWR VPWR _3645_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6364_ _7212_/Q _6089_/X _6379_/B1 _7190_/Q _6363_/X VGND VGND VPWR VPWR _6364_/X
+ sky130_fd_sc_hd__a221o_1
X_3576_ _4509_/C _3576_/B _3576_/C VGND VGND VPWR VPWR _3576_/X sky130_fd_sc_hd__and3_4
XANTENNA__3551__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3303 _6498_/X VGND VGND VPWR VPWR _7616_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3551__B2 hold52/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5315_ _5038_/A _5410_/A _4823_/B _4809_/B _5160_/C VGND VGND VPWR VPWR _5317_/C
+ sky130_fd_sc_hd__a311o_1
Xhold3314 _7640_/Q VGND VGND VPWR VPWR _6810_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6295_ _7142_/Q _6121_/C _6116_/C _6121_/B VGND VGND VPWR VPWR _6295_/X sky130_fd_sc_hd__o211a_1
XFILLER_170_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3325 _7607_/Q VGND VGND VPWR VPWR _6260_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3336 _7208_/Q VGND VGND VPWR VPWR _5580_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3347 _6890_/Q VGND VGND VPWR VPWR _4098_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2602 _4267_/X VGND VGND VPWR VPWR hold974/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2613 _7121_/Q VGND VGND VPWR VPWR hold753/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3358 _6902_/Q VGND VGND VPWR VPWR _4039_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5246_ _4622_/Y _4726_/Y _4748_/Y _4947_/Y _5245_/X VGND VGND VPWR VPWR _5247_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2624 _7451_/Q VGND VGND VPWR VPWR hold711/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3369 _6882_/Q VGND VGND VPWR VPWR _3400_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__buf_8
XFILLER_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2635 _6970_/Q VGND VGND VPWR VPWR hold777/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1901 hold353/X VGND VGND VPWR VPWR _4269_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__buf_6
XANTENNA__4500__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__buf_4
Xhold2646 _7030_/Q VGND VGND VPWR VPWR hold759/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2657 hold893/X VGND VGND VPWR VPWR _5900_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5177_ _5203_/C _5183_/C _5216_/A VGND VGND VPWR VPWR _5177_/Y sky130_fd_sc_hd__o21ai_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1912 _6969_/Q VGND VGND VPWR VPWR hold345/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1923 _7299_/Q VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2668 hold739/X VGND VGND VPWR VPWR _4466_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2679 _4445_/X VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1934 _7362_/Q VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout476_A _6428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1945 _4518_/X VGND VGND VPWR VPWR hold404/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1956 _7346_/Q VGND VGND VPWR VPWR hold367/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4128_ _6896_/Q _4128_/B VGND VGND VPWR VPWR _4128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1967 _4355_/X VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1978 _7123_/Q VGND VGND VPWR VPWR hold461/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1989 _7138_/Q VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6253__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4059_ _6892_/Q _6891_/Q _4123_/B _4058_/Y VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__o211a_1
XFILLER_24_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3909__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3429__A _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1758_A _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4319__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6459__B _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3041_A _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6492__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input37_A mgmt_gpio_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3845__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4426__C _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3781__A1 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5507__C1 _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold508 hold508/A VGND VGND VPWR VPWR _6935_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3430_ _7402_/Q VGND VGND VPWR VPWR _3430_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3533__A1 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5100_ _5100_/A _5260_/B _5107_/C VGND VGND VPWR VPWR _5100_/X sky130_fd_sc_hd__and3_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6080_ _6080_/A _6136_/B _6116_/A VGND VGND VPWR VPWR _6080_/X sky130_fd_sc_hd__and3_4
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5031_/A _5031_/B _5031_/C VGND VGND VPWR VPWR _5033_/A sky130_fd_sc_hd__nor3_1
XANTENNA__6483__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1208 hold3265/X VGND VGND VPWR VPWR hold1208/X sky130_fd_sc_hd__clkdlybuf4s25_2
Xhold1219 hold2876/X VGND VGND VPWR VPWR _7482_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3836__A2 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6235__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3521__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6982_ _7000_/CLK _6982_/D VGND VGND VPWR VPWR _6982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5933_ _5978_/A0 _5933_/A1 _5937_/S VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6250__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7565_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ _5999_/A1 _5864_/A1 _5865_/S VGND VGND VPWR VPWR _5864_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__A1 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6538__B2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4549__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7603_ _7625_/CLK _7603_/D fanout705/X VGND VGND VPWR VPWR _7603_/Q sky130_fd_sc_hd__dfrtp_1
X_4815_ _5107_/C _5059_/B _5399_/C VGND VGND VPWR VPWR _4818_/A sky130_fd_sc_hd__and3_1
XANTENNA__4352__B _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5795_ _5894_/A0 _5795_/A1 _5802_/S VGND VGND VPWR VPWR _5795_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5210__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2942_A _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7534_ _7572_/CLK hold67/X fanout736/X VGND VGND VPWR VPWR _7534_/Q sky130_fd_sc_hd__dfrtp_4
X_4746_ _4755_/A _5138_/B _4746_/C _5005_/A VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nand4_2
XFILLER_147_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7465_ _7563_/CLK _7465_/D fanout739/X VGND VGND VPWR VPWR _7465_/Q sky130_fd_sc_hd__dfrtp_4
X_4677_ _5089_/B _4675_/Y _4673_/Y _4562_/Y VGND VGND VPWR VPWR _5012_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6416_ _6466_/B _6467_/A _6651_/B _6466_/A VGND VGND VPWR VPWR _6419_/B sky130_fd_sc_hd__and4bb_1
X_3628_ _7540_/Q _3590_/C _5947_/B _3544_/X _7420_/Q VGND VGND VPWR VPWR _3628_/X
+ sky130_fd_sc_hd__a32o_1
X_7396_ _7582_/CLK _7396_/D fanout718/X VGND VGND VPWR VPWR _7396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6347_ _7053_/Q _6087_/X _6344_/X _6346_/X VGND VGND VPWR VPWR _6347_/X sky130_fd_sc_hd__a211o_1
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3559_ _7542_/Q _5947_/A _5947_/B _3558_/X _7286_/Q VGND VGND VPWR VPWR _3559_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA_fanout593_A hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3100 _7463_/Q VGND VGND VPWR VPWR hold3100/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_1_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3111 _7152_/Q VGND VGND VPWR VPWR hold3111/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3122 _6874_/Q VGND VGND VPWR VPWR hold3122/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3133 hold3133/A VGND VGND VPWR VPWR _4456_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3144 hold3144/A VGND VGND VPWR VPWR _4371_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2410 _4327_/X VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6278_ _7374_/Q _6144_/C _6388_/A3 _6110_/X _7438_/Q VGND VGND VPWR VPWR _6278_/X
+ sky130_fd_sc_hd__a32o_1
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR _4562_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_103_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5277__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3155 hold3155/A VGND VGND VPWR VPWR _4534_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR _4089_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2421 hold771/X VGND VGND VPWR VPWR _5666_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6474__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3166 hold3166/A VGND VGND VPWR VPWR _5975_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR input128/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2432 hold901/X VGND VGND VPWR VPWR _5737_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5911__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3177 _6933_/Q VGND VGND VPWR VPWR hold3177/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR _6800_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout760_A _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5229_ _4600_/Y _5091_/C _5213_/B _4916_/B VGND VGND VPWR VPWR _5231_/B sky130_fd_sc_hd__a31o_1
Xhold3188 _7222_/Q VGND VGND VPWR VPWR hold3188/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2443 _7414_/Q VGND VGND VPWR VPWR hold715/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2454 _5728_/X VGND VGND VPWR VPWR hold958/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3827__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3199 hold3199/A VGND VGND VPWR VPWR _4266_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1720 _7528_/Q VGND VGND VPWR VPWR hold347/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2465 _5835_/X VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1731 _4433_/X VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2476 hold925/X VGND VGND VPWR VPWR _5782_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1742 _7400_/Q VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2487 hold907/X VGND VGND VPWR VPWR _4547_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1753 hold276/X VGND VGND VPWR VPWR _5681_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2498 _4333_/X VGND VGND VPWR VPWR hold736/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4527__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1764 _7578_/Q VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6226__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1775 hold374/X VGND VGND VPWR VPWR _7432_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1786 _5976_/X VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1797 _6907_/Q VGND VGND VPWR VPWR _3450_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6241__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6529__A1 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__B2 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_90 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__B2 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3256_A _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6465__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5821__B _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6480__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6217__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6768__A1 _7045_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4172__B _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4600_ _4843_/A _5073_/A VGND VGND VPWR VPWR _4600_/Y sky130_fd_sc_hd__nor2_8
X_5580_ _5580_/A1 _5580_/A2 _5579_/X _5577_/Y VGND VGND VPWR VPWR _7208_/D sky130_fd_sc_hd__a211o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3754__A1 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4531_ _4531_/A0 _5585_/A0 _4532_/S VGND VGND VPWR VPWR _4531_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3754__B2 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold305 hold305/A VGND VGND VPWR VPWR _7096_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2356_A _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7250_ _7250_/CLK _7250_/D fanout692/X VGND VGND VPWR VPWR _7250_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6299__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4462_ _4462_/A0 _5912_/A1 _4466_/S VGND VGND VPWR VPWR _4462_/X sky130_fd_sc_hd__mux2_1
Xhold327 hold327/A VGND VGND VPWR VPWR _7067_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold338 hold338/A VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6201_ _7451_/Q _6112_/B _6116_/A _6089_/X _7507_/Q VGND VGND VPWR VPWR _6201_/X
+ sky130_fd_sc_hd__a32o_1
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3516__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3413_ _7538_/Q VGND VGND VPWR VPWR _3413_/Y sky130_fd_sc_hd__inv_2
X_4393_ _5736_/A1 _4393_/A1 _4393_/S VGND VGND VPWR VPWR _4393_/X sky130_fd_sc_hd__mux2_1
X_7181_ _7181_/CLK _7181_/D fanout721/X VGND VGND VPWR VPWR _7181_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _7320_/Q _6082_/X _6094_/X _7504_/Q _6131_/X VGND VGND VPWR VPWR _6132_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4628__A _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6063_ _6932_/Q _6061_/X _6067_/A _4117_/B VGND VGND VPWR VPWR _6063_/X sky130_fd_sc_hd__a211o_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 hold3015/X VGND VGND VPWR VPWR hold3016/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3532__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1016 hold3019/X VGND VGND VPWR VPWR hold3020/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _5768_/X VGND VGND VPWR VPWR _7375_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5014_ _5328_/A _5328_/B _5339_/C _5018_/B VGND VGND VPWR VPWR _5014_/Y sky130_fd_sc_hd__nand4_2
Xhold1038 hold3104/X VGND VGND VPWR VPWR _7479_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1049 hold3098/X VGND VGND VPWR VPWR hold3099/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6208__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _7179_/CLK _6965_/D fanout698/X VGND VGND VPWR VPWR _6965_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5431__A1 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5916_ _5916_/A0 _5979_/A0 _5919_/S VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__mux2_1
X_6896_ _7075_/CLK _6896_/D _6846_/X VGND VGND VPWR VPWR _6896_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3993__A1 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3993__B2 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5847_ _5847_/A0 _5991_/A1 _5847_/S VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout606_A _3444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5778_ _5994_/A1 _5778_/A1 _5784_/S VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3745__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7517_ _7565_/CLK hold69/X fanout748/X VGND VGND VPWR VPWR _7517_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3745__B2 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4729_ _4772_/A _4802_/A _4733_/B _4733_/A VGND VGND VPWR VPWR _4834_/B sky130_fd_sc_hd__and4b_2
XFILLER_181_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4302__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1456_A _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7448_ _7531_/CLK _7448_/D fanout744/X VGND VGND VPWR VPWR _7448_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6695__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold850 hold850/A VGND VGND VPWR VPWR _7054_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7379_ _7475_/CLK _7379_/D fanout729/X VGND VGND VPWR VPWR _7379_/Q sky130_fd_sc_hd__dfrtp_4
Xhold861 hold861/A VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold872 hold872/A VGND VGND VPWR VPWR _7416_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold894 hold894/A VGND VGND VPWR VPWR _7493_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3442__A _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2240 _7292_/Q VGND VGND VPWR VPWR hold695/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2251 hold571/X VGND VGND VPWR VPWR _5601_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2262 _6961_/Q VGND VGND VPWR VPWR hold555/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2273 _7273_/Q VGND VGND VPWR VPWR hold693/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input139_A wb_dat_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2284 _5955_/X VGND VGND VPWR VPWR hold576/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1550 _4439_/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2295 _5800_/X VGND VGND VPWR VPWR hold790/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1561 hold156/X VGND VGND VPWR VPWR _5845_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1572 hold138/X VGND VGND VPWR VPWR _5918_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1583 _3463_/X VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1594 _5919_/X VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold3004_A _5650_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3984__B2 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3617__A _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5489__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6686__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6438__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6453__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5661__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6750_ wire350/X wire349/X _6960_/Q _6431_/Y VGND VGND VPWR VPWR _6750_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3962_ _6962_/Q _4352_/B _5659_/B _5794_/A _7399_/Q VGND VGND VPWR VPWR _3962_/X
+ sky130_fd_sc_hd__a32o_1
X_5701_ _5701_/A0 _5953_/A1 _5703_/S VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3975__B2 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6681_ _7118_/Q _6427_/X _6679_/X _6680_/X VGND VGND VPWR VPWR _6681_/X sky130_fd_sc_hd__a211o_1
XFILLER_148_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3893_ _7536_/Q _3590_/C _5947_/B _3565_/X _7464_/Q VGND VGND VPWR VPWR _3893_/X
+ sky130_fd_sc_hd__a32o_1
X_5632_ _5992_/C _5632_/B _5992_/D VGND VGND VPWR VPWR _5633_/S sky130_fd_sc_hd__and3_1
XFILLER_164_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3727__A1 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5563_ _5563_/A1 _4722_/Y _4741_/Y _5084_/C _5379_/X VGND VGND VPWR VPWR _5564_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3527__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7302_ _7334_/CLK _7302_/D fanout710/X VGND VGND VPWR VPWR _7302_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4514_ _4514_/A0 _5817_/A1 _4514_/S VGND VGND VPWR VPWR _4514_/X sky130_fd_sc_hd__mux2_1
Xhold102 hold102/A VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5494_ _4595_/Y _4601_/Y _5495_/C1 _4834_/Y _5494_/B2 VGND VGND VPWR VPWR _5496_/C
+ sky130_fd_sc_hd__o32a_1
Xhold113 hold113/A VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold124 _3485_/X VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold135 hold135/A VGND VGND VPWR VPWR _7494_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6677__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7233_ _7255_/CLK _7233_/D fanout689/X VGND VGND VPWR VPWR _7233_/Q sky130_fd_sc_hd__dfstp_4
X_4445_ _4445_/A0 _5853_/A0 _4448_/S VGND VGND VPWR VPWR _4445_/X sky130_fd_sc_hd__mux2_1
Xhold146 hold146/A VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold157 hold157/A VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold179 hold179/A VGND VGND VPWR VPWR _7326_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7164_ _7164_/CLK _7164_/D fanout699/X VGND VGND VPWR VPWR _7164_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout615 _7593_/Q VGND VGND VPWR VPWR _6429_/C sky130_fd_sc_hd__buf_8
X_4376_ _4455_/A _4376_/B _4388_/B _4533_/B VGND VGND VPWR VPWR _4381_/S sky130_fd_sc_hd__and4_4
Xfanout626 _7111_/Q VGND VGND VPWR VPWR _4427_/D sky130_fd_sc_hd__buf_8
Xfanout637 _6930_/Q VGND VGND VPWR VPWR _6009_/B sky130_fd_sc_hd__buf_6
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ _7447_/Q _6144_/A _6120_/B _6379_/B1 _7519_/Q VGND VGND VPWR VPWR _6115_/X
+ sky130_fd_sc_hd__a32o_1
Xfanout648 _4871_/X VGND VGND VPWR VPWR _4970_/C sky130_fd_sc_hd__buf_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7095_/CLK _7095_/D fanout749/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfrtp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ _7594_/Q _6019_/A _6929_/Q _6045_/Y VGND VGND VPWR VPWR _7594_/D sky130_fd_sc_hd__o31a_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6444__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout556_A _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4805__B _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ _7314_/CLK _6948_/D fanout711/X VGND VGND VPWR VPWR _7653_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3966__B2 _7327_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6879_ _4127_/A1 _6879_/D _6830_/X VGND VGND VPWR VPWR _6879_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_139_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3718__A1 _7030_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3718__B2 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6380__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3437__A _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6668__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6132__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4143__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold680 _4490_/X VGND VGND VPWR VPWR _7146_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6683__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold691 hold691/A VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6467__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5891__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_635 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_37_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2070 hold2070/A VGND VGND VPWR VPWR _5805_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2081 hold521/X VGND VGND VPWR VPWR _5823_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5798__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2092 _7390_/Q VGND VGND VPWR VPWR hold2092/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1380 _7099_/Q VGND VGND VPWR VPWR _4447_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1391 hold1416/X VGND VGND VPWR VPWR hold1417/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6199__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3957__A1 _7479_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3957__B2 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6371__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput207 _3441_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput218 _7656_/X VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
XANTENNA__6659__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput229 _7666_/X VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
XANTENNA__6123__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4230_ _4230_/A0 _4229_/X _4232_/S VGND VGND VPWR VPWR _4230_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4161_ _6940_/Q _4161_/A1 _7260_/Q VGND VGND VPWR VPWR _4161_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ _4563_/C _4563_/D _4562_/A _4562_/B VGND VGND VPWR VPWR _4095_/C sky130_fd_sc_hd__nor4_1
XFILLER_82_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4625__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ _4427_/D _6802_/A2 _6802_/B1 _4427_/B VGND VGND VPWR VPWR _6802_/X sky130_fd_sc_hd__a22o_1
XFILLER_90_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4994_ _5158_/A _5034_/B _5180_/A VGND VGND VPWR VPWR _5035_/B sky130_fd_sc_hd__and3_1
XANTENNA__3948__A1 _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6733_ _7180_/Q _6058_/X _6728_/X _6732_/X _6430_/X VGND VGND VPWR VPWR _6733_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_3945_ _7335_/Q _3531_/X _3667_/X _7021_/Q _3944_/X VGND VGND VPWR VPWR _3961_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6664_ _7593_/Q _7117_/Q _6408_/C _6663_/X VGND VGND VPWR VPWR _6664_/X sky130_fd_sc_hd__a31o_1
X_3876_ _6989_/Q _4346_/C _5623_/B _3875_/X VGND VGND VPWR VPWR _3879_/C sky130_fd_sc_hd__a31o_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5615_ _5615_/A0 _5894_/A0 _5618_/S VGND VGND VPWR VPWR _5615_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6595_ _7396_/Q _6420_/C _6588_/X _6590_/X _6594_/X VGND VGND VPWR VPWR _6595_/X
+ sky130_fd_sc_hd__a2111o_2
XFILLER_164_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5546_ _4741_/Y _4886_/Y _4891_/Y _4894_/Y VGND VGND VPWR VPWR _5546_/X sky130_fd_sc_hd__o211a_1
XFILLER_132_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5477_ _5134_/A _5282_/B _5524_/A3 _5105_/X _5395_/X VGND VGND VPWR VPWR _5559_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_145_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4125__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7216_ _4127_/A1 _7216_/D _6868_/X VGND VGND VPWR VPWR _7216_/Q sky130_fd_sc_hd__dfrtn_1
X_4428_ _7107_/Q _4428_/B VGND VGND VPWR VPWR _4428_/Y sky130_fd_sc_hd__nand2b_4
Xfanout401 _5614_/B VGND VGND VPWR VPWR _5965_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__3479__A3 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout412 _5785_/B VGND VGND VPWR VPWR _4431_/A sky130_fd_sc_hd__buf_8
Xclkbuf_2_3__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4169_/B2
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5873__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout434 hold90/X VGND VGND VPWR VPWR _5956_/B sky130_fd_sc_hd__clkbuf_16
X_7147_ _7561_/CLK _7147_/D fanout737/X VGND VGND VPWR VPWR _7147_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout445 _3489_/Y VGND VGND VPWR VPWR _3860_/D sky130_fd_sc_hd__buf_8
X_4359_ _4359_/A0 _5876_/A1 _4363_/S VGND VGND VPWR VPWR _4359_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout456 hold76/X VGND VGND VPWR VPWR _3682_/A sky130_fd_sc_hd__buf_12
Xfanout478 _6413_/C VGND VGND VPWR VPWR _6651_/B sky130_fd_sc_hd__buf_4
X_7078_ _7095_/CLK _7078_/D fanout748/X VGND VGND VPWR VPWR _7658_/A sky130_fd_sc_hd__dfrtp_1
Xfanout489 _6078_/X VGND VGND VPWR VPWR _6116_/A sky130_fd_sc_hd__buf_12
XFILLER_59_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5625__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6029_ _6027_/X _6028_/Y _6019_/A VGND VGND VPWR VPWR _6029_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3636__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3939__A1 _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4551__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6353__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input67_A mgmt_gpio_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6105__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5616__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3890__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6041__A1 _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ _7571_/Q _5983_/A _4479_/A _4422_/S input48/X VGND VGND VPWR VPWR _3730_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3661_ _5740_/A _4515_/B _4509_/C VGND VGND VPWR VPWR _3661_/X sky130_fd_sc_hd__and3_2
XANTENNA__4180__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5001__C1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4355__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5400_ _5397_/X _5482_/A _5481_/B VGND VGND VPWR VPWR _5400_/Y sky130_fd_sc_hd__nand3b_1
X_6380_ _7005_/Q _6097_/B _6097_/C _6379_/X VGND VGND VPWR VPWR _6380_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3508__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3592_ _7437_/Q _3525_/X _3590_/X _3591_/X _3589_/X VGND VGND VPWR VPWR _3592_/X
+ sky130_fd_sc_hd__a2111o_1
X_5331_ _5495_/C1 _4759_/Y _5007_/Y _4690_/Y _5184_/X VGND VGND VPWR VPWR _5331_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5262_ _5563_/A1 _4737_/Y _5255_/X _5077_/Y _5480_/B2 VGND VGND VPWR VPWR _5564_/A
+ sky130_fd_sc_hd__o32a_1
X_7001_ _7164_/CLK _7001_/D fanout692/X VGND VGND VPWR VPWR _7001_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2806 _7266_/Q VGND VGND VPWR VPWR hold947/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4213_ _4213_/A0 _5948_/A1 _4214_/S VGND VGND VPWR VPWR _4213_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2817 _4471_/X VGND VGND VPWR VPWR hold992/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2828 hold2828/A VGND VGND VPWR VPWR _4239_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5193_ _5339_/A _5053_/C _5188_/X _5192_/X _5171_/X VGND VGND VPWR VPWR _5193_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_96_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2839 _7417_/Q VGND VGND VPWR VPWR hold2839/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3866__B1 _3549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4144_ _4144_/A _4174_/B VGND VGND VPWR VPWR _4144_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__6835__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5607__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3881__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4075_ hold196/A _4076_/B _4075_/S VGND VGND VPWR VPWR _6883_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3618__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_4_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__3633__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4977_ _5138_/A _5138_/B _5029_/A VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__and3_2
XANTENNA__6583__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6716_ _7053_/Q _6434_/B _6574_/C _6466_/X _7211_/Q VGND VGND VPWR VPWR _6716_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout421_A _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3928_ _6897_/Q _6882_/Q _7248_/Q VGND VGND VPWR VPWR _3929_/A sky130_fd_sc_hd__nor3_4
XFILLER_149_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6647_ _6647_/A _6647_/B _6647_/C _6647_/D VGND VGND VPWR VPWR _6647_/Y sky130_fd_sc_hd__nor4_4
XANTENNA__6335__A2 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3859_ _3859_/A _5992_/A _3860_/D _5992_/C VGND VGND VPWR VPWR _3859_/X sky130_fd_sc_hd__and4_2
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6578_ _7388_/Q _6413_/C _6426_/X _6577_/X VGND VGND VPWR VPWR _6578_/X sky130_fd_sc_hd__a31o_1
XFILLER_119_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4897__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3554__C1 _3551_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5529_ _5529_/A _5529_/B _5529_/C _5529_/D VGND VGND VPWR VPWR _5533_/A sky130_fd_sc_hd__and4_1
XFILLER_106_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6638__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5846__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4129__A_N _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input121_A wb_adr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4265__B _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A3 _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_csclk_A _4169_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5377__A3 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5782__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4281__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5096__B _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6326__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire654 _5282_/D VGND VGND VPWR VPWR _5115_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3560__A2 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5298__C1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3848__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4175__B input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4900_ _4601_/Y _4622_/Y _4726_/Y _4895_/Y _4896_/Y VGND VGND VPWR VPWR _4902_/A
+ sky130_fd_sc_hd__o311a_1
XTAP_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5880_ _5880_/A0 _5997_/A1 _5883_/S VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4831_ _4831_/A _4860_/A _4831_/C _4805_/B VGND VGND VPWR VPWR _4831_/Y sky130_fd_sc_hd__nor4b_2
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6565__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4191__A _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6892__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7550_ _7556_/CLK hold61/X fanout732/X VGND VGND VPWR VPWR _7550_/Q sky130_fd_sc_hd__dfrtp_2
X_4762_ _4772_/A _4801_/B _4803_/A _5404_/B VGND VGND VPWR VPWR _4763_/B sky130_fd_sc_hd__and4b_1
XANTENNA_clkbuf_leaf_6_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6501_ _7529_/Q _6058_/X _6422_/X _7289_/Q _6500_/X VGND VGND VPWR VPWR _6501_/X
+ sky130_fd_sc_hd__a221o_1
X_3713_ _7291_/Q hold90/A _5731_/B input30/X _3503_/X VGND VGND VPWR VPWR _3713_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3519__B _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7481_ _7563_/CLK _7481_/D fanout739/X VGND VGND VPWR VPWR _7481_/Q sky130_fd_sc_hd__dfrtp_4
X_4693_ _4733_/A _4733_/B _4801_/C VGND VGND VPWR VPWR _4794_/A sky130_fd_sc_hd__a21oi_4
X_6432_ _7527_/Q _6058_/X _6424_/X _7567_/Q VGND VGND VPWR VPWR _6432_/X sky130_fd_sc_hd__a22o_1
X_3644_ _7218_/Q _3643_/Y _3923_/S VGND VGND VPWR VPWR _3644_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6363_ _7054_/Q _6121_/A _6097_/C _6317_/C _7049_/Q VGND VGND VPWR VPWR _6363_/X
+ sky130_fd_sc_hd__a32o_1
X_3575_ input27/X _3488_/X _3490_/X input18/X _3574_/X VGND VGND VPWR VPWR _3575_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3535__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2818_A _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5314_ _5314_/A _5535_/A VGND VGND VPWR VPWR _5317_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5453__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3304 _7613_/Q VGND VGND VPWR VPWR _6400_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6294_ _7016_/Q _6086_/X _6121_/C _6988_/Q _6121_/X VGND VGND VPWR VPWR _6294_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3315 _7638_/Q VGND VGND VPWR VPWR _6804_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3326 _7074_/Q VGND VGND VPWR VPWR hold3326/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_170_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3337 _6880_/Q VGND VGND VPWR VPWR _4121_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2603 _7055_/Q VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5245_ _4571_/Y _4843_/A _4888_/C _4960_/A VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__o22a_1
Xhold3348 _4066_/Y VGND VGND VPWR VPWR _6891_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2614 hold753/X VGND VGND VPWR VPWR _4460_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3359 _6909_/Q VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2625 hold711/X VGND VGND VPWR VPWR _5853_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2636 hold777/X VGND VGND VPWR VPWR _4275_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1902 _4269_/X VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2647 hold759/X VGND VGND VPWR VPWR _4357_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2658 _5900_/X VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5176_ _5495_/C1 _4690_/Y _4971_/X _5014_/Y _5175_/X VGND VGND VPWR VPWR _5176_/X
+ sky130_fd_sc_hd__o311a_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1913 hold345/X VGND VGND VPWR VPWR _4274_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1924 hold212/X VGND VGND VPWR VPWR _5682_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2669 _4466_/X VGND VGND VPWR VPWR hold740/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1935 hold371/X VGND VGND VPWR VPWR _5753_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1946 _7323_/Q VGND VGND VPWR VPWR hold302/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4127_ input83/X _4127_/A1 _6896_/Q VGND VGND VPWR VPWR _4127_/X sky130_fd_sc_hd__mux2_1
Xhold1957 hold367/X VGND VGND VPWR VPWR _5735_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1968 _7307_/Q VGND VGND VPWR VPWR hold278/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6253__B2 _7509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1979 hold461/X VGND VGND VPWR VPWR _4463_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4058_ _4058_/A _4058_/B _7073_/Q VGND VGND VPWR VPWR _4058_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5896__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_5_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_5_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6556__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5764__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold214_A _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6308__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3790__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6459__C _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input169_A wb_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3845__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6244__A1 _7525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4723__B _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output290_A _6924_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3781__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold509 hold509/A VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6180__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3533__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__A1 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5030_ _5038_/A _5034_/B _5030_/C VGND VGND VPWR VPWR _5031_/B sky130_fd_sc_hd__and3_1
XANTENNA__6483__B2 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1209 hold1209/A VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_78_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3521__C _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ _7000_/CLK _6981_/D VGND VGND VPWR VPWR _6981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5932_ _5986_/A1 _5932_/A1 _5937_/S VGND VGND VPWR VPWR _5932_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5863_ _5998_/A1 _5863_/A1 _5865_/S VGND VGND VPWR VPWR _5863_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2670_A _7045_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7602_ _7625_/CLK _7602_/D fanout705/X VGND VGND VPWR VPWR _7602_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4125__S _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ _4831_/C _5260_/B _4814_/C VGND VGND VPWR VPWR _4814_/Y sky130_fd_sc_hd__nand3_4
XFILLER_166_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5794_ _5794_/A _5893_/B VGND VGND VPWR VPWR _5802_/S sky130_fd_sc_hd__nand2_8
XANTENNA__4352__C _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7533_ _7580_/CLK _7533_/D fanout733/X VGND VGND VPWR VPWR _7533_/Q sky130_fd_sc_hd__dfrtp_4
X_4745_ _5100_/A _5079_/B _5061_/B VGND VGND VPWR VPWR _4746_/C sky130_fd_sc_hd__and3_1
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7464_ _7562_/CLK _7464_/D fanout739/X VGND VGND VPWR VPWR _7464_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_190_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4676_ _4675_/A _4675_/B _4675_/C _4674_/A VGND VGND VPWR VPWR _4679_/A sky130_fd_sc_hd__a31o_2
XFILLER_119_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6415_ _6427_/A _6467_/A _6468_/C VGND VGND VPWR VPWR _6419_/A sky130_fd_sc_hd__and3_4
X_3627_ _7340_/Q _3531_/X _3532_/X input57/X _3626_/X VGND VGND VPWR VPWR _3632_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6171__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7395_ _7395_/CLK _7395_/D fanout737/X VGND VGND VPWR VPWR _7395_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6710__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6346_ _7008_/Q _6082_/X _6097_/X _7184_/Q _6345_/X VGND VGND VPWR VPWR _6346_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5183__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3558_ _5590_/A _5640_/B _5659_/B VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__and3_4
Xhold3101 hold3101/A VGND VGND VPWR VPWR _5867_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3112 hold3112/A VGND VGND VPWR VPWR _4498_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3123 hold3123/A VGND VGND VPWR VPWR _4182_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3134 _4456_/X VGND VGND VPWR VPWR hold3134/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6277_ _7422_/Q _6072_/X _6097_/X _7446_/Q _6276_/X VGND VGND VPWR VPWR _6280_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3145 _4371_/X VGND VGND VPWR VPWR hold3145/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout586_A hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3489_ _3507_/A _3576_/C VGND VGND VPWR VPWR _3489_/Y sky130_fd_sc_hd__nor2_4
Xhold2400 hold867/X VGND VGND VPWR VPWR _4390_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR _4562_/A sky130_fd_sc_hd__clkbuf_2
Xhold2411 _7316_/Q VGND VGND VPWR VPWR hold903/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3156 _7046_/Q VGND VGND VPWR VPWR hold3156/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR input118/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2422 _5666_/X VGND VGND VPWR VPWR hold772/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6474__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5277__A2 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3167 _5975_/X VGND VGND VPWR VPWR hold3167/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5228_ _5228_/A _5228_/B _5228_/C _5228_/D VGND VGND VPWR VPWR _5231_/A sky130_fd_sc_hd__nand4_1
XANTENNA__6474__B2 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR _4564_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3178 hold3178/A VGND VGND VPWR VPWR _4218_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2433 _7483_/Q VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3189 hold3189/A VGND VGND VPWR VPWR _5588_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2444 hold715/X VGND VGND VPWR VPWR _5811_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4808__B _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1710 _5892_/X VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2455 hold958/X VGND VGND VPWR VPWR _7340_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3827__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1721 hold347/X VGND VGND VPWR VPWR _5940_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2466 _7114_/Q VGND VGND VPWR VPWR hold861/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1732 _6914_/Q VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2477 _5782_/X VGND VGND VPWR VPWR hold926/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1743 hold391/X VGND VGND VPWR VPWR _5796_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5159_ _5410_/A _4706_/A _5453_/B _5158_/X VGND VGND VPWR VPWR _5160_/D sky130_fd_sc_hd__a31o_1
XANTENNA_fanout753_A input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2488 _4547_/X VGND VGND VPWR VPWR hold908/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1754 _5681_/X VGND VGND VPWR VPWR hold277/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2499 _7505_/Q VGND VGND VPWR VPWR hold863/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1765 hold154/X VGND VGND VPWR VPWR _5996_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1776 _7670_/A VGND VGND VPWR VPWR hold282/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1787 _7376_/Q VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1798 _3450_/X VGND VGND VPWR VPWR _3451_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6631__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6529__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5201__A2 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3763__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _6304_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6465__A1 _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5821__C hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6768__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4734__A _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output303_A _3578_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5976__A0 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4530_ _4530_/A0 _4548_/A0 _4532_/S VGND VGND VPWR VPWR _4530_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3754__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6153__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4461_ _4473_/A _4551_/A _4551_/C _4533_/B VGND VGND VPWR VPWR _4466_/S sky130_fd_sc_hd__and4_4
Xhold317 hold317/A VGND VGND VPWR VPWR _7090_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold328 hold328/A VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6099__C _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6200_ _7467_/Q _6121_/A _6116_/A _6317_/C _7515_/Q VGND VGND VPWR VPWR _6200_/X
+ sky130_fd_sc_hd__a32o_1
Xhold339 hold339/A VGND VGND VPWR VPWR _7048_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3412_ _7546_/Q VGND VGND VPWR VPWR _3412_/Y sky130_fd_sc_hd__inv_2
X_7180_ _7180_/CLK _7180_/D fanout728/X VGND VGND VPWR VPWR _7180_/Q sky130_fd_sc_hd__dfrtp_4
X_4392_ _5647_/A0 _4392_/A1 _4393_/S VGND VGND VPWR VPWR _4392_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _7408_/Q _6144_/C _6097_/B _6270_/C1 VGND VGND VPWR VPWR _6131_/X sky130_fd_sc_hd__o211a_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__A1 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6009_/Y _6019_/Y _6061_/X _6932_/Q VGND VGND VPWR VPWR _6062_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5731__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 _5984_/X VGND VGND VPWR VPWR _7567_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1017 hold3021/X VGND VGND VPWR VPWR _7455_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__B _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5013_ _5158_/A _5339_/A _5013_/C VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__and3_2
Xhold1028 hold3079/X VGND VGND VPWR VPWR hold3080/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1039 hold3044/X VGND VGND VPWR VPWR hold3045/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3690__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6759__A2 _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ _7179_/CLK _6964_/D fanout698/X VGND VGND VPWR VPWR _6964_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5915_ _5915_/A0 _5978_/A0 _5919_/S VGND VGND VPWR VPWR _5915_/X sky130_fd_sc_hd__mux2_1
X_6895_ _4127_/A1 _6895_/D _6845_/X VGND VGND VPWR VPWR _6895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5719__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5846_ _5846_/A0 _5990_/A1 _5847_/S VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6392__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5777_ _5993_/A1 _5777_/A1 _5784_/S VGND VGND VPWR VPWR _5777_/X sky130_fd_sc_hd__mux2_1
X_4728_ _5260_/C _5387_/D _5059_/B VGND VGND VPWR VPWR _4763_/A sky130_fd_sc_hd__and3_1
XANTENNA_fanout501_A _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3745__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7516_ _7565_/CLK _7516_/D fanout746/X VGND VGND VPWR VPWR _7516_/Q sky130_fd_sc_hd__dfrtp_4
X_7447_ _7561_/CLK _7447_/D fanout738/X VGND VGND VPWR VPWR _7447_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_162_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4659_ _5248_/A _5248_/B VGND VGND VPWR VPWR _4659_/Y sky130_fd_sc_hd__nand2_4
XFILLER_135_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6695__A1 _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold840 hold840/A VGND VGND VPWR VPWR _7449_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7378_ _7575_/CLK _7378_/D fanout734/X VGND VGND VPWR VPWR _7378_/Q sky130_fd_sc_hd__dfrtp_4
Xhold851 hold851/A VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold862 hold862/A VGND VGND VPWR VPWR _7114_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold873 hold873/A VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold884 hold884/A VGND VGND VPWR VPWR _6989_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6329_ _6958_/Q _6036_/Y _6067_/A VGND VGND VPWR VPWR _6329_/X sky130_fd_sc_hd__o21a_1
Xhold895 hold895/A VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2230 _7302_/Q VGND VGND VPWR VPWR hold569/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2241 hold695/X VGND VGND VPWR VPWR _5674_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2252 _7537_/Q VGND VGND VPWR VPWR hold629/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2263 hold555/X VGND VGND VPWR VPWR _4264_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2274 hold693/X VGND VGND VPWR VPWR _5653_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2285 _7476_/Q VGND VGND VPWR VPWR hold767/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1540 _5935_/X VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2296 _7370_/Q VGND VGND VPWR VPWR hold615/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1551 _6955_/Q VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1562 _5845_/X VGND VGND VPWR VPWR hold157/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1573 _5918_/X VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1584 hold88/X VGND VGND VPWR VPWR _3504_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1595 _7529_/Q VGND VGND VPWR VPWR hold206/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3984__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input97_A usr2_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3617__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6135__B1 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6150__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7522_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6438__A1 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7491_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ _3961_/A _3961_/B _3961_/C _3961_/D VGND VGND VPWR VPWR _3995_/B sky130_fd_sc_hd__nor4_1
XFILLER_189_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5994__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5700_ _5700_/A0 _5952_/A1 _5703_/S VGND VGND VPWR VPWR _5700_/X sky130_fd_sc_hd__mux2_1
X_6680_ _7052_/Q _6434_/B _6771_/A3 _6463_/X _7163_/Q VGND VGND VPWR VPWR _6680_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3892_ _7360_/Q _5803_/A _5965_/B _3891_/X VGND VGND VPWR VPWR _3892_/X sky130_fd_sc_hd__a31o_1
X_5631_ _5640_/D _5631_/B VGND VGND VPWR VPWR _5631_/X sky130_fd_sc_hd__and2_1
XFILLER_188_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5295__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2466_A _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3727__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5562_ _5393_/X _5478_/B _5562_/C _5562_/D VGND VGND VPWR VPWR _5562_/Y sky130_fd_sc_hd__nand4bb_1
X_7301_ _7334_/CLK _7301_/D fanout710/X VGND VGND VPWR VPWR _7301_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3527__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4513_ _4513_/A0 _5585_/A0 _4514_/S VGND VGND VPWR VPWR _4513_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6126__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 hold103/A VGND VGND VPWR VPWR hold103/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5493_ _4595_/Y _4832_/Y _5528_/A3 _5492_/X VGND VGND VPWR VPWR _5493_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_144_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold114 _7227_/Q VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold125 _3598_/B VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7232_ _7232_/CLK _7232_/D _4128_/B VGND VGND VPWR VPWR _7232_/Q sky130_fd_sc_hd__dfrtp_4
X_4444_ _4444_/A0 _5996_/A1 _4448_/S VGND VGND VPWR VPWR _4444_/X sky130_fd_sc_hd__mux2_1
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold147 hold147/A VGND VGND VPWR VPWR _7318_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6838__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6141__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold169 hold169/A VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7163_ _7212_/CLK _7163_/D fanout723/X VGND VGND VPWR VPWR _7163_/Q sky130_fd_sc_hd__dfrtp_4
X_4375_ _5853_/A0 _4375_/A1 _4375_/S VGND VGND VPWR VPWR _4375_/X sky130_fd_sc_hd__mux2_1
Xfanout605 _3444_/Y VGND VGND VPWR VPWR _6121_/C sky130_fd_sc_hd__buf_6
XANTENNA__3543__A _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout616 _7592_/Q VGND VGND VPWR VPWR _6332_/B sky130_fd_sc_hd__buf_6
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6114_ _7383_/Q _6109_/X _6110_/X _7431_/Q _6113_/X VGND VGND VPWR VPWR _6114_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout627 _7110_/Q VGND VGND VPWR VPWR _4427_/C sky130_fd_sc_hd__buf_8
Xfanout638 _6751_/S VGND VGND VPWR VPWR _6649_/S sky130_fd_sc_hd__buf_6
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7094_ _7095_/CLK _7094_/D fanout749/X VGND VGND VPWR VPWR _7094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6434_/B _6466_/C _6019_/A VGND VGND VPWR VPWR _6045_/Y sky130_fd_sc_hd__o21ai_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__A1 _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6854__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_A _4446_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__A1 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__B2 _7525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4093__B _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6947_ _7306_/CLK _6947_/D _4079_/A VGND VGND VPWR VPWR _6947_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4612__B1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3966__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6878_ _7201_/CLK _6878_/D fanout726/X VGND VGND VPWR VPWR _6878_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4821__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5829_ _5829_/A0 hold20/X hold33/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__mux2_1
XFILLER_139_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3718__A2 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4143__A2 _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold670 hold670/A VGND VGND VPWR VPWR _7136_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold681 hold681/A VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold692 hold692/A VGND VGND VPWR VPWR _7045_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1900_A _6965_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input151_A wb_dat_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2060 _7395_/Q VGND VGND VPWR VPWR hold389/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2071 _5805_/X VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2082 _7368_/Q VGND VGND VPWR VPWR hold515/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2093 hold2093/A VGND VGND VPWR VPWR _5784_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1370 _6792_/A1 VGND VGND VPWR VPWR hold3029/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1381 hold1441/X VGND VGND VPWR VPWR hold1442/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input12_A mask_rev_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1392 hold2092/X VGND VGND VPWR VPWR hold2093/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3957__A2 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6356__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4223__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6371__A3 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput208 _3440_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XANTENNA__6659__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput219 _7657_/X VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5331__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _7282_/Q input1/X _4159_/Y VGND VGND VPWR VPWR _4160_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__4178__B _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3893__B2 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4091_ _4562_/C _4562_/D _4091_/C input116/X VGND VGND VPWR VPWR _4093_/D sky130_fd_sc_hd__nor4b_1
XFILLER_56_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4625__C _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6801_ _6800_/X hold485/A _6822_/S VGND VGND VPWR VPWR _7637_/D sky130_fd_sc_hd__mux2_1
XFILLER_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5398__A1 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4993_ _5203_/C _5034_/B _5180_/A VGND VGND VPWR VPWR _5035_/A sky130_fd_sc_hd__and3_1
XFILLER_90_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_700 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3944_ _6897_/Q _6882_/Q _7248_/Q _5619_/A _5619_/B VGND VGND VPWR VPWR _3944_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__3948__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6732_ _7130_/Q _6424_/X _6730_/X _6731_/X VGND VGND VPWR VPWR _6732_/X sky130_fd_sc_hd__a211o_1
X_6663_ _7172_/Q _6747_/B _6747_/C _6408_/A _7147_/Q VGND VGND VPWR VPWR _6663_/X
+ sky130_fd_sc_hd__a32o_1
X_3875_ _6928_/Q hold90/A _5640_/C _3861_/X VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__a31o_1
XFILLER_149_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3538__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4133__S _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5614_ _5731_/A _5614_/B _5947_/C VGND VGND VPWR VPWR _5614_/X sky130_fd_sc_hd__and3_2
XFILLER_176_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6594_ _7516_/Q _6435_/X _6591_/X _6593_/X VGND VGND VPWR VPWR _6594_/X sky130_fd_sc_hd__a211o_1
XFILLER_164_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5545_ _5545_/A _5545_/B _5545_/C _5545_/D VGND VGND VPWR VPWR _5548_/B sky130_fd_sc_hd__nor4_1
XFILLER_191_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3581__B1 _3549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_0_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_5476_ _5476_/A _5476_/B _5476_/C VGND VGND VPWR VPWR _5478_/B sky130_fd_sc_hd__nand3_1
X_4427_ _7107_/Q _4427_/B _4427_/C _4427_/D VGND VGND VPWR VPWR _4430_/C sky130_fd_sc_hd__nor4_4
X_7215_ _4127_/A1 _7215_/D _6867_/X VGND VGND VPWR VPWR _7215_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_132_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout499_A _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout402 hold1802/X VGND VGND VPWR VPWR _5614_/B sky130_fd_sc_hd__buf_12
Xfanout413 _3933_/A VGND VGND VPWR VPWR _5785_/B sky130_fd_sc_hd__buf_6
X_7146_ _7213_/CLK _7146_/D fanout700/X VGND VGND VPWR VPWR _7146_/Q sky130_fd_sc_hd__dfrtp_4
X_4358_ _4473_/A _4551_/C _4509_/C _4533_/B VGND VGND VPWR VPWR _4363_/S sky130_fd_sc_hd__and4_4
XFILLER_160_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout435 hold89/X VGND VGND VPWR VPWR hold90/A sky130_fd_sc_hd__buf_8
XANTENNA__3884__A1 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5899__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout446 _5830_/C VGND VGND VPWR VPWR _4455_/A sky130_fd_sc_hd__buf_6
XANTENNA_input4_A mask_rev_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout457 _5612_/A VGND VGND VPWR VPWR _4551_/A sky130_fd_sc_hd__buf_12
XFILLER_171_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7077_ _7095_/CLK _7077_/D fanout748/X VGND VGND VPWR VPWR _7657_/A sky130_fd_sc_hd__dfrtp_1
Xfanout479 _6561_/A2 VGND VGND VPWR VPWR _6413_/C sky130_fd_sc_hd__buf_6
XFILLER_101_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4289_ _3570_/Y _4289_/A1 _4289_/S VGND VGND VPWR VPWR _6979_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6028_ _7589_/Q _7588_/Q _6081_/C VGND VGND VPWR VPWR _6028_/Y sky130_fd_sc_hd__nor3_1
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3636__A1 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3636__B2 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4816__B _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4551__B _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7139__SET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6105__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3627__B2 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6577__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6041__A2 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6329__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4461__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3660_ _4455_/A _3860_/D _5614_/B VGND VGND VPWR VPWR _4467_/A sky130_fd_sc_hd__and3_4
XANTENNA__4180__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6344__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5552__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3591_ input59/X _3933_/A _5614_/B _5704_/A _7325_/Q VGND VGND VPWR VPWR _3591_/X
+ sky130_fd_sc_hd__a32o_1
X_5330_ _5495_/C1 _4759_/Y _5007_/Y _4690_/Y _5173_/X VGND VGND VPWR VPWR _5554_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5261_ _5480_/B2 _4727_/Y _5516_/A3 _5077_/Y _5260_/Y VGND VGND VPWR VPWR _5265_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5304__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6501__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7000_ _7000_/CLK _7000_/D VGND VGND VPWR VPWR _7000_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ hold90/X _5640_/C _5640_/D VGND VGND VPWR VPWR _4214_/S sky130_fd_sc_hd__and3_1
Xhold2807 hold947/X VGND VGND VPWR VPWR _5645_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5192_ _5034_/C _5188_/X _5190_/X _5191_/X VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__a211o_1
Xhold2818 _6989_/Q VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2829 _4239_/X VGND VGND VPWR VPWR hold2829/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4143_ _7570_/Q _4142_/A _4142_/Y VGND VGND VPWR VPWR _4143_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA_clkbuf_leaf_2_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4074_ hold4/A hold196/A _4074_/S VGND VGND VPWR VPWR _6884_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3618__B2 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5083__A3 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6568__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _4956_/A _4956_/B _4975_/X _4826_/Y VGND VGND VPWR VPWR _5438_/B sky130_fd_sc_hd__a211o_1
XANTENNA__5240__B1 wire649/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6583__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6715_ _6969_/Q _6420_/A _6704_/X _6714_/X VGND VGND VPWR VPWR _6715_/X sky130_fd_sc_hd__a211o_1
X_3927_ _7263_/Q _5640_/A _5640_/B _5640_/C VGND VGND VPWR VPWR _3927_/X sky130_fd_sc_hd__and4_2
XANTENNA__5791__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3858_ _3858_/A1 _3996_/A _3856_/Y _3857_/X VGND VGND VPWR VPWR _7216_/D sky130_fd_sc_hd__a22o_1
X_6646_ _7462_/Q _6455_/X _6645_/X _6644_/X _6643_/X VGND VGND VPWR VPWR _6647_/D
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__6335__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6577_ _7484_/Q _6447_/C _6459_/C _6421_/X _7324_/Q VGND VGND VPWR VPWR _6577_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6740__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3789_ _7346_/Q _3590_/C _4352_/A _3525_/X _7434_/Q VGND VGND VPWR VPWR _3789_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3554__B1 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4897__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5528_ _4595_/Y _4832_/Y _5528_/A3 _5422_/D _5294_/A VGND VGND VPWR VPWR _5529_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5459_ _5222_/A _5134_/A _5248_/A _5458_/X VGND VGND VPWR VPWR _5459_/X sky130_fd_sc_hd__a31o_1
XFILLER_133_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7129_ _7395_/CLK _7129_/D fanout737/X VGND VGND VPWR VPWR _7129_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4827__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_15__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X VGND VGND VPWR VPWR _7646_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4265__C _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input114_A wb_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6559__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3279_A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire655 _4831_/Y VGND VGND VPWR VPWR _5282_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_7_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6731__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3848__A1 _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4737__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6262__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4273__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4830_ _4830_/A _4830_/B _4830_/C VGND VGND VPWR VPWR _4837_/A sky130_fd_sc_hd__nor3_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4903__C _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4761_ _4831_/C _4801_/B _5404_/B VGND VGND VPWR VPWR _4761_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__4191__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5773__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6500_ _7369_/Q _6651_/B _6651_/C _6457_/X _7473_/Q VGND VGND VPWR VPWR _6500_/X
+ sky130_fd_sc_hd__a32o_1
X_3712_ _7515_/Q _5920_/A _3704_/X _3706_/X _3711_/X VGND VGND VPWR VPWR _3732_/B
+ sky130_fd_sc_hd__a2111o_2
X_7480_ _7531_/CLK _7480_/D fanout739/X VGND VGND VPWR VPWR _7480_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3519__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4692_ _5038_/A _5328_/A _5328_/B VGND VGND VPWR VPWR _4692_/Y sky130_fd_sc_hd__nand3_4
XFILLER_146_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_6_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6431_ _6431_/A _6431_/B _6431_/C VGND VGND VPWR VPWR _6431_/Y sky130_fd_sc_hd__nand3_4
X_3643_ _3643_/A _3643_/B _3643_/C VGND VGND VPWR VPWR _3643_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6722__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4411__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3536__B1 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6362_ _6357_/X _6362_/B _6362_/C VGND VGND VPWR VPWR _6362_/Y sky130_fd_sc_hd__nand3b_4
X_3574_ _7573_/Q _3872_/A2 _5965_/A _5974_/A _7565_/Q VGND VGND VPWR VPWR _3574_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_161_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3535__B _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5313_ _4723_/Y _4796_/Y _4978_/Y _4793_/Y _5312_/X VGND VGND VPWR VPWR _5535_/A
+ sky130_fd_sc_hd__o221a_1
X_6293_ _7021_/Q _6070_/X _6087_/X _7051_/Q _6292_/X VGND VGND VPWR VPWR _6293_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3551__A3 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3305 _7625_/Q VGND VGND VPWR VPWR _6751_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3316 _7600_/Q VGND VGND VPWR VPWR _6064_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3327 _7604_/Q VGND VGND VPWR VPWR _6170_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5244_ _5367_/B _5545_/A _5244_/C VGND VGND VPWR VPWR _5247_/B sky130_fd_sc_hd__nor3_1
Xhold3338 _6899_/Q VGND VGND VPWR VPWR _4047_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3349 _7583_/Q VGND VGND VPWR VPWR _6002_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2604 hold657/X VGND VGND VPWR VPWR _4387_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3839__A1 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2615 _4460_/X VGND VGND VPWR VPWR hold754/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3839__B2 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2626 _5853_/X VGND VGND VPWR VPWR hold712/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5175_ _4956_/B _5174_/Y _5012_/Y VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__a21o_1
Xhold2637 _4275_/X VGND VGND VPWR VPWR hold778/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1903 _7314_/Q VGND VGND VPWR VPWR hold318/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2648 _4357_/X VGND VGND VPWR VPWR hold760/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2659 _7015_/Q VGND VGND VPWR VPWR hold729/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1914 _4274_/X VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1925 _7274_/Q VGND VGND VPWR VPWR hold377/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1936 _5753_/X VGND VGND VPWR VPWR hold372/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4126_ _6897_/Q _4128_/B VGND VGND VPWR VPWR _4126_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1947 hold302/X VGND VGND VPWR VPWR _5709_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1958 _5735_/X VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1969 hold278/X VGND VGND VPWR VPWR _5691_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4057_ _4057_/A0 _4076_/B _4057_/S VGND VGND VPWR VPWR _6893_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4264__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout531_A _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4382__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6556__A3 _6428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4813__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4959_ _5248_/A _5248_/B _5453_/C _4953_/X _5113_/A VGND VGND VPWR VPWR _4959_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3775__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6308__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6629_ _7542_/Q _6408_/D _6435_/X hold52/A VGND VGND VPWR VPWR _6629_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3790__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4321__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6492__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4255__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3766__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3781__A3 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4231__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6180__A1 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6180__B2 _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3533__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__A2 _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4494__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5691__A0 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5997__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6235__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4246__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6980_ _7000_/CLK _6980_/D VGND VGND VPWR VPWR _6980_/Q sky130_fd_sc_hd__dfxtp_1
X_5931_ _5976_/A0 _5931_/A1 _5937_/S VGND VGND VPWR VPWR _5931_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4914__B _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5994__A1 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5862_ _5997_/A1 _5862_/A1 _5865_/S VGND VGND VPWR VPWR _5862_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6538__A3 _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7601_ _7601_/CLK _7601_/D _6873_/A VGND VGND VPWR VPWR _7601_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5746__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4813_ _4984_/B _5260_/B _4814_/C VGND VGND VPWR VPWR _4983_/C sky130_fd_sc_hd__and3_2
X_5793_ _5793_/A0 hold20/X hold48/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__mux2_1
XANTENNA__3757__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5210__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7532_ _7574_/CLK _7532_/D fanout730/X VGND VGND VPWR VPWR _7532_/Q sky130_fd_sc_hd__dfrtp_4
X_4744_ _5282_/A _5282_/B VGND VGND VPWR VPWR _4744_/Y sky130_fd_sc_hd__nand2_4
XFILLER_147_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4675_ _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4675_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__7200__RESET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7463_ _7562_/CLK _7463_/D fanout739/X VGND VGND VPWR VPWR _7463_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3509__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6414_ _6466_/A _6466_/B _6463_/A _6462_/C VGND VGND VPWR VPWR _6420_/C sky130_fd_sc_hd__and4_4
X_3626_ _7428_/Q hold32/A _5965_/B _5704_/A _7324_/Q VGND VGND VPWR VPWR _3626_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_134_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6171__A1 _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6171__B2 _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7394_ _7578_/CLK _7394_/D fanout747/X VGND VGND VPWR VPWR _7394_/Q sky130_fd_sc_hd__dfrtp_4
X_6345_ _7048_/Q _6332_/B _6317_/C _6110_/X _7174_/Q VGND VGND VPWR VPWR _6345_/X
+ sky130_fd_sc_hd__a32o_1
X_3557_ _3511_/C hold46/X _3557_/C VGND VGND VPWR VPWR _3557_/X sky130_fd_sc_hd__and3b_2
Xhold3102 _7479_/Q VGND VGND VPWR VPWR hold3102/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3113 _7172_/Q VGND VGND VPWR VPWR hold3113/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6276_ _7494_/Q _6080_/A _6276_/A3 _6119_/X _7406_/Q VGND VGND VPWR VPWR _6276_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3124 _4182_/X VGND VGND VPWR VPWR hold3124/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3135 _7122_/Q VGND VGND VPWR VPWR hold3135/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3488_ _5640_/A _4328_/A _5612_/B VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__and3_4
Xhold2401 _4390_/X VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3146 _7471_/Q VGND VGND VPWR VPWR hold3146/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR _4562_/D sky130_fd_sc_hd__clkbuf_2
Xhold2412 hold903/X VGND VGND VPWR VPWR _5701_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3157 hold3157/A VGND VGND VPWR VPWR _4377_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5227_ _4775_/C _4885_/X _4907_/X VGND VGND VPWR VPWR _5228_/D sky130_fd_sc_hd__a21oi_2
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR input119/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3168 _7127_/Q VGND VGND VPWR VPWR hold3168/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2423 _7261_/Q VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3179 _4218_/X VGND VGND VPWR VPWR hold3179/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2434 hold625/X VGND VGND VPWR VPWR _5889_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1700 hold190/X VGND VGND VPWR VPWR _4434_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2445 _5811_/X VGND VGND VPWR VPWR hold716/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout579_A _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1711 _7301_/Q VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2456 _7043_/Q VGND VGND VPWR VPWR hold829/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1722 _5940_/X VGND VGND VPWR VPWR hold348/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5158_ _5158_/A _5158_/B _5410_/A VGND VGND VPWR VPWR _5158_/X sky130_fd_sc_hd__and3_1
Xhold2467 hold861/X VGND VGND VPWR VPWR _4452_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1733 hold152/X VGND VGND VPWR VPWR _4195_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2478 _7070_/Q VGND VGND VPWR VPWR hold749/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2489 _7366_/Q VGND VGND VPWR VPWR hold713/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1744 _5796_/X VGND VGND VPWR VPWR hold392/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1755 _7512_/Q VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6226__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4109_ _4427_/B _4084_/X _4425_/A VGND VGND VPWR VPWR _7109_/D sky130_fd_sc_hd__a21o_1
Xhold1766 _5996_/X VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1777 hold282/X VGND VGND VPWR VPWR _5646_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5089_ _5091_/C _5089_/B _5089_/C _5089_/D VGND VGND VPWR VPWR _5089_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__5700__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1788 hold349/X VGND VGND VPWR VPWR _5769_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1799 _3451_/Y VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5985__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3748__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_70 _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _7068_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6162__A1 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input42_A mgmt_gpio_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6465__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6882__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5673__A0 _5673_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4476__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2990 _6949_/Q VGND VGND VPWR VPWR hold2990/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5425__B1 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5728__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7215__CLK_N _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4460_ _4460_/A0 _5853_/A0 _4460_/S VGND VGND VPWR VPWR _4460_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold307 hold307/A VGND VGND VPWR VPWR _7484_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold318 hold318/A VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3411_ _7554_/Q VGND VGND VPWR VPWR _3411_/Y sky130_fd_sc_hd__inv_2
Xhold329 hold329/A VGND VGND VPWR VPWR _7007_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4391_ _4548_/A0 _4391_/A1 _4391_/S VGND VGND VPWR VPWR _4391_/X sky130_fd_sc_hd__mux2_1
X_6130_ _7472_/Q _6032_/Y _6276_/A3 _7488_/Q _6129_/X VGND VGND VPWR VPWR _6130_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_124_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4909__B _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6061_ _7585_/Q _7584_/Q _7586_/Q _7587_/Q VGND VGND VPWR VPWR _6061_/X sky130_fd_sc_hd__a211o_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6456__A2 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2411_A _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5012_/A _5328_/B _5013_/C VGND VGND VPWR VPWR _5012_/Y sky130_fd_sc_hd__nand3_2
Xhold1007 hold3006/X VGND VGND VPWR VPWR hold3007/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3532__C _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1018 hold3085/X VGND VGND VPWR VPWR hold3086/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1029 hold3081/X VGND VGND VPWR VPWR _7511_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4219__A1 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3690__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6759__A3 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5967__A1 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ _7180_/CLK _6963_/D fanout721/X VGND VGND VPWR VPWR _6963_/Q sky130_fd_sc_hd__dfrtp_4
X_5914_ _5914_/A0 _5914_/A1 _5919_/S VGND VGND VPWR VPWR _5914_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6894_ _4127_/A1 _6894_/D _6844_/X VGND VGND VPWR VPWR _6894_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5845_ _5845_/A0 _5998_/A1 _5847_/S VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3993__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ _5776_/A _5956_/C VGND VGND VPWR VPWR _5784_/S sky130_fd_sc_hd__nand2_8
XFILLER_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7515_ _7531_/CLK _7515_/D fanout740/X VGND VGND VPWR VPWR _7515_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4727_ _5260_/C _5387_/D VGND VGND VPWR VPWR _4727_/Y sky130_fd_sc_hd__nand2_2
XFILLER_135_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7446_ _7525_/CLK _7446_/D fanout745/X VGND VGND VPWR VPWR _7446_/Q sky130_fd_sc_hd__dfrtp_4
X_4658_ _4954_/A _5248_/A _5213_/A VGND VGND VPWR VPWR _4952_/B sky130_fd_sc_hd__and3_2
XFILLER_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR _4142_/B sky130_fd_sc_hd__clkbuf_4
Xhold830 hold830/A VGND VGND VPWR VPWR _7043_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3609_ _3608_/X _3609_/A1 _3996_/A VGND VGND VPWR VPWR _7220_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6695__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7377_ _7528_/CLK _7377_/D fanout729/X VGND VGND VPWR VPWR _7377_/Q sky130_fd_sc_hd__dfrtp_4
X_4589_ _4825_/A _4674_/A VGND VGND VPWR VPWR _5115_/B sky130_fd_sc_hd__and2b_4
XANTENNA_fanout696_A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold852 hold852/A VGND VGND VPWR VPWR _7029_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold863 hold863/A VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6328_ _6312_/X _6314_/X _6327_/Y VGND VGND VPWR VPWR _6328_/X sky130_fd_sc_hd__a21bo_4
Xhold874 hold874/A VGND VGND VPWR VPWR _6876_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold885 hold885/A VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold896 hold896/A VGND VGND VPWR VPWR _7405_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4819__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2220 _4308_/X VGND VGND VPWR VPWR hold538/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6259_ _7285_/Q _6036_/Y _6623_/B1 VGND VGND VPWR VPWR _6259_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4458__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5655__A0 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2231 hold569/X VGND VGND VPWR VPWR _5685_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2242 _5674_/X VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2253 hold629/X VGND VGND VPWR VPWR _5950_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2264 _7297_/Q VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1530 _7436_/Q VGND VGND VPWR VPWR hold192/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2275 _5653_/X VGND VGND VPWR VPWR hold694/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2286 hold767/X VGND VGND VPWR VPWR _5881_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1541 _7445_/Q VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2297 hold615/X VGND VGND VPWR VPWR _5762_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1552 hold85/X VGND VGND VPWR VPWR _4257_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1563 hold157/X VGND VGND VPWR VPWR _7444_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1574 _7024_/Q VGND VGND VPWR VPWR hold93/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3681__A2 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1585 _3504_/Y VGND VGND VPWR VPWR hold1585/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5407__B1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1596 hold206/X VGND VGND VPWR VPWR _5941_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5958__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4630__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4570__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5186__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3617__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6686__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5894__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6438__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5646__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4745__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5949__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6610__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3960_ _7122_/Q _3665_/X _3952_/X _3954_/X _3959_/X VGND VGND VPWR VPWR _3961_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_189_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3891_ _7193_/Q _4545_/A _3669_/X _6968_/Q _3890_/X VGND VGND VPWR VPWR _3891_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_189_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5630_ _5630_/A0 _5732_/A1 _5630_/S VGND VGND VPWR VPWR _5630_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5177__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4911__C _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _5561_/A1 _4814_/Y _5471_/X _5278_/B VGND VGND VPWR VPWR _5562_/D sky130_fd_sc_hd__o31a_1
XFILLER_163_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7300_ _7334_/CLK _7300_/D fanout710/X VGND VGND VPWR VPWR _7300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4512_ _4512_/A0 _4548_/A0 _4514_/S VGND VGND VPWR VPWR _4512_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6126__A1 _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3527__C _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5492_ _5486_/Y _5488_/Y _5532_/B _5492_/D VGND VGND VPWR VPWR _5492_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__6126__B2 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold104 _3505_/C VGND VGND VPWR VPWR _3504_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold115 hold115/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7231_ _7232_/CLK _7231_/D fanout689/X VGND VGND VPWR VPWR _7231_/Q sky130_fd_sc_hd__dfrtp_4
Xhold126 _4207_/S VGND VGND VPWR VPWR _4211_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6677__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4443_ hold7/X _5635_/A0 _4448_/S VGND VGND VPWR VPWR _4443_/X sky130_fd_sc_hd__mux2_1
Xhold137 hold137/A VGND VGND VPWR VPWR _7525_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold148 hold148/A VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold159 hold159/A VGND VGND VPWR VPWR _7569_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7162_ _7211_/CLK _7162_/D fanout700/X VGND VGND VPWR VPWR _7162_/Q sky130_fd_sc_hd__dfrtp_4
X_4374_ _4555_/A0 _4374_/A1 _4375_/S VGND VGND VPWR VPWR _4374_/X sky130_fd_sc_hd__mux2_1
Xfanout606 _3444_/Y VGND VGND VPWR VPWR _6119_/D sky130_fd_sc_hd__buf_6
XFILLER_113_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3543__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout617 _7592_/Q VGND VGND VPWR VPWR _6112_/C sky130_fd_sc_hd__buf_6
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6113_ _7367_/Q _6082_/C _6388_/A3 _6112_/X _7479_/Q VGND VGND VPWR VPWR _6113_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 _7109_/Q VGND VGND VPWR VPWR _4427_/B sky130_fd_sc_hd__buf_12
X_7093_ _7095_/CLK _7093_/D fanout747/X VGND VGND VPWR VPWR _7093_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout639 _6930_/Q VGND VGND VPWR VPWR _6751_/S sky130_fd_sc_hd__clkbuf_4
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5637__A0 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4358__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _7594_/Q _6429_/C VGND VGND VPWR VPWR _6443_/B sky130_fd_sc_hd__and2b_2
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6601__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6946_ _7581_/CLK _6946_/D fanout715/X VGND VGND VPWR VPWR _7652_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__6870__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_A _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4612__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3966__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6877_ _7201_/CLK _6877_/D fanout725/X VGND VGND VPWR VPWR _6877_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5828_ _5828_/A0 _5999_/A1 hold33/X VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout709_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4821__C _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3718__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5759_ _5993_/A1 _5759_/A1 hold27/X VGND VGND VPWR VPWR _5759_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6117__B2 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7429_ _7581_/CLK _7429_/D fanout716/X VGND VGND VPWR VPWR _7429_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold660 _5648_/X VGND VGND VPWR VPWR _7269_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold671 hold671/A VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold682 hold682/A VGND VGND VPWR VPWR _7418_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold693 hold693/A VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input144_A wb_dat_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2050 _4469_/X VGND VGND VPWR VPWR hold472/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4300__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2061 hold389/X VGND VGND VPWR VPWR _5790_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2072 _7133_/Q VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2083 hold515/X VGND VGND VPWR VPWR _5760_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_92_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2094 _5784_/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1360 _4312_/A1 VGND VGND VPWR VPWR hold3010/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1371 _6791_/A1 VGND VGND VPWR VPWR hold3036/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1382 hold1443/X VGND VGND VPWR VPWR hold1444/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1393 hold2160/X VGND VGND VPWR VPWR hold2161/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5800__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput209 _3439_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XANTENNA__6659__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5331__A2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3893__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4090_ _4564_/C _4564_/D _4563_/A _4563_/B VGND VGND VPWR VPWR _4095_/B sky130_fd_sc_hd__nor4_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6292__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4906__C _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6800_ _4427_/B _6800_/A2 _6800_/B1 _4426_/Y _6799_/X VGND VGND VPWR VPWR _6800_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5398__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4992_ _5038_/A _5183_/A _5038_/B _5053_/C VGND VGND VPWR VPWR _4992_/Y sky130_fd_sc_hd__nand4_1
XFILLER_90_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6731_ _7004_/Q _6419_/D _6446_/X _7190_/Q VGND VGND VPWR VPWR _6731_/X sky130_fd_sc_hd__a22o_1
X_3943_ input71/X _4231_/S _3934_/X _3935_/X _3942_/X VGND VGND VPWR VPWR _3961_/A
+ sky130_fd_sc_hd__a2111o_4
XANTENNA__4831__D_N _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4414__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6662_ _6874_/Q _6600_/B _6459_/C _6661_/X VGND VGND VPWR VPWR _6662_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3874_ _7280_/Q _5731_/A _5659_/B _3598_/X VGND VGND VPWR VPWR _3879_/B sky130_fd_sc_hd__a31o_4
XFILLER_176_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5613_ _5613_/A0 _5894_/A0 _5613_/S VGND VGND VPWR VPWR _5613_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3538__B _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6593_ _7548_/Q _6419_/A _6419_/C _7564_/Q _6592_/X VGND VGND VPWR VPWR _6593_/X
+ sky130_fd_sc_hd__a221o_1
X_5544_ _5453_/C _5180_/B _5248_/B _5453_/A VGND VGND VPWR VPWR _5545_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3581__B2 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ _4722_/Y _4748_/Y _4806_/Y _5561_/A1 VGND VGND VPWR VPWR _5476_/C sky130_fd_sc_hd__a211o_1
XFILLER_160_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5858__A0 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7214_ _4150_/A1 _7214_/D _6866_/X VGND VGND VPWR VPWR _7214_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_105_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4426_ _4427_/B _4427_/C _4427_/D VGND VGND VPWR VPWR _4426_/Y sky130_fd_sc_hd__nor3_4
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout403 _3590_/C VGND VGND VPWR VPWR _5947_/A sky130_fd_sc_hd__buf_8
X_7145_ _7191_/CLK _7145_/D fanout700/X VGND VGND VPWR VPWR _7145_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout414 _3472_/X VGND VGND VPWR VPWR _3933_/A sky130_fd_sc_hd__buf_8
XFILLER_99_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4357_ _4357_/A0 _5817_/A1 _4357_/S VGND VGND VPWR VPWR _4357_/X sky130_fd_sc_hd__mux2_1
Xfanout436 _4491_/C VGND VGND VPWR VPWR _5596_/B sky130_fd_sc_hd__buf_12
XANTENNA__3884__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout447 _3483_/X VGND VGND VPWR VPWR _5830_/C sky130_fd_sc_hd__buf_6
Xfanout458 _5612_/A VGND VGND VPWR VPWR _5992_/A sky130_fd_sc_hd__buf_6
X_7076_ _7095_/CLK _7076_/D fanout748/X VGND VGND VPWR VPWR _7656_/A sky130_fd_sc_hd__dfrtp_1
X_4288_ _3607_/Y _4288_/A1 _4289_/S VGND VGND VPWR VPWR _6978_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_4_14__f_wb_clk_i clkbuf_3_7_0_wb_clk_i/X VGND VGND VPWR VPWR _7641_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6283__B1 _6281_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6027_ _7589_/Q _7588_/Q _6081_/C VGND VGND VPWR VPWR _6027_/X sky130_fd_sc_hd__o21a_1
XFILLER_100_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout561_A _5726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3636__A2 _3486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7587_/CLK _6929_/D _6873_/A VGND VGND VPWR VPWR _6929_/Q sky130_fd_sc_hd__dfstp_4
Xclkbuf_leaf_31_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7514_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3939__A3 _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_46_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7435_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5561__A2 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3572__A1 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold490 hold490/A VGND VGND VPWR VPWR _6939_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3875__A2 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6274__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3627__A2 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 _4206_/X VGND VGND VPWR VPWR _6921_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4234__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4180__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3590_ _7477_/Q hold32/A _3590_/C VGND VGND VPWR VPWR _3590_/X sky130_fd_sc_hd__and3_1
XANTENNA__5552__A2 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5260_ _5260_/A _5260_/B _5260_/C _5260_/D VGND VGND VPWR VPWR _5260_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__5304__A2 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6501__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6501__B2 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4211_ _4211_/A0 _5955_/A1 _4211_/S VGND VGND VPWR VPWR _4211_/X sky130_fd_sc_hd__mux2_1
X_5191_ _4924_/B _5180_/A _5180_/B _5035_/C VGND VGND VPWR VPWR _5191_/X sky130_fd_sc_hd__a31o_1
Xhold2808 _7185_/Q VGND VGND VPWR VPWR hold993/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2819 hold883/X VGND VGND VPWR VPWR _4305_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3866__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4142_ _4142_/A _4142_/B VGND VGND VPWR VPWR _4142_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6265__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4073_ hold12/A hold4/A _4074_/S VGND VGND VPWR VPWR _6885_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4409__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3618__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6568__B2 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4975_ _4984_/B _4984_/A _4660_/Y _4672_/X VGND VGND VPWR VPWR _4975_/X sky130_fd_sc_hd__a211o_1
XANTENNA_hold2860_A _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3549__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6714_ _6990_/Q _6420_/B _6706_/X _6710_/X _6713_/X VGND VGND VPWR VPWR _6714_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_149_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3926_ _6874_/Q hold31/A _3514_/X _3494_/X _7471_/Q VGND VGND VPWR VPWR _3926_/X
+ sky130_fd_sc_hd__a32o_1
X_6645_ _7438_/Q _6747_/B _6747_/C VGND VGND VPWR VPWR _6645_/X sky130_fd_sc_hd__and3_1
X_3857_ _3924_/A1 _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3857_/X sky130_fd_sc_hd__o211a_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_A _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6576_ _7380_/Q _6408_/B _6423_/X _7332_/Q _6575_/X VGND VGND VPWR VPWR _6576_/X
+ sky130_fd_sc_hd__a221o_1
X_3788_ _7170_/Q _3647_/X _4340_/A _7019_/Q _3787_/X VGND VGND VPWR VPWR _3788_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3554__A1 _4176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4751__B1 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__B2 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5527_ hold29/A _5580_/A2 _5560_/B _5526_/X _5515_/X VGND VGND VPWR VPWR _7206_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5458_ _5134_/A _5248_/A _5089_/D _5252_/B VGND VGND VPWR VPWR _5458_/X sky130_fd_sc_hd__a31o_1
XFILLER_105_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4409_ _4409_/A0 _4408_/X _4423_/S VGND VGND VPWR VPWR _4409_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout776_A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5389_ _4601_/Y _4700_/Y _4844_/Y _4789_/Y VGND VGND VPWR VPWR _5518_/C sky130_fd_sc_hd__a31o_1
XANTENNA__5703__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7128_ _7395_/CLK _7128_/D fanout737/X VGND VGND VPWR VPWR _7128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4319__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ _7191_/CLK _7059_/D fanout701/X VGND VGND VPWR VPWR _7059_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4795__A_N _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6271__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__A1 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__B2 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input107_A wb_adr_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input72_A mgmt_gpio_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3848__A2 _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6247__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4229__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5470__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _5139_/D _4760_/B _4760_/C _4760_/D VGND VGND VPWR VPWR _4763_/C sky130_fd_sc_hd__nand4_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4191__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3784__A1 _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3711_ input24/X _3488_/X _3707_/X _3708_/X _3710_/X VGND VGND VPWR VPWR _3711_/X
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__3784__B2 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4691_ _5038_/A _5012_/A _5328_/B VGND VGND VPWR VPWR _5297_/A sky130_fd_sc_hd__and3_2
XFILLER_174_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_24_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6430_ _6431_/A _6431_/B _6431_/C VGND VGND VPWR VPWR _6430_/X sky130_fd_sc_hd__and3_4
XFILLER_146_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3642_ _3642_/A _3642_/B _3642_/C _3642_/D VGND VGND VPWR VPWR _3642_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__6722__A1 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5525__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6722__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6361_ _7039_/Q _6111_/X _6121_/X _6991_/Q _6360_/X VGND VGND VPWR VPWR _6362_/C
+ sky130_fd_sc_hd__a221oi_4
X_3573_ _3572_/X _3573_/A1 _3996_/A VGND VGND VPWR VPWR _7221_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7477__RESET_B fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5312_ _4667_/A _4692_/Y _4768_/Y _4796_/Y _4755_/Y VGND VGND VPWR VPWR _5312_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3535__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6292_ _7197_/Q _6332_/B _6079_/X _6094_/X _7209_/Q VGND VGND VPWR VPWR _6292_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_154_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3306 _7617_/Q VGND VGND VPWR VPWR _6523_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6486__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3317 _7602_/Q VGND VGND VPWR VPWR _6124_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3328 _7615_/Q VGND VGND VPWR VPWR _6473_/B2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5243_ _5248_/B _5453_/A _5243_/C VGND VGND VPWR VPWR _5367_/B sky130_fd_sc_hd__and3_1
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3339 _6905_/Q VGND VGND VPWR VPWR _4023_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2605 _4387_/X VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2616 _7577_/Q VGND VGND VPWR VPWR hold929/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2627 _7181_/Q VGND VGND VPWR VPWR hold721/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__buf_4
X_5174_ _4888_/C _5011_/B _5183_/C VGND VGND VPWR VPWR _5174_/Y sky130_fd_sc_hd__a21oi_4
Xhold2638 _7116_/Q VGND VGND VPWR VPWR hold705/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1904 hold318/X VGND VGND VPWR VPWR _5699_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2649 _7165_/Q VGND VGND VPWR VPWR hold825/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1915 _7363_/Q VGND VGND VPWR VPWR hold284/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4139__S _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1926 hold377/X VGND VGND VPWR VPWR _5654_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4125_ input84/X _4168_/D _6897_/Q VGND VGND VPWR VPWR _4125_/X sky130_fd_sc_hd__mux2_2
XFILLER_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1937 _7422_/Q VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6789__A1 _6789_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1948 _5709_/X VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1959 _7318_/Q VGND VGND VPWR VPWR hold146/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6253__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4056_ _6910_/Q _6909_/Q _6908_/Q _7071_/Q VGND VGND VPWR VPWR _4057_/S sky130_fd_sc_hd__and4bb_1
XFILLER_36_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4382__B _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _4958_/A _4958_/B _4958_/C VGND VGND VPWR VPWR _4962_/A sky130_fd_sc_hd__nand3_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3775__A1 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3775__B2 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3909_ _6963_/Q _4352_/B _4265_/B _5794_/A _7400_/Q VGND VGND VPWR VPWR _3909_/X
+ sky130_fd_sc_hd__a32o_1
X_4889_ _4889_/A _4889_/B VGND VGND VPWR VPWR _4891_/D sky130_fd_sc_hd__nor2_1
XFILLER_165_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6628_ _7310_/Q _6420_/B _6463_/X _7430_/Q _6627_/X VGND VGND VPWR VPWR _6628_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6559_ _7323_/Q _6421_/X _6462_/X _7363_/Q _6558_/X VGND VGND VPWR VPWR _6559_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_hold1541_A _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6477__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4557__B _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3766__A1 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_832 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6704__A1 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6180__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__A _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6483__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4467__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5443__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6640__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5930_ _5975_/A0 _5930_/A1 _5937_/S VGND VGND VPWR VPWR _7519_/D sky130_fd_sc_hd__mux2_1
XFILLER_46_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ _5978_/A0 _5861_/A1 _5865_/S VGND VGND VPWR VPWR _5861_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7600_ _7601_/CLK _7600_/D fanout692/X VGND VGND VPWR VPWR _7600_/Q sky130_fd_sc_hd__dfrtp_1
X_4812_ _4812_/A _4812_/B _4812_/C VGND VGND VPWR VPWR _4818_/C sky130_fd_sc_hd__nand3_1
X_5792_ _5792_/A0 _5999_/A1 hold48/X VGND VGND VPWR VPWR _5792_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7531_ _7531_/CLK _7531_/D fanout741/X VGND VGND VPWR VPWR _7531_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_159_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3757__B2 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4743_ _4910_/D _4856_/A _5073_/B VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__nor3_2
XFILLER_187_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4422__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7462_ _7556_/CLK hold63/X fanout731/X VGND VGND VPWR VPWR _7462_/Q sky130_fd_sc_hd__dfrtp_2
X_4674_ _4674_/A _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4679_/C sky130_fd_sc_hd__nand4_4
XFILLER_119_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6413_ _6434_/B _6468_/C _6413_/C VGND VGND VPWR VPWR _6420_/B sky130_fd_sc_hd__and3_4
X_3625_ _7460_/Q _5857_/A hold77/A _7524_/Q _3624_/X VGND VGND VPWR VPWR _3632_/A
+ sky130_fd_sc_hd__a221o_1
X_7393_ _7395_/CLK _7393_/D fanout737/X VGND VGND VPWR VPWR _7393_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6171__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4182__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6344_ _7038_/Q _6121_/C _6388_/A3 _6112_/X _6876_/Q VGND VGND VPWR VPWR _6344_/X
+ sky130_fd_sc_hd__a32o_1
X_3556_ _5612_/A _5640_/A _3562_/C VGND VGND VPWR VPWR _5704_/A sky130_fd_sc_hd__and3_4
Xhold3103 hold3103/A VGND VGND VPWR VPWR _5885_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_170_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6275_ _7470_/Q _6087_/X _6094_/X _7510_/Q _6274_/X VGND VGND VPWR VPWR _6280_/B
+ sky130_fd_sc_hd__a221o_1
Xhold3114 hold3114/A VGND VGND VPWR VPWR _4522_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3125 _7147_/Q VGND VGND VPWR VPWR hold3125/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3487_ _7406_/Q _5794_/A _3486_/X input10/X _3479_/X VGND VGND VPWR VPWR _3487_/X
+ sky130_fd_sc_hd__a221o_1
Xhold3136 hold3136/A VGND VGND VPWR VPWR _4462_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3562__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2402 _7161_/Q VGND VGND VPWR VPWR hold689/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3147 hold3147/A VGND VGND VPWR VPWR _5876_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR _4562_/C sky130_fd_sc_hd__clkbuf_2
Xhold2413 _5701_/X VGND VGND VPWR VPWR hold904/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3158 _4377_/X VGND VGND VPWR VPWR hold3158/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5226_ _4933_/B _4907_/B _4918_/D _5102_/B wire658/X VGND VGND VPWR VPWR _5226_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5131__B1 _5028_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6474__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3169 hold3169/A VGND VGND VPWR VPWR _4468_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2424 hold701/X VGND VGND VPWR VPWR _5638_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2435 _5889_/X VGND VGND VPWR VPWR hold626/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5682__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1701 _4434_/X VGND VGND VPWR VPWR hold191/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2446 _7191_/Q VGND VGND VPWR VPWR hold663/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2457 hold829/X VGND VGND VPWR VPWR _4373_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1712 hold182/X VGND VGND VPWR VPWR _5684_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5157_ _5107_/C _5059_/B _5453_/B _4977_/X _4823_/B VGND VGND VPWR VPWR _5160_/C
+ sky130_fd_sc_hd__a32o_1
Xhold1723 _7484_/Q VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2468 _4452_/X VGND VGND VPWR VPWR hold862/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1734 _4195_/X VGND VGND VPWR VPWR hold153/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2479 hold749/X VGND VGND VPWR VPWR _4405_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1745 _7004_/Q VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1756 hold415/X VGND VGND VPWR VPWR _5922_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4108_ _6009_/B _6427_/A _4105_/B _4107_/Y _4100_/X VGND VGND VPWR VPWR _6932_/D
+ sky130_fd_sc_hd__a41o_1
Xhold1767 hold155/X VGND VGND VPWR VPWR _7578_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1778 _5646_/X VGND VGND VPWR VPWR hold283/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5088_ _4600_/Y _5086_/B _5087_/Y VGND VGND VPWR VPWR _5088_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1789 _5769_/X VGND VGND VPWR VPWR hold350/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4039_ _4039_/A0 _4038_/X _4040_/A VGND VGND VPWR VPWR _6902_/D sky130_fd_sc_hd__mux2_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1589_A _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3748__A1 _7354_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4840__B _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__A _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_60 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_82 _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_93 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1923_A _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3920__A1 _7520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4568__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3472__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5673__A1 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input35_A mask_rev_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3684__B1 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2980 _6983_/Q VGND VGND VPWR VPWR _4296_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2991 hold2991/A VGND VGND VPWR VPWR _4251_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5425__A1 _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5399__A _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3987__A1 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3739__A1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4242__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7069__RESET_B _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6689__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold319 hold319/A VGND VGND VPWR VPWR _7314_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4164__A1 _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4390_ _4547_/A0 _4390_/A1 _4393_/S VGND VGND VPWR VPWR _4390_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2237_A _7281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6060_ _6060_/A1 _6019_/Y _6059_/X _6067_/B VGND VGND VPWR VPWR _7598_/D sky130_fd_sc_hd__a22o_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5664__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5011_ _5011_/A _5011_/B _5328_/B _5328_/A VGND VGND VPWR VPWR _5011_/Y sky130_fd_sc_hd__nand4_1
Xhold1008 hold3008/X VGND VGND VPWR VPWR _7543_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_140_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1019 hold3087/X VGND VGND VPWR VPWR _7351_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5801__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6208__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6613__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3690__A3 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6962_ _7160_/CLK _6962_/D fanout700/X VGND VGND VPWR VPWR _6962_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_93_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5913_ _5913_/A0 _5922_/A0 _5919_/S VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__mux2_1
X_6893_ _4127_/A1 _6893_/D _6843_/X VGND VGND VPWR VPWR _6893_/Q sky130_fd_sc_hd__dfrtp_4
X_5844_ _5844_/A0 _5853_/A0 _5847_/S VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5775_ _5775_/A0 hold20/X _5775_/S VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__mux2_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6392__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7514_ _7514_/CLK _7514_/D fanout744/X VGND VGND VPWR VPWR _7514_/Q sky130_fd_sc_hd__dfrtp_4
X_4726_ _4726_/A _4726_/B _4726_/C _5005_/A VGND VGND VPWR VPWR _4726_/Y sky130_fd_sc_hd__nand4_4
XFILLER_108_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7445_ _7525_/CLK _7445_/D fanout745/X VGND VGND VPWR VPWR _7445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4657_ _4657_/A _4657_/B _4657_/C _4657_/D VGND VGND VPWR VPWR _5248_/B sky130_fd_sc_hd__and4_4
XFILLER_135_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4155__A1 _4135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput80 spi_sck VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__clkbuf_2
X_3608_ _3645_/A1 _3607_/Y _3923_/S VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__mux2_1
Xhold820 _4523_/X VGND VGND VPWR VPWR _7173_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7376_ _7528_/CLK _7376_/D fanout729/X VGND VGND VPWR VPWR _7376_/Q sky130_fd_sc_hd__dfstp_4
X_4588_ _4562_/Y _4585_/Y _4593_/A _4674_/A VGND VGND VPWR VPWR _5295_/A sky130_fd_sc_hd__a2bb2o_4
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold842 _5842_/X VGND VGND VPWR VPWR _7441_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3902__A1 _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold853 hold853/A VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6327_ _6327_/A _6327_/B _6327_/C _6327_/D VGND VGND VPWR VPWR _6327_/Y sky130_fd_sc_hd__nor4_1
XFILLER_116_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold864 _5914_/X VGND VGND VPWR VPWR _7505_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold875 hold875/A VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4388__A _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3539_ _7430_/Q _3537_/X hold77/A _7526_/Q _3536_/X VGND VGND VPWR VPWR _3539_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmgmt_gpio_15_buff_inst _4161_/X VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_8
Xhold886 hold886/A VGND VGND VPWR VPWR _7168_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold897 hold897/A VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6258_ _6243_/X _6245_/X _6257_/Y VGND VGND VPWR VPWR _6258_/X sky130_fd_sc_hd__a21bo_1
Xhold2210 hold627/X VGND VGND VPWR VPWR _5716_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2221 _7241_/Q VGND VGND VPWR VPWR hold579/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2232 _7300_/Q VGND VGND VPWR VPWR hold707/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5209_ _4943_/B _4915_/C _4946_/Y _4774_/Y VGND VGND VPWR VPWR _5228_/A sky130_fd_sc_hd__o2bb2a_1
Xhold2243 _6915_/Q VGND VGND VPWR VPWR hold551/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2254 _5950_/X VGND VGND VPWR VPWR hold630/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6189_ _6181_/X _6075_/A _6186_/X _6184_/X _6188_/X VGND VGND VPWR VPWR _6189_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2265 hold649/X VGND VGND VPWR VPWR _5680_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5711__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1520 hold181/X VGND VGND VPWR VPWR _7580_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2276 _7347_/Q VGND VGND VPWR VPWR hold597/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1531 hold192/X VGND VGND VPWR VPWR _5836_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2287 _7406_/Q VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1542 hold144/X VGND VGND VPWR VPWR _5846_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1553 _4257_/X VGND VGND VPWR VPWR hold86/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2298 _5762_/X VGND VGND VPWR VPWR hold616/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1564 _6883_/Q VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__A1 _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1575 hold93/X VGND VGND VPWR VPWR _4350_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__7221__CLK_N _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1586 _5590_/X VGND VGND VPWR VPWR _5595_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1597 _5941_/X VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5012__A _5012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3969__A1 _7026_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4630__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5947__A _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6383__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6135__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6686__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4298__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4879__A_N _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4237__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5857__A _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3890_ _7178_/Q _4376_/B _5619_/B _3525_/X _7432_/Q VGND VGND VPWR VPWR _3890_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6374__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5295__C _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5560_ _5560_/A _5560_/B _5560_/C VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__and3_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4511_ _4511_/A0 _4547_/A0 _4514_/S VGND VGND VPWR VPWR _4511_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6126__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5491_ _5491_/A _5531_/B _5491_/C _5531_/C VGND VGND VPWR VPWR _5492_/D sky130_fd_sc_hd__and4_1
XFILLER_145_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7230_ _7255_/CLK _7230_/D fanout688/X VGND VGND VPWR VPWR _7230_/Q sky130_fd_sc_hd__dfstp_4
Xhold105 _3647_/A VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4442_ _4442_/A0 _5985_/A1 _4448_/S VGND VGND VPWR VPWR _4442_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold116 _7234_/Q VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold127 hold127/A VGND VGND VPWR VPWR _6924_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold138 hold138/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold149 hold149/A VGND VGND VPWR VPWR _7091_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5885__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7161_ _7268_/CLK _7161_/D _6861_/A VGND VGND VPWR VPWR _7161_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4373_ _5914_/A1 _4373_/A1 _4375_/S VGND VGND VPWR VPWR _4373_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3896__B1 _3862_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6119_/B _6112_/B _6112_/C _6119_/A VGND VGND VPWR VPWR _6112_/X sky130_fd_sc_hd__and4b_4
Xfanout607 _6082_/C VGND VGND VPWR VPWR _6144_/C sky130_fd_sc_hd__buf_6
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout618 _6110_/A VGND VGND VPWR VPWR _6317_/B sky130_fd_sc_hd__clkbuf_8
Xfanout629 _7084_/Q VGND VGND VPWR VPWR _4181_/S sky130_fd_sc_hd__buf_8
X_7092_ _7565_/CLK hold59/X fanout748/X VGND VGND VPWR VPWR _7092_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4358__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X VGND VGND VPWR VPWR _4164_/A1 sky130_fd_sc_hd__clkbuf_16
X_6043_ _7594_/Q _6429_/C VGND VGND VPWR VPWR _6447_/B sky130_fd_sc_hd__nor2_8
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ _7421_/CLK _6945_/D fanout715/X VGND VGND VPWR VPWR _7651_/A sky130_fd_sc_hd__dfrtp_1
X_6876_ _7201_/CLK _6876_/D fanout725/X VGND VGND VPWR VPWR _6876_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__3820__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_A _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5827_ _5827_/A0 _5881_/A1 hold33/X VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6365__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5758_ _5758_/A hold26/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__nand2_1
XFILLER_136_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4709_ _4748_/A _4844_/B _5387_/B VGND VGND VPWR VPWR _4709_/Y sky130_fd_sc_hd__nand3_4
XANTENNA_clkbuf_leaf_72_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6117__A2 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5689_ _5995_/A1 _5689_/A1 _5694_/S VGND VGND VPWR VPWR _5689_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5706__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7428_ _7576_/CLK _7428_/D fanout717/X VGND VGND VPWR VPWR _7428_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5325__B1 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6668__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5876__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7359_ _7360_/CLK _7359_/D fanout703/X VGND VGND VPWR VPWR _7359_/Q sky130_fd_sc_hd__dfstp_2
Xhold650 _5680_/X VGND VGND VPWR VPWR _7297_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold661 hold661/A VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6110__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold672 hold672/A VGND VGND VPWR VPWR _7333_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold683 hold683/A VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold694 hold694/A VGND VGND VPWR VPWR _7273_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5628__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2040 _5994_/X VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2051 _7118_/Q VGND VGND VPWR VPWR hold467/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2062 _7183_/Q VGND VGND VPWR VPWR hold475/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2073 hold491/X VGND VGND VPWR VPWR _4475_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input137_A wb_dat_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2084 _7374_/Q VGND VGND VPWR VPWR hold2084/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1350 _4320_/A1 VGND VGND VPWR VPWR hold2996/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2095 _7430_/Q VGND VGND VPWR VPWR hold2095/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 _4294_/B VGND VGND VPWR VPWR hold2994/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1372 _6790_/A1 VGND VGND VPWR VPWR hold3018/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 hold1445/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1394 _7338_/Q VGND VGND VPWR VPWR _5726_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4581__A _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3575__C1 _3574_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5867__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3893__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__A _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6292__A1 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4991_ _5183_/A _5183_/B _5034_/B _5158_/A VGND VGND VPWR VPWR _5037_/B sky130_fd_sc_hd__nand4_1
XANTENNA__6595__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5398__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5587__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6730_ _7150_/Q _6408_/A _6420_/A _6970_/Q _6729_/X VGND VGND VPWR VPWR _6730_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4491__A _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6895__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3942_ input61/X _5643_/A _3938_/X _3939_/X _3941_/X VGND VGND VPWR VPWR _3942_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3802__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ _6967_/Q _6420_/A _6421_/X _7006_/Q _6660_/X VGND VGND VPWR VPWR _6661_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6347__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3873_ _7544_/Q _3519_/X _3866_/X _3868_/X _3872_/X VGND VGND VPWR VPWR _3879_/A
+ sky130_fd_sc_hd__a2111o_2
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5612_ _5612_/A _5612_/B _5612_/C _5947_/C VGND VGND VPWR VPWR _5613_/S sky130_fd_sc_hd__and4_1
XANTENNA__3538__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6592_ _7468_/Q _6434_/B _6771_/A3 _6466_/X _7508_/Q VGND VGND VPWR VPWR _6592_/X
+ sky130_fd_sc_hd__a32o_1
X_5543_ _5543_/A _5543_/B _5543_/C VGND VGND VPWR VPWR _5543_/X sky130_fd_sc_hd__and3_1
XANTENNA__3581__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5474_ _5521_/B _5564_/B _5474_/C _5518_/A VGND VGND VPWR VPWR _5478_/A sky130_fd_sc_hd__nand4_2
XFILLER_105_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7213_ _7213_/CLK _7213_/D fanout701/X VGND VGND VPWR VPWR _7213_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4425_ _4425_/A _4425_/B _4425_/C _4424_/Y VGND VGND VPWR VPWR _4430_/B sky130_fd_sc_hd__nor4b_2
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7144_ _7266_/CLK _7144_/D fanout692/X VGND VGND VPWR VPWR _7144_/Q sky130_fd_sc_hd__dfstp_2
Xfanout404 _3590_/C VGND VGND VPWR VPWR _5731_/A sky130_fd_sc_hd__buf_4
X_4356_ _4356_/A0 _5585_/A0 _4357_/S VGND VGND VPWR VPWR _4356_/X sky130_fd_sc_hd__mux2_1
Xfanout415 _4364_/A VGND VGND VPWR VPWR _5803_/A sky130_fd_sc_hd__buf_8
Xfanout426 _5339_/A VGND VGND VPWR VPWR _5183_/A sky130_fd_sc_hd__buf_6
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout437 _4491_/C VGND VGND VPWR VPWR _4509_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout448 _3483_/X VGND VGND VPWR VPWR _4328_/A sky130_fd_sc_hd__clkbuf_16
X_7075_ _7075_/CLK _7075_/D _6865_/X VGND VGND VPWR VPWR _7075_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout459 _3464_/X VGND VGND VPWR VPWR _5612_/A sky130_fd_sc_hd__buf_12
XFILLER_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4287_ _3643_/Y _4287_/A1 _4289_/S VGND VGND VPWR VPWR _6977_/D sky130_fd_sc_hd__mux2_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6026_ _6019_/A _6929_/Q _7589_/Q _6025_/Y VGND VGND VPWR VPWR _7589_/D sky130_fd_sc_hd__o31a_1
XFILLER_74_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6586__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6440__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6928_ _7327_/CLK _6928_/D fanout703/X VGND VGND VPWR VPWR _6928_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6859_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6859_/X sky130_fd_sc_hd__and2_1
XANTENNA__6338__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1571_A _7509_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4551__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4349__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6121__A _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6510__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold480 _4499_/X VGND VGND VPWR VPWR _7153_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold491 hold491/A VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6274__A1 hold52/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1180 hold2868/X VGND VGND VPWR VPWR _7289_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1191 hold2877/X VGND VGND VPWR VPWR hold2878/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6577__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6329__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4461__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3655__A _7672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6501__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4210_ _4210_/A0 _5954_/A1 _4211_/S VGND VGND VPWR VPWR _4210_/X sky130_fd_sc_hd__mux2_1
XFILLER_130_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5190_ _5030_/C _5188_/X _5189_/X _5187_/X VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__a211o_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2809 hold993/X VGND VGND VPWR VPWR _4537_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4141_ _7578_/Q _4142_/A _4140_/Y VGND VGND VPWR VPWR _4141_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_122_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4917__C _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6265__B2 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4072_ hold1/A hold12/A _4074_/S VGND VGND VPWR VPWR _6886_/D sky130_fd_sc_hd__mux2_1
XFILLER_110_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6568__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4974_ _4996_/A _4974_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _5342_/C sky130_fd_sc_hd__and4_1
XANTENNA__7073__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5240__A2 _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6713_ _7003_/Q _6455_/B _6466_/C _6462_/C _6712_/X VGND VGND VPWR VPWR _6713_/X
+ sky130_fd_sc_hd__a41o_1
X_3925_ _7046_/Q _5830_/C _4539_/C _4388_/B VGND VGND VPWR VPWR _3925_/X sky130_fd_sc_hd__and4_1
XFILLER_189_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold2853_A _6913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6644_ _7502_/Q _6447_/C _6769_/A3 _6420_/C _7398_/Q VGND VGND VPWR VPWR _6644_/X
+ sky130_fd_sc_hd__a32o_1
X_3856_ _3856_/A _3856_/B VGND VGND VPWR VPWR _3856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6575_ _7356_/Q _6413_/C _6459_/C _6462_/X _7364_/Q VGND VGND VPWR VPWR _6575_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3787_ _7247_/Q _5947_/A _5614_/B _3515_/X _7238_/Q VGND VGND VPWR VPWR _3787_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3565__A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6740__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4751__A1 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__A2 _3552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5526_ _5038_/A _5282_/C _5282_/D _5525_/X VGND VGND VPWR VPWR _5526_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6910__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5457_ _5457_/A _5457_/B VGND VGND VPWR VPWR _5457_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4408_ _4441_/A0 _5975_/A0 _4422_/S VGND VGND VPWR VPWR _4408_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5388_ _4596_/X _5387_/C _5387_/D _5081_/A _5387_/X VGND VGND VPWR VPWR _5521_/A
+ sky130_fd_sc_hd__a41oi_4
XFILLER_87_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7127_ _7395_/CLK _7127_/D fanout737/X VGND VGND VPWR VPWR _7127_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4339_ _4339_/A0 _5817_/A1 _4339_/S VGND VGND VPWR VPWR _4339_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout769_A _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6256__A1 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4827__C _4983_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7058_ _7179_/CLK _7058_/D fanout699/X VGND VGND VPWR VPWR _7058_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6009_ _6932_/Q _6009_/B VGND VGND VPWR VPWR _6009_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7416__CLK _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__A _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6731__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire679 _4833_/A VGND VGND VPWR VPWR _5295_/D sky130_fd_sc_hd__buf_4
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input65_A mgmt_gpio_in[36] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6786__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5298__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3848__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6247__B2 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4245__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3710_ _7579_/Q _3501_/X _4248_/S _4150_/A1 _3709_/X VGND VGND VPWR VPWR _3710_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3784__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4690_ _5328_/A _5328_/B VGND VGND VPWR VPWR _4690_/Y sky130_fd_sc_hd__nand2_8
X_3641_ _7372_/Q _5758_/A _3527_/X _6916_/Q _3640_/X VGND VGND VPWR VPWR _3642_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6183__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6722__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5930__A0 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6360_ _7009_/Q _6082_/C _6081_/X _6097_/X _7185_/Q VGND VGND VPWR VPWR _6360_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3536__A2 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3572_ _3609_/A1 _3570_/Y _3923_/S VGND VGND VPWR VPWR _3572_/X sky130_fd_sc_hd__mux2_1
X_5311_ _5311_/A _5311_/B _5488_/A VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__and3_1
XFILLER_142_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ _7061_/Q _6032_/Y _6081_/X _7192_/Q _6290_/X VGND VGND VPWR VPWR _6291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5804__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5289__A2 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3307 _7605_/Q VGND VGND VPWR VPWR _6192_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6486__B2 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5242_ _5222_/A _5248_/B _5453_/A _4941_/B VGND VGND VPWR VPWR _5545_/A sky130_fd_sc_hd__a31o_1
Xhold3318 _7626_/Q VGND VGND VPWR VPWR _6776_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_114_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3329 _6473_/X VGND VGND VPWR VPWR _7615_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_30_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7531_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2606 _7154_/Q VGND VGND VPWR VPWR hold967/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2617 hold929/X VGND VGND VPWR VPWR _5995_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5173_ _5495_/C1 _5528_/A3 _5046_/A _5046_/B _4690_/Y VGND VGND VPWR VPWR _5173_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_96_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2628 hold721/X VGND VGND VPWR VPWR _4532_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2639 hold705/X VGND VGND VPWR VPWR _4454_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1905 _5699_/X VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1916 hold284/X VGND VGND VPWR VPWR _5754_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4124_ _4058_/B _4123_/B _4123_/Y _7073_/Q VGND VGND VPWR VPWR _7073_/D sky130_fd_sc_hd__a22o_1
Xhold1927 _5654_/X VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1938 hold164/X VGND VGND VPWR VPWR _5820_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1949 _7570_/Q VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xinput1 debug_mode VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_4
XFILLER_110_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4055_ _4076_/B _4058_/A _3856_/A _4054_/X VGND VGND VPWR VPWR _6894_/D sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_45_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7572_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4155__S _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4382__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4957_ _4953_/X _4956_/Y _4955_/X VGND VGND VPWR VPWR _4958_/C sky130_fd_sc_hd__a21oi_1
X_3908_ _7230_/Q _3617_/X _3682_/X _7225_/Q _3907_/X VGND VGND VPWR VPWR _3913_/B
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3775__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4972__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4888_ _4840_/D _4888_/B _4888_/C _4910_/D VGND VGND VPWR VPWR _4888_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_131_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6627_ _7358_/Q _6459_/B _6428_/X _6408_/B _7382_/Q VGND VGND VPWR VPWR _6627_/X
+ sky130_fd_sc_hd__a32o_1
X_3839_ _7043_/Q _4370_/A _3673_/X _7199_/Q VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5516__A3 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5921__A0 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6558_ _7443_/Q _6574_/B _6574_/C _6466_/X _7507_/Q VGND VGND VPWR VPWR _6558_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5509_ _4726_/Y _4796_/Y _5509_/A3 _4930_/B _5237_/C VGND VGND VPWR VPWR _5510_/C
+ sky130_fd_sc_hd__o311a_1
X_6489_ _7552_/Q _6408_/A _6408_/D _7536_/Q _6488_/X VGND VGND VPWR VPWR _6494_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6477__A1 _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6477__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4488__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4838__B _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6229__A1 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6244__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5204__A2 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3766__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4963__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6165__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6180__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3933__A _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4748__B _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5979__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2015_A _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__A1 _7446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5443__A2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__B2 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3454__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ _5995_/A1 _5860_/A1 _5865_/S VGND VGND VPWR VPWR _5860_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_817 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4811_ _5158_/B _5138_/A _5138_/B _4811_/D VGND VGND VPWR VPWR _4812_/C sky130_fd_sc_hd__nand4_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ _5791_/A0 _5881_/A1 hold48/X VGND VGND VPWR VPWR _5791_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7530_ _7565_/CLK _7530_/D fanout748/X VGND VGND VPWR VPWR _7530_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3757__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4742_ _5407_/A1 _5282_/A VGND VGND VPWR VPWR _5073_/B sky130_fd_sc_hd__nand2b_4
X_7461_ _7478_/CLK _7461_/D fanout715/X VGND VGND VPWR VPWR _7461_/Q sky130_fd_sc_hd__dfrtp_4
X_4673_ _4674_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _4673_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__6156__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6412_ _6463_/A _6468_/C _6413_/C VGND VGND VPWR VPWR _6420_/A sky130_fd_sc_hd__and3_4
XANTENNA__5903__A0 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3624_ _7300_/Q _3848_/A2 _3562_/C _5776_/A _7388_/Q VGND VGND VPWR VPWR _3624_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3509__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7392_ _7562_/CLK _7392_/D fanout739/X VGND VGND VPWR VPWR _7392_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_190_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6343_ _7018_/Q _6121_/C _6086_/X _6342_/X VGND VGND VPWR VPWR _6343_/X sky130_fd_sc_hd__a31o_1
X_3555_ _5740_/A _4551_/A _5938_/A VGND VGND VPWR VPWR _5776_/A sky130_fd_sc_hd__and3_4
XFILLER_155_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6274_ hold52/A _6080_/A _6274_/A3 _6085_/X _7502_/Q VGND VGND VPWR VPWR _6274_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3104 _5885_/X VGND VGND VPWR VPWR hold3104/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3486_ _5590_/A _4328_/A _5612_/B VGND VGND VPWR VPWR _3486_/X sky130_fd_sc_hd__and3_4
Xhold3115 _6997_/Q VGND VGND VPWR VPWR _4317_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3126 hold3126/A VGND VGND VPWR VPWR _4492_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3562__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3137 _4462_/X VGND VGND VPWR VPWR hold3137/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5131__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5225_ _4933_/B _4907_/B _4918_/D _5102_/B wire658/X VGND VGND VPWR VPWR _5228_/C
+ sky130_fd_sc_hd__a32oi_4
Xhold2403 hold689/X VGND VGND VPWR VPWR _4508_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3148 _7423_/Q VGND VGND VPWR VPWR hold3148/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2414 _7211_/Q VGND VGND VPWR VPWR hold855/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3159 _7167_/Q VGND VGND VPWR VPWR hold3159/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2425 _5638_/X VGND VGND VPWR VPWR hold702/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2436 _7173_/Q VGND VGND VPWR VPWR hold819/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1702 _7513_/Q VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2447 hold663/X VGND VGND VPWR VPWR _4544_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5156_ _5156_/A _5156_/B _5156_/C VGND VGND VPWR VPWR _5160_/B sky130_fd_sc_hd__nand3_1
Xhold2458 _4373_/X VGND VGND VPWR VPWR hold830/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1713 _5684_/X VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3693__A1 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1724 hold306/X VGND VGND VPWR VPWR _5890_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2469 _6876_/Q VGND VGND VPWR VPWR hold873/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1735 _7094_/Q VGND VGND VPWR VPWR hold355/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4107_ _4107_/A _4117_/B VGND VGND VPWR VPWR _4107_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1746 hold292/X VGND VGND VPWR VPWR _4326_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1757 _5922_/X VGND VGND VPWR VPWR hold416/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5087_ _4717_/Y _4960_/A _5086_/Y _5085_/Y VGND VGND VPWR VPWR _5087_/Y sky130_fd_sc_hd__o211ai_1
Xhold1768 _7339_/Q VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1779 hold283/X VGND VGND VPWR VPWR _7267_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4038_ _4037_/Y _4029_/X _4025_/A _6901_/Q VGND VGND VPWR VPWR _4038_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6395__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5709__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5989_/A0 _5998_/A1 _5991_/S VGND VGND VPWR VPWR _5989_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3748__A2 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3737__B _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_50 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7659_ _7659_/A VGND VGND VPWR VPWR _7659_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_61 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _7499_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1749_A _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3920__A2 hold77/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input167_A wb_sel_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput190 _3422_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XANTENNA__3684__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3684__B2 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2970 _4403_/X VGND VGND VPWR VPWR hold2970/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input28_A mask_rev_in[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2981 hold2981/A VGND VGND VPWR VPWR hold2981/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2992 _4251_/X VGND VGND VPWR VPWR hold2992/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_leaf_67_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5425__A2 _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5399__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3987__A2 _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5189__A1 _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6386__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3928__A _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3739__A2 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4750__C _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3647__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6689__A1 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6153__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold309 hold309/A VGND VGND VPWR VPWR _7039_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4759__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3663__A _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_4_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3911__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_12__f_wb_clk_i clkbuf_3_6_0_wb_clk_i/X VGND VGND VPWR VPWR _7111_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5010_ _4996_/A _5339_/C _5216_/A VGND VGND VPWR VPWR _5011_/A sky130_fd_sc_hd__o21a_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 hold3026/X VGND VGND VPWR VPWR hold3027/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6961_ _7238_/CLK _6961_/D fanout691/X VGND VGND VPWR VPWR _6961_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_53_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5912_ _5912_/A0 _5912_/A1 _5919_/S VGND VGND VPWR VPWR _5912_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3978__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6892_ _7075_/CLK _6892_/D _6842_/X VGND VGND VPWR VPWR _6892_/Q sky130_fd_sc_hd__dfrtp_4
X_5843_ _5843_/A0 _5978_/A0 _5847_/S VGND VGND VPWR VPWR _5843_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6377__B1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5774_ _5774_/A0 _5999_/A1 _5775_/S VGND VGND VPWR VPWR _5774_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7513_ _7531_/CLK _7513_/D fanout744/X VGND VGND VPWR VPWR _7513_/Q sky130_fd_sc_hd__dfrtp_4
X_4725_ _5222_/B _4726_/B _4726_/C _5005_/A VGND VGND VPWR VPWR _4725_/X sky130_fd_sc_hd__and4_2
XANTENNA__6129__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4656_ _4667_/A _4899_/A2 _4657_/C _4657_/B VGND VGND VPWR VPWR _4889_/A sky130_fd_sc_hd__o211ai_2
X_7444_ _7565_/CLK _7444_/D fanout748/X VGND VGND VPWR VPWR _7444_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3607_ _3575_/X _3607_/B _3607_/C VGND VGND VPWR VPWR _3607_/Y sky130_fd_sc_hd__nand3b_4
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR _4176_/B sky130_fd_sc_hd__buf_4
Xinput81 spi_sdo VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__buf_2
Xhold810 _4502_/X VGND VGND VPWR VPWR _7156_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4587_ _4674_/A _4593_/A _4687_/B VGND VGND VPWR VPWR _4755_/A sky130_fd_sc_hd__a21boi_4
Xhold821 hold821/A VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7375_ _7528_/CLK _7375_/D fanout729/X VGND VGND VPWR VPWR _7375_/Q sky130_fd_sc_hd__dfstp_2
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR _4140_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold832 hold832/A VGND VGND VPWR VPWR _6877_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold843 hold843/A VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__A2 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6326_ _7052_/Q _6087_/X _6120_/X _7017_/Q _6325_/X VGND VGND VPWR VPWR _6327_/D
+ sky130_fd_sc_hd__a221o_1
X_3538_ _4551_/A _3682_/A _5938_/C VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__and3_4
Xhold854 _4362_/X VGND VGND VPWR VPWR _7034_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4388__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold865 hold865/A VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold876 _5934_/X VGND VGND VPWR VPWR _7523_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold887 hold887/A VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold898 _5755_/X VGND VGND VPWR VPWR _7364_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5104__A1 _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6257_ _6257_/A _6257_/B _6257_/C _6257_/D VGND VGND VPWR VPWR _6257_/Y sky130_fd_sc_hd__nor4_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2200 hold645/X VGND VGND VPWR VPWR _5878_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6301__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3469_ _6901_/Q _6900_/Q _4007_/B VGND VGND VPWR VPWR _3469_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout584_A _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2211 _5716_/X VGND VGND VPWR VPWR hold628/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2222 hold579/X VGND VGND VPWR VPWR _5610_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5208_ _5561_/A1 _4796_/Y _5516_/A3 _4930_/C VGND VGND VPWR VPWR _5208_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2233 hold707/X VGND VGND VPWR VPWR _5683_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2244 hold551/X VGND VGND VPWR VPWR _4196_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6188_ _7442_/Q _6097_/X _6121_/X _7306_/Q _6187_/X VGND VGND VPWR VPWR _6188_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1510 _7545_/Q VGND VGND VPWR VPWR hold176/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2255 _7554_/Q VGND VGND VPWR VPWR hold651/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1521 _7569_/Q VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2266 _6923_/Q VGND VGND VPWR VPWR hold577/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5139_ _5013_/X _5139_/B _5139_/C _5139_/D VGND VGND VPWR VPWR _5139_/X sky130_fd_sc_hd__and4b_1
Xhold2277 hold597/X VGND VGND VPWR VPWR _5736_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1532 _5836_/X VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2288 hold601/X VGND VGND VPWR VPWR _5802_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1543 _5846_/X VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2299 _6952_/Q VGND VGND VPWR VPWR hold667/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1554 _6956_/Q VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1565 hold196/X VGND VGND VPWR VPWR _4183_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1576 _4350_/X VGND VGND VPWR VPWR hold94/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5407__A2 _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1587 _5594_/X VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1598 _7521_/Q VGND VGND VPWR VPWR hold230/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5012__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3969__A2 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5947__B _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6368__B1 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5591__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4579__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6540__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3247_A _7327_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4854__B1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4745__C _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output301_A _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5857__B _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6359__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4510_ _4510_/A0 _5582_/A0 _4514_/S VGND VGND VPWR VPWR _4510_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3593__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5490_ _4997_/A _4952_/B _5052_/B _5489_/X VGND VGND VPWR VPWR _5532_/B sky130_fd_sc_hd__a211oi_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold106 _5938_/X VGND VGND VPWR VPWR _5946_/S sky130_fd_sc_hd__buf_6
X_4441_ _4441_/A0 _5993_/A1 _4448_/S VGND VGND VPWR VPWR _4441_/X sky130_fd_sc_hd__mux2_1
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold139 hold139/A VGND VGND VPWR VPWR _7509_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7160_ _7160_/CLK _7160_/D fanout700/X VGND VGND VPWR VPWR _7160_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ _4553_/A0 _4372_/A1 _4375_/S VGND VGND VPWR VPWR _4372_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6112_/C _6119_/B _6121_/A _6119_/A VGND VGND VPWR VPWR _6111_/X sky130_fd_sc_hd__and4bb_4
Xfanout608 _3444_/Y VGND VGND VPWR VPWR _6082_/C sky130_fd_sc_hd__buf_8
X_7091_ _7522_/CLK _7091_/D fanout748/X VGND VGND VPWR VPWR _7091_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _7592_/Q VGND VGND VPWR VPWR _6110_/A sky130_fd_sc_hd__buf_6
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__C1 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6042_ _7594_/Q _6429_/C VGND VGND VPWR VPWR _6042_/X sky130_fd_sc_hd__and2_4
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5113__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6944_ _7314_/CLK _6944_/D _4079_/A VGND VGND VPWR VPWR _7650_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__4952__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5767__B _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3820__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6875_ _7201_/CLK _6875_/D fanout725/X VGND VGND VPWR VPWR _6875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_179_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5826_ _5826_/A0 _5826_/A1 hold33/X VGND VGND VPWR VPWR _5826_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5757_ _5757_/A0 _5955_/A1 _5757_/S VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6770__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4708_ _4887_/B _4945_/A _5387_/B VGND VGND VPWR VPWR _4811_/D sky130_fd_sc_hd__and3_4
X_5688_ _5949_/A1 _5688_/A1 _5694_/S VGND VGND VPWR VPWR _5688_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6117__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7427_ _7471_/CLK _7427_/D fanout729/X VGND VGND VPWR VPWR _7427_/Q sky130_fd_sc_hd__dfrtp_2
X_4639_ _4667_/A _5494_/B2 _4636_/Y VGND VGND VPWR VPWR _4641_/B sky130_fd_sc_hd__o21ai_4
XANTENNA_hold1447_A _4085_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold640 hold640/A VGND VGND VPWR VPWR _7515_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7358_ _7576_/CLK _7358_/D fanout731/X VGND VGND VPWR VPWR _7358_/Q sky130_fd_sc_hd__dfrtp_4
Xhold651 hold651/A VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold662 hold662/A VGND VGND VPWR VPWR _7369_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6110__C _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5007__B _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold673 hold673/A VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold684 hold684/A VGND VGND VPWR VPWR _7201_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6309_ _7012_/Q _6384_/A4 _6120_/B _6317_/B VGND VGND VPWR VPWR _6309_/X sky130_fd_sc_hd__a31o_1
Xhold695 hold695/A VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmgmt_gpio_30_buff_inst _4164_/X VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__clkbuf_8
X_7289_ _7327_/CLK _7289_/D fanout703/X VGND VGND VPWR VPWR _7289_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2030 hold443/X VGND VGND VPWR VPWR _5708_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__B2 _7673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2041 _7186_/Q VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2052 hold467/X VGND VGND VPWR VPWR _4457_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7416__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2063 hold475/X VGND VGND VPWR VPWR _4535_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2074 _7488_/Q VGND VGND VPWR VPWR hold513/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1340 hold3210/X VGND VGND VPWR VPWR _7066_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2085 hold2085/A VGND VGND VPWR VPWR _5766_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6038__C1 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1351 _4319_/A1 VGND VGND VPWR VPWR hold2989/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2096 hold2096/A VGND VGND VPWR VPWR _5829_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1362 _4291_/B VGND VGND VPWR VPWR hold2972/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1373 _6786_/B VGND VGND VPWR VPWR hold3023/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6589__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1384 _6788_/B VGND VGND VPWR VPWR hold3265/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1395 hold1435/X VGND VGND VPWR VPWR hold1436/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4581__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3811__A1 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3478__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6356__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input95_A usr1_vcc_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6761__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3575__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3925__B _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5316__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5316__B2 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3878__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4756__B _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3660__B _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4248__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4055__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4990_ _5183_/A _5203_/C _5034_/B _5183_/B VGND VGND VPWR VPWR _5037_/C sky130_fd_sc_hd__nand4_1
XANTENNA__5587__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3941_ _7551_/Q _3508_/X _4422_/S input43/X _3940_/X VGND VGND VPWR VPWR _3941_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4491__B _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6660_ _7112_/Q _6651_/B _6426_/X _6659_/X VGND VGND VPWR VPWR _6660_/X sky130_fd_sc_hd__a31o_1
X_3872_ _7568_/Q _3872_/A2 _3637_/C _3869_/X _3871_/X VGND VGND VPWR VPWR _3872_/X
+ sky130_fd_sc_hd__a311o_4
XFILLER_149_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5611_ _5611_/A0 _5955_/A1 _5611_/S VGND VGND VPWR VPWR _5611_/X sky130_fd_sc_hd__mux2_1
X_6591_ _7452_/Q _6443_/X _6446_/X _7524_/Q _6574_/X VGND VGND VPWR VPWR _6591_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_192_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5807__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5542_ _4622_/Y _4726_/Y _4748_/Y _5512_/A _5462_/X VGND VGND VPWR VPWR _5543_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_129_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6504__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5473_ _4791_/A _5473_/B _5473_/C _5473_/D VGND VGND VPWR VPWR _5518_/A sky130_fd_sc_hd__and4b_1
XANTENNA__5307__B2 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3581__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7212_ _7212_/CLK _7212_/D fanout721/X VGND VGND VPWR VPWR _7212_/Q sky130_fd_sc_hd__dfrtp_4
X_4424_ _7102_/Q _4424_/B VGND VGND VPWR VPWR _4424_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7143_ _7266_/CLK _7143_/D fanout692/X VGND VGND VPWR VPWR _7143_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4355_ _4355_/A0 _5788_/A1 _4357_/S VGND VGND VPWR VPWR _4355_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout405 _3492_/X VGND VGND VPWR VPWR _3590_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_98_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout416 hold47/X VGND VGND VPWR VPWR _4364_/A sky130_fd_sc_hd__buf_8
XFILLER_101_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout427 _4997_/B VGND VGND VPWR VPWR _5339_/A sky130_fd_sc_hd__buf_6
X_7074_ _4127_/A1 _7074_/D _6864_/X VGND VGND VPWR VPWR _7074_/Q sky130_fd_sc_hd__dfrtp_1
Xfanout438 hold1585/X VGND VGND VPWR VPWR _4491_/C sky130_fd_sc_hd__buf_8
Xfanout449 _5938_/B VGND VGND VPWR VPWR _5640_/B sky130_fd_sc_hd__buf_8
XFILLER_59_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4286_ _4289_/S _6789_/A2 _4285_/Y VGND VGND VPWR VPWR _6976_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__4666__B _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6025_ _6112_/B _6136_/B _6019_/A VGND VGND VPWR VPWR _6025_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout547_A hold1428/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6927_ _7327_/CLK _6927_/D fanout703/X VGND VGND VPWR VPWR _6927_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6858_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6858_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout714_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6338__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold125_A _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5809_ _5809_/A0 _5953_/A1 _5811_/S VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6743__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6789_ _6789_/A1 _6789_/A2 _6788_/Y VGND VGND VPWR VPWR _7633_/D sky130_fd_sc_hd__o21ai_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6121__B _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6510__A3 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold470 _5808_/X VGND VGND VPWR VPWR _7411_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold481 hold481/A VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold492 _4475_/X VGND VGND VPWR VPWR _7133_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1170 hold1170/A VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XANTENNA_input10_A mask_rev_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1181 hold3226/X VGND VGND VPWR VPWR hold3227/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1192 _5593_/X VGND VGND VPWR VPWR _7226_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6577__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_786 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6734__B1 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3655__B _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6031__B _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3671__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4140_ _4142_/A _4140_/B VGND VGND VPWR VPWR _4140_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_hold2045_A _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4917__D _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6265__A2 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4071_ hold15/A hold1/A _4074_/S VGND VGND VPWR VPWR _6887_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4276__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2212_A _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4933__C _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4973_ _5480_/B2 _4748_/Y _4814_/Y _4826_/Y VGND VGND VPWR VPWR _5200_/C sky130_fd_sc_hd__a211o_2
XANTENNA__3787__B1 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6712_ _7169_/Q _6408_/D _6427_/X _7119_/Q _6711_/X VGND VGND VPWR VPWR _6712_/X
+ sky130_fd_sc_hd__a221o_4
X_3924_ _3923_/X _3924_/A1 _3996_/A VGND VGND VPWR VPWR _7215_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3549__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6643_ _7550_/Q _6419_/A _6467_/X _7422_/Q _6642_/X VGND VGND VPWR VPWR _6643_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6725__B1 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3855_ _3855_/A _3855_/B _3855_/C VGND VGND VPWR VPWR _3856_/B sky130_fd_sc_hd__and3_4
XFILLER_149_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3539__B1 hold77/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4441__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4200__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3786_ _7165_/Q _3663_/X _3666_/X _7014_/Q _3785_/X VGND VGND VPWR VPWR _3792_/C
+ sky130_fd_sc_hd__a221o_1
X_6574_ _7444_/Q _6574_/B _6574_/C VGND VGND VPWR VPWR _6574_/X sky130_fd_sc_hd__and3_1
XANTENNA__6740__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3565__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5525_ _4817_/X _5453_/C _5395_/X _5521_/Y _5524_/X VGND VGND VPWR VPWR _5525_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4751__A2 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5456_ _5545_/C _5541_/D _5456_/C _5543_/A VGND VGND VPWR VPWR _5457_/A sky130_fd_sc_hd__and4b_1
XFILLER_59_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5161__C1 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4407_ _4422_/S _4215_/X _4406_/Y _5956_/C VGND VGND VPWR VPWR _4423_/S sky130_fd_sc_hd__o211a_4
XANTENNA__5700__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5387_ _4748_/A _5387_/B _5387_/C _5387_/D VGND VGND VPWR VPWR _5387_/X sky130_fd_sc_hd__and4b_1
XANTENNA_fanout497_A _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7126_ _7186_/CLK _7126_/D _6839_/A VGND VGND VPWR VPWR _7126_/Q sky130_fd_sc_hd__dfrtp_4
X_4338_ _4338_/A0 _5585_/A0 _4339_/S VGND VGND VPWR VPWR _4338_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A debug_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6256__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4269_ _4269_/A0 _5647_/A0 _4270_/S VGND VGND VPWR VPWR _4269_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7057_ _7181_/CLK _7057_/D fanout724/X VGND VGND VPWR VPWR _7057_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4267__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6008_ _6005_/Y _6006_/X _6018_/A VGND VGND VPWR VPWR _7584_/D sky130_fd_sc_hd__o21a_1
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6716__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire603 _4058_/Y VGND VGND VPWR VPWR _4075_/S sky130_fd_sc_hd__buf_4
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1946_A _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire658 _4715_/Y VGND VGND VPWR VPWR wire658/X sky130_fd_sc_hd__buf_2
Xwire669 _5118_/A VGND VGND VPWR VPWR _4810_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input58_A mgmt_gpio_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4258__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5910__S hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5470__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3410__1 _4127_/A1 VGND VGND VPWR VPWR _6881_/CLK sky130_fd_sc_hd__inv_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6707__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3784__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3666__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _7396_/Q _5803_/A _3933_/A _3564_/X _7364_/Q VGND VGND VPWR VPWR _3640_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ _6893_/Q _7073_/Q VGND VGND VPWR VPWR _3996_/A sky130_fd_sc_hd__nand2_8
XANTENNA__3536__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3941__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5310_ _5494_/B2 _4783_/Y _4789_/Y _4744_/Y _5153_/B VGND VGND VPWR VPWR _5488_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6290_ _7187_/Q _6099_/D _6081_/C _6136_/B _6121_/C VGND VGND VPWR VPWR _6290_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_182_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6486__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3308 _6192_/X VGND VGND VPWR VPWR _7605_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5241_ _4935_/X _5243_/C _5239_/X VGND VGND VPWR VPWR _5244_/C sky130_fd_sc_hd__a21o_1
XFILLER_142_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3319 hold44/A VGND VGND VPWR VPWR _4024_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5694__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5172_ _4877_/A _4970_/C _5018_/B _5180_/A VGND VGND VPWR VPWR _5172_/X sky130_fd_sc_hd__a22o_1
Xhold2607 hold967/X VGND VGND VPWR VPWR _4500_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2618 _5995_/X VGND VGND VPWR VPWR hold930/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2629 _4532_/X VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6238__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4123_ _4123_/A _4123_/B _4123_/C VGND VGND VPWR VPWR _4123_/Y sky130_fd_sc_hd__nand3_1
Xhold1906 _7160_/Q VGND VGND VPWR VPWR hold296/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1917 _7275_/Q VGND VGND VPWR VPWR hold265/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5820__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1928 _7048_/Q VGND VGND VPWR VPWR hold338/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1939 _5820_/X VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 debug_oeb VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4054_ _6910_/Q _6909_/Q _6908_/Q _4062_/A _4054_/B1 VGND VGND VPWR VPWR _4054_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5997__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4382__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4960__A _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ _4956_/A _4956_/B VGND VGND VPWR VPWR _4956_/Y sky130_fd_sc_hd__nand2_2
X_3907_ _7408_/Q _4364_/A _5947_/A _4485_/A _7143_/Q VGND VGND VPWR VPWR _3907_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4972__A2 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4887_ _4840_/D _4887_/B _4945_/A _4887_/D VGND VGND VPWR VPWR _4887_/X sky130_fd_sc_hd__and4b_2
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3576__A _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6626_ _7534_/Q _6058_/X _6409_/X _7406_/Q VGND VGND VPWR VPWR _6626_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout412_A _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6174__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3838_ _7377_/Q _5740_/A _5983_/A _3658_/X _7114_/Q VGND VGND VPWR VPWR _3838_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6713__A3 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6557_ _7563_/Q _6419_/C _6434_/X _7467_/Q _6556_/X VGND VGND VPWR VPWR _6557_/X
+ sky130_fd_sc_hd__a221o_2
X_3769_ input29/X _3503_/X _3520_/X _7442_/Q _3768_/X VGND VGND VPWR VPWR _3769_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_152_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3932__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5508_ _5508_/A _5508_/B _5508_/C VGND VGND VPWR VPWR _5575_/A sky130_fd_sc_hd__and3_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6488_ _7472_/Q _6466_/C _6441_/X _6423_/X _7328_/Q VGND VGND VPWR VPWR _6488_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6477__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5439_ _5059_/A _5203_/A _5180_/B _5049_/C _5058_/C VGND VGND VPWR VPWR _5439_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_2__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7109_ _4164_/A1 _7109_/D fanout751/X VGND VGND VPWR VPWR _7109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5730__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_user_clock clkbuf_0_user_clock/X VGND VGND VPWR VPWR _4163_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_75_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5988__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4573__C _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input112_A wb_adr_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4412__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3766__A3 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3486__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire433 _5158_/B VGND VGND VPWR VPWR _5295_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_128_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5905__S hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3933__B _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_775 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X VGND VGND VPWR VPWR _7630_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_124_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3652__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5140__A2 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6640__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6900__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4810_ _5138_/A _5138_/B _4810_/C _5453_/B VGND VGND VPWR VPWR _4812_/B sky130_fd_sc_hd__nand4_1
XFILLER_22_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _5790_/A0 _5826_/A1 hold48/X VGND VGND VPWR VPWR _5790_/X sky130_fd_sc_hd__mux2_1
X_4741_ _5074_/B _4814_/C VGND VGND VPWR VPWR _4741_/Y sky130_fd_sc_hd__nand2_8
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2377_A _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7460_ _7556_/CLK _7460_/D fanout731/X VGND VGND VPWR VPWR _7460_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4672_ _4861_/A _4861_/B _4667_/Y _4669_/X VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__a211o_4
XFILLER_174_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6411_ _6467_/A _6462_/C _6409_/X _6410_/X _6466_/D VGND VGND VPWR VPWR _6411_/Y
+ sky130_fd_sc_hd__a2111oi_2
X_3623_ _3623_/A _3623_/B _3623_/C _3623_/D VGND VGND VPWR VPWR _3643_/A sky130_fd_sc_hd__nor4_2
XANTENNA__3509__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7391_ _7562_/CLK _7391_/D fanout739/X VGND VGND VPWR VPWR _7391_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5815__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3914__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6342_ _7058_/Q _6332_/B _6388_/A3 _6121_/X _6990_/Q VGND VGND VPWR VPWR _6342_/X
+ sky130_fd_sc_hd__a32o_1
X_3554_ _4176_/B _3552_/X _3553_/X input42/X _3551_/X VGND VGND VPWR VPWR _3568_/C
+ sky130_fd_sc_hd__a221o_1
X_3485_ _3511_/C hold46/X _3485_/C VGND VGND VPWR VPWR _3485_/X sky130_fd_sc_hd__and3b_4
X_6273_ _7462_/Q _6080_/X _6269_/X _6270_/X _6272_/X VGND VGND VPWR VPWR _6280_/A
+ sky130_fd_sc_hd__a2111o_1
Xhold3105 _7132_/Q VGND VGND VPWR VPWR hold3105/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3116 hold3116/A VGND VGND VPWR VPWR hold3116/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3127 _7026_/Q VGND VGND VPWR VPWR hold3127/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_143_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5224_ _5224_/A _5349_/A _5224_/C VGND VGND VPWR VPWR _5228_/B sky130_fd_sc_hd__nor3_1
XANTENNA__3562__C _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3138 _7031_/Q VGND VGND VPWR VPWR hold3138/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2404 _4508_/X VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3149 hold3149/A VGND VGND VPWR VPWR _5822_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2415 hold855/X VGND VGND VPWR VPWR _5584_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2426 _7020_/Q VGND VGND VPWR VPWR hold687/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2437 hold819/X VGND VGND VPWR VPWR _4523_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1703 hold216/X VGND VGND VPWR VPWR _5923_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2448 _4544_/X VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5155_ _4625_/Y _4690_/Y _4802_/Y _4796_/Y _4706_/Y VGND VGND VPWR VPWR _5156_/C
+ sky130_fd_sc_hd__o32a_1
Xhold1714 _7544_/Q VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2459 _7163_/Q VGND VGND VPWR VPWR hold915/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3693__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1725 _5890_/X VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1736 hold355/X VGND VGND VPWR VPWR _4442_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4106_ _7585_/Q _7584_/Q _7586_/Q _7587_/Q VGND VGND VPWR VPWR _4107_/A sky130_fd_sc_hd__nand4bb_4
X_5086_ _5094_/A _5086_/B VGND VGND VPWR VPWR _5086_/Y sky130_fd_sc_hd__nand2_1
Xhold1747 _4326_/X VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1758 _7538_/Q VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1769 hold118/X VGND VGND VPWR VPWR _5727_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4166__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4037_ _6901_/Q _6900_/Q _6902_/Q VGND VGND VPWR VPWR _4037_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6631__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ _5988_/A0 _5997_/A1 _5991_/S VGND VGND VPWR VPWR _5988_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _4954_/A _5453_/A _4939_/C _4940_/D VGND VGND VPWR VPWR _4941_/A sky130_fd_sc_hd__and4_1
XANTENNA__4840__D _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_40 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3737__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7658_ _7658_/A VGND VGND VPWR VPWR _7658_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_51 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _5627_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ _7301_/Q _6420_/A _6421_/X _7325_/Q _6608_/X VGND VGND VPWR VPWR _6609_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_84 _6967_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7589_ _7594_/CLK _7589_/D fanout694/X VGND VGND VPWR VPWR _7589_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5725__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6162__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5370__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5658__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput180 _3431_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
Xoutput191 _3421_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3684__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2960 _4391_/X VGND VGND VPWR VPWR hold2960/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2971 _6980_/Q VGND VGND VPWR VPWR _4291_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2982 _6985_/Q VGND VGND VPWR VPWR _4300_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2993 _6982_/Q VGND VGND VPWR VPWR _4294_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6083__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6622__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5291__D1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5189__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6386__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6386__B2 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5043__D1 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4397__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3739__A3 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4105__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3647__C _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6689__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_44_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7573_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3663__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3911__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7541_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6613__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6960_ _6991_/CLK _6960_/D fanout693/X VGND VGND VPWR VPWR _6960_/Q sky130_fd_sc_hd__dfstp_2
X_5911_ _5983_/A _5938_/C _5992_/D VGND VGND VPWR VPWR _5919_/S sky130_fd_sc_hd__and3_4
X_6891_ _7075_/CLK _6891_/D _6841_/X VGND VGND VPWR VPWR _6891_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3978__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5842_ _5842_/A0 _5914_/A1 _5847_/S VGND VGND VPWR VPWR _5842_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5773_ _5773_/A0 _5881_/A1 _5775_/S VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__mux2_1
X_7512_ _7514_/CLK _7512_/D fanout744/X VGND VGND VPWR VPWR _7512_/Q sky130_fd_sc_hd__dfstp_4
X_4724_ _4088_/Y _4558_/X _4726_/A VGND VGND VPWR VPWR _4948_/C sky130_fd_sc_hd__o21a_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6129__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6129__B2 _7520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7443_ _7519_/CLK _7443_/D fanout741/X VGND VGND VPWR VPWR _7443_/Q sky130_fd_sc_hd__dfrtp_4
X_4655_ _4667_/A _4571_/Y _5387_/B _4657_/C _4657_/B VGND VGND VPWR VPWR _5213_/A
+ sky130_fd_sc_hd__o311a_4
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__buf_2
Xhold800 _5756_/X VGND VGND VPWR VPWR _7365_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3606_ _3606_/A _3606_/B _3606_/C _3606_/D VGND VGND VPWR VPWR _3607_/C sky130_fd_sc_hd__nor4_2
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__buf_2
X_7374_ _7579_/CLK hold28/X fanout731/X VGND VGND VPWR VPWR _7374_/Q sky130_fd_sc_hd__dfrtp_4
Xhold811 hold811/A VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ _4675_/A _4675_/B _4586_/C _5089_/B VGND VGND VPWR VPWR _4687_/B sky130_fd_sc_hd__nand4_4
Xinput82 spi_sdoenb VGND VGND VPWR VPWR _4144_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold822 hold822/A VGND VGND VPWR VPWR _7277_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 trap VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__buf_6
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold844 hold844/A VGND VGND VPWR VPWR _7212_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6325_ _7198_/Q _6317_/B _6079_/X _6099_/X _7027_/Q VGND VGND VPWR VPWR _6325_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold855 hold855/A VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3537_ _3682_/A hold32/A _4509_/C VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__and3_4
XFILLER_131_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3902__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold866 hold866/A VGND VGND VPWR VPWR _6966_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4388__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold877 hold877/A VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold888 hold888/A VGND VGND VPWR VPWR _7124_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold899 hold899/A VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6256_ _7533_/Q _6092_/X _6252_/X _6253_/X _6255_/X VGND VGND VPWR VPWR _6257_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6301__B2 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3468_ _4181_/S _3468_/A2 hold341/X _3465_/Y VGND VGND VPWR VPWR _3505_/A sky130_fd_sc_hd__a22o_1
XFILLER_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2201 _7025_/Q VGND VGND VPWR VPWR hold543/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2212 _7294_/Q VGND VGND VPWR VPWR hold559/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4312__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2223 _5610_/X VGND VGND VPWR VPWR hold580/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5207_ _4956_/A _5480_/B2 _4659_/Y VGND VGND VPWR VPWR _5419_/A sky130_fd_sc_hd__a21o_1
Xhold2234 _7333_/Q VGND VGND VPWR VPWR hold671/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6187_ _7490_/Q _6075_/A _6276_/A3 _6100_/X _7474_/Q VGND VGND VPWR VPWR _6187_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout577_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1500 _5609_/X VGND VGND VPWR VPWR hold169/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2245 _7369_/Q VGND VGND VPWR VPWR hold661/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3399_ _6900_/Q VGND VGND VPWR VPWR _3399_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4863__A1 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1511 hold176/X VGND VGND VPWR VPWR _5959_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2256 hold651/X VGND VGND VPWR VPWR _5969_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2267 hold577/X VGND VGND VPWR VPWR _4208_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1522 hold158/X VGND VGND VPWR VPWR _5986_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2278 _5736_/X VGND VGND VPWR VPWR hold598/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1533 hold193/X VGND VGND VPWR VPWR _7436_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5138_ _5138_/A _5138_/B _5138_/C _5138_/D VGND VGND VPWR VPWR _5138_/Y sky130_fd_sc_hd__nand4_1
XANTENNA_clkbuf_leaf_11_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1544 hold145/X VGND VGND VPWR VPWR _7445_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2289 _5802_/X VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1555 hold56/X VGND VGND VPWR VPWR _4258_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6604__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5407__A3 _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1566 _4183_/X VGND VGND VPWR VPWR hold197/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1577 hold94/X VGND VGND VPWR VPWR _7024_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout744_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1588 hold115/X VGND VGND VPWR VPWR _7227_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5069_ _5091_/A _5072_/B _5107_/C VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__and3_4
Xhold1599 hold230/X VGND VGND VPWR VPWR _5932_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3969__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5947__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6368__B2 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1859_A _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6540__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input40_A mgmt_gpio_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4595__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3930__C _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2790 _4453_/X VGND VGND VPWR VPWR hold970/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3658__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3674__A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4440_ _5650_/A1 hold365/X _4168_/D _4422_/S _5956_/C VGND VGND VPWR VPWR _4448_/S
+ sky130_fd_sc_hd__o311a_4
Xhold107 hold107/A VGND VGND VPWR VPWR _7533_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold118 hold118/A VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6531__B2 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold129 hold129/A VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_wire378_A _4145_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4371_ _5912_/A1 _4371_/A1 _4375_/S VGND VGND VPWR VPWR _4371_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3896__A2 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _6110_/A _6121_/A _6144_/B VGND VGND VPWR VPWR _6110_/X sky130_fd_sc_hd__and3_4
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7090_ _7522_/CLK _7090_/D fanout748/X VGND VGND VPWR VPWR _7669_/A sky130_fd_sc_hd__dfrtp_1
Xfanout609 _3408_/Y VGND VGND VPWR VPWR _6067_/A sky130_fd_sc_hd__buf_8
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6295__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6041_ _6429_/C _6067_/B _6040_/Y VGND VGND VPWR VPWR _7593_/D sky130_fd_sc_hd__a21oi_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6943_ _7314_/CLK _6943_/D _4079_/A VGND VGND VPWR VPWR _7649_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__4444__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5270__B2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ _7186_/CLK _6874_/D fanout725/X VGND VGND VPWR VPWR _6874_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3820__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5825_ _5825_/A0 _5969_/A1 hold33/X VGND VGND VPWR VPWR _5825_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5756_ _5756_/A0 _5954_/A1 _5757_/S VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6770__B2 _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4707_ _5091_/C _5387_/C VGND VGND VPWR VPWR _4707_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3584__B2 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5687_ _5894_/A0 _5687_/A1 _5694_/S VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__mux2_1
X_7426_ _7551_/CLK _7426_/D fanout734/X VGND VGND VPWR VPWR _7426_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4638_ _4667_/A _5494_/B2 _4636_/Y VGND VGND VPWR VPWR _4801_/C sky130_fd_sc_hd__o21a_4
Xhold630 hold630/A VGND VGND VPWR VPWR _7537_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7357_ _7421_/CLK _7357_/D fanout715/X VGND VGND VPWR VPWR _7357_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout694_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4569_ _4831_/A _4984_/B _4805_/B VGND VGND VPWR VPWR _4615_/A sky130_fd_sc_hd__and3_2
XFILLER_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold652 _5969_/X VGND VGND VPWR VPWR _7554_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold663 hold663/A VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6308_ _7002_/Q _6097_/B _6120_/B _6332_/C _7032_/Q VGND VGND VPWR VPWR _6308_/X
+ sky130_fd_sc_hd__a32o_1
Xhold674 hold674/A VGND VGND VPWR VPWR _6971_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold685 hold685/A VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7288_ _7329_/CLK _7288_/D fanout704/X VGND VGND VPWR VPWR _7288_/Q sky130_fd_sc_hd__dfstp_4
Xhold696 hold696/A VGND VGND VPWR VPWR _7292_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6239_ _7373_/Q _6084_/X _6276_/A3 _7365_/Q VGND VGND VPWR VPWR _6239_/X sky130_fd_sc_hd__a22o_1
Xhold2020 _4451_/X VGND VGND VPWR VPWR hold460/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2031 _5708_/X VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3639__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2042 hold298/X VGND VGND VPWR VPWR _4538_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2053 _4457_/X VGND VGND VPWR VPWR hold468/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2064 _7384_/Q VGND VGND VPWR VPWR hold501/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1330 _4365_/X VGND VGND VPWR VPWR _7036_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2075 hold513/X VGND VGND VPWR VPWR _5895_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6038__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1341 hold3266/X VGND VGND VPWR VPWR hold3267/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2086 _5766_/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1352 _4293_/A1 VGND VGND VPWR VPWR hold3002/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2097 _7382_/Q VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1363 _4281_/B VGND VGND VPWR VPWR hold3014/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1374 _6783_/A1 VGND VGND VPWR VPWR hold3059/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 _7643_/Q VGND VGND VPWR VPWR _4199_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1396 hold1488/X VGND VGND VPWR VPWR hold1489/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5261__A1 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5677__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4581__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3811__A2 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3478__B _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold3092_A _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6210__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5974__A _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6761__B2 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input88_A spimemio_flash_io1_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3494__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3925__C _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6513__A1 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6513__B2 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6277__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3660__C _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6292__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3669__A _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5587__C _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3940_ _7567_/Q _5983_/A _3637_/C _3501_/X _7575_/Q VGND VGND VPWR VPWR _3940_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3802__A2 _3486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4491__C _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3871_ input47/X _4248_/S _4467_/A _7128_/Q _3870_/X VGND VGND VPWR VPWR _3871_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6201__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5884__A _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5610_ _5610_/A0 _5954_/A1 _5611_/S VGND VGND VPWR VPWR _5610_/X sky130_fd_sc_hd__mux2_1
X_6590_ _7348_/Q _6452_/X _6467_/X _7420_/Q _6589_/X VGND VGND VPWR VPWR _6590_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3566__B2 _7470_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5541_ _4955_/X _5459_/X _5541_/C _5541_/D VGND VGND VPWR VPWR _5543_/B sky130_fd_sc_hd__and4bb_1
X_5472_ _4774_/Y _5471_/X _5386_/X _5256_/X _5267_/X VGND VGND VPWR VPWR _5474_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__6504__B2 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7211_ _7211_/CLK _7211_/D fanout699/X VGND VGND VPWR VPWR _7211_/Q sky130_fd_sc_hd__dfstp_1
X_4423_ _4423_/A0 _4422_/X _4423_/S VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5823__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2624_A _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7142_ _7266_/CLK _7142_/D fanout692/X VGND VGND VPWR VPWR _7142_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_125_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4354_ _4354_/A0 _4547_/A0 _4357_/S VGND VGND VPWR VPWR _4354_/X sky130_fd_sc_hd__mux2_1
Xfanout406 hold125/X VGND VGND VPWR VPWR _5619_/A sky130_fd_sc_hd__buf_6
XFILLER_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout417 _5740_/A VGND VGND VPWR VPWR _4473_/A sky130_fd_sc_hd__buf_6
Xfanout428 _4689_/Y VGND VGND VPWR VPWR _4997_/B sky130_fd_sc_hd__buf_8
X_7073_ _4127_/A1 _7073_/D _6863_/X VGND VGND VPWR VPWR _7073_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout439 _3502_/X VGND VGND VPWR VPWR _4388_/B sky130_fd_sc_hd__buf_12
X_4285_ _4289_/S _4285_/B VGND VGND VPWR VPWR _4285_/Y sky130_fd_sc_hd__nand2_1
X_6024_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6121_/A sky130_fd_sc_hd__and2_4
XFILLER_140_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6926_ _7264_/CLK _6926_/D fanout688/X VGND VGND VPWR VPWR _6926_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6857_ _6861_/A _6869_/B VGND VGND VPWR VPWR _6857_/X sky130_fd_sc_hd__and2_1
XANTENNA__5794__A _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5808_ _5808_/A0 _5952_/A1 _5811_/S VGND VGND VPWR VPWR _5808_/X sky130_fd_sc_hd__mux2_1
X_6788_ _6792_/S _6788_/B VGND VGND VPWR VPWR _6788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ _5739_/A0 _5955_/A1 _5739_/S VGND VGND VPWR VPWR _5739_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4203__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7409_ _7497_/CLK _7409_/D fanout709/X VGND VGND VPWR VPWR _7409_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold460 hold460/A VGND VGND VPWR VPWR _7113_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold487_A hold487/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold482 hold482/A VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4857__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold493 hold493/A VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5034__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input142_A wb_dat_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6274__A3 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1160 hold2839/X VGND VGND VPWR VPWR hold2840/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1171 hold2850/X VGND VGND VPWR VPWR hold2851/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1182 hold3228/X VGND VGND VPWR VPWR hold3229/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold3105_A _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 hold2853/X VGND VGND VPWR VPWR hold2854/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__B2 _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5908__S hold42/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6734__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3655__C _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_2__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4150_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3671__B _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4070_ hold9/A hold15/A _4074_/S VGND VGND VPWR VPWR _6888_/D sky130_fd_sc_hd__mux2_1
XFILLER_95_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_58_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4972_ _5113_/A _5089_/D _5399_/C _5282_/C VGND VGND VPWR VPWR _5324_/A sky130_fd_sc_hd__o211a_2
XANTENNA__3787__A1 _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6711_ _7149_/Q _6408_/A _6424_/X _7129_/Q _6702_/X VGND VGND VPWR VPWR _6711_/X
+ sky130_fd_sc_hd__a221o_1
X_3923_ _3997_/A1 _3922_/Y _3923_/S VGND VGND VPWR VPWR _3923_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5818__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2574_A _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6642_ _7486_/Q _6447_/C _6428_/X _6419_/C _7566_/Q VGND VGND VPWR VPWR _6642_/X
+ sky130_fd_sc_hd__a32o_1
X_3854_ _3854_/A _3854_/B _3854_/C _3854_/D VGND VGND VPWR VPWR _3855_/C sky130_fd_sc_hd__and4_1
XFILLER_177_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6573_ _6572_/X _6598_/A2 _6573_/S VGND VGND VPWR VPWR _7619_/D sky130_fd_sc_hd__mux2_1
X_3785_ _7180_/Q _4376_/B _3738_/B _3675_/X _7190_/Q VGND VGND VPWR VPWR _3785_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3565__C _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ _5059_/A _5282_/B _5524_/A3 _5559_/C _5523_/X VGND VGND VPWR VPWR _5524_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_145_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6489__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5455_ _4947_/Y _5245_/X _5366_/X VGND VGND VPWR VPWR _5543_/A sky130_fd_sc_hd__o21ba_1
X_4406_ _5650_/A1 hold365/X _4168_/D _4422_/S VGND VGND VPWR VPWR _4406_/Y sky130_fd_sc_hd__o31ai_2
X_5386_ _5480_/A1 _5509_/A3 _4716_/Y _5563_/A1 VGND VGND VPWR VPWR _5386_/X sky130_fd_sc_hd__a211o_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3711__A1 input24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7125_ _7186_/CLK _7125_/D fanout726/X VGND VGND VPWR VPWR _7125_/Q sky130_fd_sc_hd__dfrtp_4
X_4337_ _4337_/A0 _4548_/A0 _4339_/S VGND VGND VPWR VPWR _4337_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout392_A _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7056_ _7160_/CLK _7056_/D fanout700/X VGND VGND VPWR VPWR _7056_/Q sky130_fd_sc_hd__dfrtp_4
X_4268_ _4268_/A0 _4548_/A0 _4270_/S VGND VGND VPWR VPWR _4268_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6007_ _6932_/Q _6009_/B _6019_/A _7584_/Q _4117_/Y VGND VGND VPWR VPWR _6017_/D
+ sky130_fd_sc_hd__o311a_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6661__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4199_ _4199_/A0 _4199_/A1 _4429_/B VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout657_A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6116__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _4127_/A1 _6909_/D _6859_/X VGND VGND VPWR VPWR _6909_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5728__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5519__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6413__A _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6192__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5029__A _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10__f_wb_clk_i clkbuf_3_5_0_wb_clk_i/X VGND VGND VPWR VPWR _7636_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold290 hold290/A VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout770 _4844_/B VGND VGND VPWR VPWR _4945_/A sky130_fd_sc_hd__buf_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6652__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5207__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__A1 input29/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__B2 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__C1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3666__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6042__B _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4194__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3570_ _3491_/X _3570_/B _3570_/C VGND VGND VPWR VPWR _3570_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__3682__A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5240_ _5091_/A _5072_/B wire649/X _5282_/A VGND VGND VPWR VPWR _5243_/C sky130_fd_sc_hd__a22o_2
XANTENNA__6486__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3309 _7107_/Q VGND VGND VPWR VPWR _4171_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4497__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2608 _7389_/Q VGND VGND VPWR VPWR hold899/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5171_ _5038_/A _5038_/B _5180_/A _5038_/C _4928_/B VGND VGND VPWR VPWR _5171_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2619 _7149_/Q VGND VGND VPWR VPWR hold933/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4122_ _6909_/Q _4076_/C _4121_/Y _4058_/B _4010_/Y VGND VGND VPWR VPWR _7074_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1907 hold296/X VGND VGND VPWR VPWR _4507_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3733__A_N _3686_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5105__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1918 hold265/X VGND VGND VPWR VPWR _5655_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6643__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1929 hold338/X VGND VGND VPWR VPWR _4379_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ _3998_/Y _4123_/B _4052_/X _4053_/B2 _4062_/A VGND VGND VPWR VPWR _6895_/D
+ sky130_fd_sc_hd__o221a_1
Xinput3 debug_out VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_2
XFILLER_25_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4955_ _5248_/A _5248_/B _5089_/D _4953_/X _5222_/A VGND VGND VPWR VPWR _4955_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3906_ input15/X _3503_/X _3666_/X _7012_/Q _3905_/X VGND VGND VPWR VPWR _3913_/A
+ sky130_fd_sc_hd__a221o_1
X_4886_ _5222_/A _5065_/A VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_177_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6625_ _6624_/X _6649_/A1 _6777_/S VGND VGND VPWR VPWR _6625_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3837_ _3837_/A _3837_/B _3837_/C _3837_/D VGND VGND VPWR VPWR _3854_/B sky130_fd_sc_hd__nor4_1
XANTENNA__6174__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6556_ _7355_/Q _6459_/B _6428_/X _6420_/C _7395_/Q VGND VGND VPWR VPWR _6556_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout405_A _3492_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3768_ _7418_/Q _4551_/B _5956_/B _3669_/X _6970_/Q VGND VGND VPWR VPWR _3768_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5507_ _4716_/Y _5065_/Y _5210_/X _5185_/C _5355_/A VGND VGND VPWR VPWR _5508_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3932__B2 _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6487_ _7296_/Q _6420_/A _6467_/X _7416_/Q _6486_/X VGND VGND VPWR VPWR _6494_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3699_ _7355_/Q _5740_/A _5956_/B _3498_/X _7379_/Q VGND VGND VPWR VPWR _3699_/X
+ sky130_fd_sc_hd__a32o_1
X_5438_ _5438_/A _5438_/B _5438_/C _5438_/D VGND VGND VPWR VPWR _5441_/C sky130_fd_sc_hd__and4_1
XFILLER_105_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput340 hold1072/X VGND VGND VPWR VPWR hold1073/A sky130_fd_sc_hd__buf_6
XFILLER_160_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5685__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout774_A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5369_ _4601_/Y _4956_/A _4956_/B _4960_/B VGND VGND VPWR VPWR _5457_/B sky130_fd_sc_hd__a31o_1
XFILLER_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ _7641_/CLK _7108_/D fanout751/X VGND VGND VPWR VPWR _7108_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6634__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ _7164_/CLK _7039_/D fanout698/X VGND VGND VPWR VPWR _7039_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6408__A _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A wb_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3620__B1 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3486__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input70_A mgmt_gpio_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3923__A1 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6322__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3687__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5222__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6640__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6752__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5600__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4740_ _4786_/D _4805_/B _4831_/C _4767_/A VGND VGND VPWR VPWR _5077_/B sky130_fd_sc_hd__and4bb_4
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__B1 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4671_ _4667_/A _4667_/B _4667_/C _4974_/D _4974_/B VGND VGND VPWR VPWR _5063_/D
+ sky130_fd_sc_hd__o311a_2
X_6410_ _7594_/Q _6455_/B _6462_/C VGND VGND VPWR VPWR _6410_/X sky130_fd_sc_hd__and3_1
X_3622_ _7234_/Q _3617_/X _3618_/X _3616_/X _3621_/X VGND VGND VPWR VPWR _3623_/D
+ sky130_fd_sc_hd__a2111o_4
XFILLER_190_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7390_ _7579_/CLK hold21/X fanout731/X VGND VGND VPWR VPWR _7390_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6341_ _6332_/B _6333_/X _6340_/X _6339_/X VGND VGND VPWR VPWR _6341_/X sky130_fd_sc_hd__a211o_1
X_3553_ _5938_/A _5938_/B _5992_/C VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__and3_4
XFILLER_127_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2537_A _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6272_ _7358_/Q _6099_/X _6112_/X _7486_/Q _6271_/X VGND VGND VPWR VPWR _6272_/X
+ sky130_fd_sc_hd__a221o_1
X_3484_ _3507_/A hold38/X _5830_/C VGND VGND VPWR VPWR _3484_/X sky130_fd_sc_hd__and3_2
Xhold3106 hold3106/A VGND VGND VPWR VPWR _4474_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5667__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3117 _6967_/Q VGND VGND VPWR VPWR hold3117/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5223_ _5223_/A _5223_/B _5223_/C _5223_/D VGND VGND VPWR VPWR _5224_/C sky130_fd_sc_hd__nand4_1
XFILLER_170_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3128 hold3128/A VGND VGND VPWR VPWR _4353_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3139 hold3139/A VGND VGND VPWR VPWR _4359_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2405 _7418_/Q VGND VGND VPWR VPWR hold681/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5831__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2416 _5584_/X VGND VGND VPWR VPWR hold856/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2427 hold687/X VGND VGND VPWR VPWR _4345_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5154_ _4687_/Y _4793_/Y _4821_/Y _4796_/Y _4723_/Y VGND VGND VPWR VPWR _5156_/B
+ sky130_fd_sc_hd__o32a_1
Xhold2438 _7478_/Q VGND VGND VPWR VPWR hold723/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1704 _5923_/X VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2449 _7317_/Q VGND VGND VPWR VPWR hold879/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6616__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1715 hold334/X VGND VGND VPWR VPWR _5958_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4105_ _6427_/A _4105_/B VGND VGND VPWR VPWR _4105_/Y sky130_fd_sc_hd__nand2_1
Xhold1726 _7280_/Q VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3693__A3 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1737 _4442_/X VGND VGND VPWR VPWR hold356/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5085_ _4600_/Y _5387_/C _4717_/B _5084_/Y VGND VGND VPWR VPWR _5085_/Y sky130_fd_sc_hd__a31oi_1
Xhold1748 hold293/X VGND VGND VPWR VPWR _7004_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1759 hold274/X VGND VGND VPWR VPWR _5951_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4036_ _4036_/A0 _4035_/X _4040_/A VGND VGND VPWR VPWR _6903_/D sky130_fd_sc_hd__mux2_1
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3850__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4690__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _5987_/A0 _5996_/A1 _5991_/S VGND VGND VPWR VPWR _5987_/X sky130_fd_sc_hd__mux2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4938_ _4882_/Y _4936_/Y _4937_/Y _4934_/Y VGND VGND VPWR VPWR _4941_/C sky130_fd_sc_hd__o211ai_1
XANTENNA__3602__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _4646_/A _4608_/Y _4617_/Y _4860_/B VGND VGND VPWR VPWR _4889_/B sky130_fd_sc_hd__o211ai_4
X_7657_ _7657_/A VGND VGND VPWR VPWR _7657_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_41 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_63 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4158__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6608_ _7389_/Q _6413_/C _6426_/X _6451_/X _7485_/Q VGND VGND VPWR VPWR _6608_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_74 _4179_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7588_ _7610_/CLK _7588_/D fanout692/X VGND VGND VPWR VPWR _7588_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_85 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3905__A1 _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6539_ _7546_/Q _6419_/A _6435_/X _7514_/Q _6538_/X VGND VGND VPWR VPWR _6544_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_180_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4849__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5741__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput181 _3430_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 _3420_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XANTENNA__4330__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2950 _7179_/Q VGND VGND VPWR VPWR hold2950/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6607__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3684__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2961 _7038_/Q VGND VGND VPWR VPWR hold2961/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2972 hold2972/A VGND VGND VPWR VPWR hold2972/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2983 hold2983/A VGND VGND VPWR VPWR hold2983/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2994 hold2994/A VGND VGND VPWR VPWR hold2994/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6083__B2 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6386__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3497__A hold40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4105__B _4105_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6138__A2 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4149__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output274_A _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3663__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4775__B _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4267__S _4270_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4085__B1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6898__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5910_ hold20/X _5910_/A1 hold42/X VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__mux2_1
X_6890_ _7075_/CLK _6890_/D _6840_/X VGND VGND VPWR VPWR _6890_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3832__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ _5841_/A0 _5922_/A0 _5847_/S VGND VGND VPWR VPWR _5841_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5585__A0 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5772_ _5772_/A0 _5997_/A1 _5775_/S VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4723_ _5068_/B _5059_/B VGND VGND VPWR VPWR _4723_/Y sky130_fd_sc_hd__nand2_4
X_7511_ _7531_/CLK _7511_/D fanout743/X VGND VGND VPWR VPWR _7511_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_159_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6129__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5826__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7442_ _7514_/CLK _7442_/D fanout744/X VGND VGND VPWR VPWR _7442_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4654_ _4644_/Y _4646_/Y _4833_/A VGND VGND VPWR VPWR _4654_/Y sky130_fd_sc_hd__o21ai_4
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__buf_4
X_3605_ input9/X _3486_/X _3508_/X _7557_/Q _3604_/X VGND VGND VPWR VPWR _3606_/D
+ sky130_fd_sc_hd__a221o_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__buf_2
X_7373_ _7478_/CLK _7373_/D fanout715/X VGND VGND VPWR VPWR _7373_/Q sky130_fd_sc_hd__dfrtp_2
X_4585_ _4585_/A _4643_/C _4823_/D _5089_/B VGND VGND VPWR VPWR _4585_/Y sky130_fd_sc_hd__nand4_2
Xhold801 hold801/A VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold812 _5880_/X VGND VGND VPWR VPWR _7475_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold823 hold823/A VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__clkbuf_4
Xhold834 hold834/A VGND VGND VPWR VPWR _7199_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2919_A _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput94 uart_enabled VGND VGND VPWR VPWR _4173_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_6324_ _7007_/Q _6082_/X _6094_/X _7210_/Q _6323_/X VGND VGND VPWR VPWR _6327_/C
+ sky130_fd_sc_hd__a221o_1
X_3536_ _7494_/Q _5938_/C _5965_/B _3535_/X _7486_/Q VGND VGND VPWR VPWR _3536_/X
+ sky130_fd_sc_hd__a32o_1
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold856 hold856/A VGND VGND VPWR VPWR _7211_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold867 hold867/A VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold878 hold878/A VGND VGND VPWR VPWR _7012_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6255_ _7325_/Q _6082_/X _6110_/X _7437_/Q _6254_/X VGND VGND VPWR VPWR _6255_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_89_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold889 hold889/A VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3467_ _4181_/S _3468_/A2 _3466_/X _3465_/Y VGND VGND VPWR VPWR _3467_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_107_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2202 hold543/X VGND VGND VPWR VPWR _4351_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5206_ _5202_/X _5204_/X _5205_/X VGND VGND VPWR VPWR _5206_/Y sky130_fd_sc_hd__a21oi_1
Xhold2213 hold559/X VGND VGND VPWR VPWR _5676_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2224 _7305_/Q VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6186_ _7498_/Q _6085_/X _6112_/X _7482_/Q _6185_/X VGND VGND VPWR VPWR _6186_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2235 hold671/X VGND VGND VPWR VPWR _5720_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1501 hold169/X VGND VGND VPWR VPWR _7240_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2246 hold661/X VGND VGND VPWR VPWR _5761_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1512 _5959_/X VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5137_ _4695_/Y _4735_/Y _4821_/Y _4687_/Y VGND VGND VPWR VPWR _5139_/C sky130_fd_sc_hd__a211o_1
Xhold2257 _7254_/Q VGND VGND VPWR VPWR hold587/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2268 _7546_/Q VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1523 _5986_/X VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2279 _7284_/Q VGND VGND VPWR VPWR hold801/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1534 _7548_/Q VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1545 _7532_/Q VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1556 _4258_/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1567 hold197/X VGND VGND VPWR VPWR hold1567/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5068_ _5091_/C _5068_/B _5453_/C VGND VGND VPWR VPWR _5573_/D sky130_fd_sc_hd__nand3_1
XANTENNA__6604__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1578 _7500_/Q VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1589 _7565_/Q VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_38_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4019_ _4040_/D _4014_/B _3450_/X _4017_/Y VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6368__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4379__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6540__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3135_A _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input33_A mask_rev_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3930__D _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2780 hold815/X VGND VGND VPWR VPWR _5862_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2791 _6920_/Q VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6359__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3658__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5646__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3593__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3674__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6050__B _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold108 hold108/A VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6531__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold119 hold119/A VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4370_ _4370_/A _4551_/D VGND VGND VPWR VPWR _4375_/S sky130_fd_sc_hd__nand2_4
XFILLER_171_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6040_ _6429_/C _6067_/B _6929_/Q VGND VGND VPWR VPWR _6040_/Y sky130_fd_sc_hd__nor3_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ _7306_/CLK _6942_/D _4079_/A VGND VGND VPWR VPWR _6942_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6873_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6873_/X sky130_fd_sc_hd__and2_1
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3820__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2869_A _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ _5824_/A0 _5968_/A1 hold33/X VGND VGND VPWR VPWR _5824_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5755_ _5755_/A0 _5953_/A1 _5757_/S VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6770__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3584__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4706_ _4706_/A _5107_/C VGND VGND VPWR VPWR _4706_/Y sky130_fd_sc_hd__nand2_4
X_5686_ _5686_/A _5947_/C VGND VGND VPWR VPWR _5694_/S sky130_fd_sc_hd__nand2_8
X_7425_ _7489_/CLK _7425_/D fanout719/X VGND VGND VPWR VPWR _7425_/Q sky130_fd_sc_hd__dfrtp_2
X_4637_ _4772_/A _4814_/C VGND VGND VPWR VPWR _4836_/C sky130_fd_sc_hd__nor2_8
XFILLER_190_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold620 _5771_/X VGND VGND VPWR VPWR _7378_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold631 hold631/A VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7356_ _7421_/CLK _7356_/D fanout715/X VGND VGND VPWR VPWR _7356_/Q sky130_fd_sc_hd__dfrtp_4
X_4568_ _4831_/A _4984_/B VGND VGND VPWR VPWR _4568_/Y sky130_fd_sc_hd__nand2_4
Xhold642 hold642/A VGND VGND VPWR VPWR _7546_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold653 hold653/A VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6307_ _6306_/X _6330_/A2 _6777_/S VGND VGND VPWR VPWR _6307_/X sky130_fd_sc_hd__mux2_1
X_3519_ hold40/A _5965_/A _5596_/B VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__and3_2
Xhold664 hold664/A VGND VGND VPWR VPWR _7191_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7287_ _7327_/CLK _7287_/D fanout703/X VGND VGND VPWR VPWR _7287_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_103_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold675 hold675/A VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold686 hold686/A VGND VGND VPWR VPWR _7434_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4499_ _4553_/A0 _4499_/A1 _4502_/S VGND VGND VPWR VPWR _4499_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout687_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold697 hold697/A VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6238_ _6260_/A2 _4116_/X _6067_/X _6237_/X VGND VGND VPWR VPWR _7607_/D sky130_fd_sc_hd__o31a_1
Xhold2010 _7393_/Q VGND VGND VPWR VPWR hold455/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2021 _7561_/Q VGND VGND VPWR VPWR hold419/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2032 _7312_/Q VGND VGND VPWR VPWR hold497/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2043 _7427_/Q VGND VGND VPWR VPWR hold330/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6649_/S _6169_/A2 _6573_/S _6168_/X VGND VGND VPWR VPWR _6169_/X sky130_fd_sc_hd__a211o_1
XFILLER_134_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2054 _7153_/Q VGND VGND VPWR VPWR hold479/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1320 hold3176/X VGND VGND VPWR VPWR _7209_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2065 hold501/X VGND VGND VPWR VPWR _5778_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1502_A _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1331 hold3159/X VGND VGND VPWR VPWR hold3160/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2076 _7472_/Q VGND VGND VPWR VPWR hold517/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6119__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1342 _5795_/X VGND VGND VPWR VPWR _7399_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2087 _7454_/Q VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1353 _4301_/A1 VGND VGND VPWR VPWR hold3000/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2098 hold50/X VGND VGND VPWR VPWR _5775_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_27_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1364 _4289_/A1 VGND VGND VPWR VPWR hold2964/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6589__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1375 _6784_/B VGND VGND VPWR VPWR hold3054/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1386 hold2095/X VGND VGND VPWR VPWR hold2096/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__A0 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1397 _7641_/Q VGND VGND VPWR VPWR _4189_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7556_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1871_A _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3811__A3 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3478__C _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7365_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6761__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3575__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3494__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3925__D _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6513__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5721__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4524__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4742__A_N _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6277__A1 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6277__B2 _7446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4288__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6682__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output237_A _4148_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4772__C _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3669__B _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5587__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4491__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3870_ _7138_/Q _3637_/C _3576_/X _5974_/A _7560_/Q VGND VGND VPWR VPWR _3870_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6201__A1 _7451_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5884__B _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4280__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3566__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5540_ _4953_/X _4956_/Y _5248_/X _5371_/X _4959_/X VGND VGND VPWR VPWR _5541_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_54_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5471_ _4879_/D _4747_/B _5073_/A _4748_/Y VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__o31a_2
XANTENNA__6504__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4422_ _4448_/A0 _4422_/A1 _4422_/S VGND VGND VPWR VPWR _4422_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5712__A0 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7210_ _7210_/CLK _7210_/D fanout702/X VGND VGND VPWR VPWR _7210_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7141_ _7197_/CLK _7141_/D fanout728/X VGND VGND VPWR VPWR _7141_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold41_A hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4353_ _4353_/A0 _5876_/A1 _4357_/S VGND VGND VPWR VPWR _4353_/X sky130_fd_sc_hd__mux2_1
Xfanout407 _3598_/B VGND VGND VPWR VPWR _5612_/B sky130_fd_sc_hd__buf_8
XANTENNA__6000__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout418 hold47/X VGND VGND VPWR VPWR _5740_/A sky130_fd_sc_hd__buf_8
X_7072_ _7075_/CLK _7072_/D _6862_/X VGND VGND VPWR VPWR _7072_/Q sky130_fd_sc_hd__dfrtp_1
X_4284_ _4289_/S _3795_/B _4283_/Y VGND VGND VPWR VPWR _6975_/D sky130_fd_sc_hd__o21ai_1
Xfanout429 _5342_/A VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__buf_8
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6023_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6089_/C sky130_fd_sc_hd__nor2_8
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6881__D _6881_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5779__A0 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6925_ _7264_/CLK _6925_/D fanout688/X VGND VGND VPWR VPWR _6925_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_81_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6856_ _6861_/A _6869_/B VGND VGND VPWR VPWR _6856_/X sky130_fd_sc_hd__and2_1
XFILLER_80_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5794__B _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5807_ _5807_/A0 _5951_/A1 _5811_/S VGND VGND VPWR VPWR _5807_/X sky130_fd_sc_hd__mux2_1
X_3999_ _4058_/A _4058_/B _7073_/Q _6908_/Q VGND VGND VPWR VPWR _4006_/A sky130_fd_sc_hd__o31a_2
XANTENNA__6743__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6787_ _6792_/S _3795_/B _6786_/Y VGND VGND VPWR VPWR _7632_/D sky130_fd_sc_hd__o21ai_1
X_5738_ _5738_/A0 _5954_/A1 _5739_/S VGND VGND VPWR VPWR _5738_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4203__B _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5669_ hold487/X _5669_/A1 _5676_/S VGND VGND VPWR VPWR _5669_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7408_ _7497_/CLK _7408_/D fanout707/X VGND VGND VPWR VPWR _7408_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_191_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold450 _5968_/X VGND VGND VPWR VPWR _7553_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7339_ _7537_/CLK _7339_/D fanout707/X VGND VGND VPWR VPWR _7339_/Q sky130_fd_sc_hd__dfrtp_4
Xhold461 hold461/A VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold472 hold472/A VGND VGND VPWR VPWR _7128_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold483 hold483/A VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold494 hold494/A VGND VGND VPWR VPWR _6938_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input135_A wb_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1150 hold3091/X VGND VGND VPWR VPWR hold1150/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1161 hold2841/X VGND VGND VPWR VPWR _7417_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1172 hold2852/X VGND VGND VPWR VPWR _7023_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1183 hold3220/X VGND VGND VPWR VPWR hold1183/X sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1194 _4194_/X VGND VGND VPWR VPWR _6913_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5050__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6734__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_690 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3671__C _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3720__A2 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4971_ _4571_/Y _4843_/A _4709_/Y VGND VGND VPWR VPWR _4971_/X sky130_fd_sc_hd__o21a_4
XFILLER_91_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6710_ _7018_/Q _6425_/X _6454_/X _7068_/Q _6709_/X VGND VGND VPWR VPWR _6710_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3787__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3922_ _3922_/A _3922_/B _3922_/C VGND VGND VPWR VPWR _3922_/Y sky130_fd_sc_hd__nand3_4
X_3853_ _7023_/Q _3667_/X _3849_/X _3850_/X _3852_/X VGND VGND VPWR VPWR _3854_/D
+ sky130_fd_sc_hd__a2111oi_2
X_6641_ _7326_/Q _6421_/X _6462_/X _7366_/Q _6640_/X VGND VGND VPWR VPWR _6647_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6186__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3619__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5528__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3539__A2 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6572_ _6649_/S _6572_/A2 _6570_/Y _6571_/X VGND VGND VPWR VPWR _6572_/X sky130_fd_sc_hd__a22o_1
X_3784_ _7538_/Q _3590_/C _5938_/C _3565_/X _7466_/Q VGND VGND VPWR VPWR _3792_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3944__C1 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5523_ _5282_/B _5399_/C _5399_/D _5324_/A VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__a31o_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5834__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ _5180_/B _4935_/X _5238_/X _5453_/X _5347_/X VGND VGND VPWR VPWR _5545_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_173_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3862__B _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4405_ _4405_/A0 _4544_/A1 _4405_/S VGND VGND VPWR VPWR _4405_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5161__A1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5385_ _4600_/Y _4810_/C _4743_/Y _5067_/C _5086_/B VGND VGND VPWR VPWR _5385_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_114_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3711__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4336_ _4336_/A0 _4547_/A0 _4339_/S VGND VGND VPWR VPWR _4336_/X sky130_fd_sc_hd__mux2_1
X_7124_ _7186_/CLK _7124_/D fanout726/X VGND VGND VPWR VPWR _7124_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_87_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7055_ _7176_/CLK _7055_/D fanout723/X VGND VGND VPWR VPWR _7055_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4267_ _4267_/A0 _4547_/A0 _4270_/S VGND VGND VPWR VPWR _4267_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout385_A _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6006_ _6006_/A _7584_/Q VGND VGND VPWR VPWR _6006_/X sky130_fd_sc_hd__and2_1
XFILLER_28_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4198_ hold142/X _5627_/A1 _4202_/S VGND VGND VPWR VPWR _4198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3475__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ _7075_/CLK _6908_/D _6858_/X VGND VGND VPWR VPWR _6908_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3778__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6839_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6839_/X sky130_fd_sc_hd__and2_1
XANTENNA__6177__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6716__A2 _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire649 _4856_/Y VGND VGND VPWR VPWR wire649/X sky130_fd_sc_hd__buf_2
XFILLER_109_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5744__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1834_A _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3950__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold291 hold291/A VGND VGND VPWR VPWR _7195_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3702__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6101__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout760 _4831_/C VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__buf_12
Xfanout771 input121/X VGND VGND VPWR VPWR _4844_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_93_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6652__A1 _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6652__B2 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5207__A2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3769__A2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6707__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3666__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5391__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3941__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3682__B _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6340__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5170_ _5339_/D _5180_/B _5030_/C _5039_/B VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__a31o_1
Xhold2609 hold899/X VGND VGND VPWR VPWR _5783_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4121_ _4121_/A _6882_/Q VGND VGND VPWR VPWR _4121_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1908 _4507_/X VGND VGND VPWR VPWR hold297/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1919 _5655_/X VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_717 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4052_ _4058_/A _4058_/B _7073_/Q _6893_/Q VGND VGND VPWR VPWR _4052_/X sky130_fd_sc_hd__o31a_1
XANTENNA__6643__B2 _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3457__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4406__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5829__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4954_ _4954_/A _5248_/A _4954_/C VGND VGND VPWR VPWR _4960_/B sky130_fd_sc_hd__nand3_4
XFILLER_33_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3905_ _7158_/Q _5947_/B _3514_/X _3544_/X _7416_/Q VGND VGND VPWR VPWR _3905_/X
+ sky130_fd_sc_hd__a32o_1
X_7673_ _7673_/A VGND VGND VPWR VPWR _7673_/X sky130_fd_sc_hd__clkbuf_2
X_4885_ _5222_/A _4942_/A _4948_/C VGND VGND VPWR VPWR _4885_/X sky130_fd_sc_hd__and3_2
XFILLER_177_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6624_ _6649_/S _7620_/Q _6622_/X _6623_/X VGND VGND VPWR VPWR _6624_/X sky130_fd_sc_hd__a22o_1
X_3836_ _7237_/Q _3515_/X _4394_/A _7063_/Q _3835_/X VGND VGND VPWR VPWR _3837_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5382__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3767_ _7330_/Q _5713_/A _3562_/X _7298_/Q _3766_/X VGND VGND VPWR VPWR _3767_/X
+ sky130_fd_sc_hd__a221o_1
X_6555_ _7435_/Q _6747_/B _6747_/C _6460_/X _7387_/Q VGND VGND VPWR VPWR _6555_/X
+ sky130_fd_sc_hd__a32o_1
X_5506_ _5205_/X _5506_/B _5506_/C _5506_/D VGND VGND VPWR VPWR _5550_/C sky130_fd_sc_hd__and4b_1
XANTENNA__3932__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6486_ _7368_/Q _6413_/C _6651_/C _6422_/X _7288_/Q VGND VGND VPWR VPWR _6486_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_133_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3698_ _7395_/Q _3473_/X _4533_/A _7186_/Q _3697_/X VGND VGND VPWR VPWR _3698_/X
+ sky130_fd_sc_hd__a221o_1
X_5437_ _5183_/B _5329_/X _5436_/X VGND VGND VPWR VPWR _5438_/D sky130_fd_sc_hd__a21oi_2
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput330 hold1115/X VGND VGND VPWR VPWR hold1116/A sky130_fd_sc_hd__buf_6
Xoutput341 hold1062/X VGND VGND VPWR VPWR hold1063/A sky130_fd_sc_hd__buf_6
XFILLER_161_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5368_ _4654_/Y _4936_/Y _5245_/X _5419_/A VGND VGND VPWR VPWR _5512_/A sky130_fd_sc_hd__o31a_2
XFILLER_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7107_ _7646_/CLK _7107_/D fanout751/X VGND VGND VPWR VPWR _7107_/Q sky130_fd_sc_hd__dfrtp_4
X_4319_ _3643_/Y _4319_/A1 _4321_/S VGND VGND VPWR VPWR _6998_/D sky130_fd_sc_hd__mux2_1
X_5299_ _4705_/Y _4722_/Y _4737_/Y _4746_/Y _5298_/X VGND VGND VPWR VPWR _5538_/A
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6229__A4 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6634__A1 _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7038_ _7179_/CLK _7038_/D fanout698/X VGND VGND VPWR VPWR _7038_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6408__B _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3853__D1 _3852_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4660__A3 _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1784_A _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__B1 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3620__A1 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3486__C _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6165__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire424 _4696_/B VGND VGND VPWR VPWR _4850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold3165_A _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input63_A mgmt_gpio_in[34] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6322__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout590 hold487/X VGND VGND VPWR VPWR _5975_/A0 sky130_fd_sc_hd__clkbuf_8
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5649__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4780__C _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4670_ _4568_/Y _4984_/C _4860_/A VGND VGND VPWR VPWR _4974_/D sky130_fd_sc_hd__o21ai_4
XFILLER_159_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3621_ _7404_/Q _5794_/A _3542_/X _6924_/Q _3620_/X VGND VGND VPWR VPWR _3621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_186_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5364__A1 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6561__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3552_ _5722_/B _5612_/C _5614_/B VGND VGND VPWR VPWR _3552_/X sky130_fd_sc_hd__and3_4
X_6340_ _7179_/Q _6092_/X _6119_/X _7134_/Q _6334_/X VGND VGND VPWR VPWR _6340_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3914__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6271_ _7430_/Q _6080_/A _6074_/X _6120_/X _7342_/Q VGND VGND VPWR VPWR _6271_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5116__A1 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6313__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3483_ _3504_/A _3504_/B VGND VGND VPWR VPWR _3483_/X sky130_fd_sc_hd__and2b_2
XANTENNA__5116__B2 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5222_ _5222_/A _5222_/B _5222_/C _5387_/D VGND VGND VPWR VPWR _5223_/C sky130_fd_sc_hd__nand4_2
XFILLER_103_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3107 _4474_/X VGND VGND VPWR VPWR hold3107/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3118 hold3118/A VGND VGND VPWR VPWR _4272_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3129 _4353_/X VGND VGND VPWR VPWR hold3129/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2406 hold681/X VGND VGND VPWR VPWR _5816_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2417 _7507_/Q VGND VGND VPWR VPWR hold655/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5153_ _5153_/A _5153_/B _5153_/C VGND VGND VPWR VPWR _5156_/A sky130_fd_sc_hd__and3_1
Xhold2428 _4345_/X VGND VGND VPWR VPWR hold688/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2439 hold723/X VGND VGND VPWR VPWR _5883_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1705 _7496_/Q VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4104_ _6429_/C _6441_/D _6433_/D _7594_/Q VGND VGND VPWR VPWR _4105_/B sky130_fd_sc_hd__and4bb_4
XANTENNA__6616__A1 _7445_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1716 _5958_/X VGND VGND VPWR VPWR hold335/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5084_ _5084_/A _5467_/A _5084_/C _5084_/D VGND VGND VPWR VPWR _5084_/Y sky130_fd_sc_hd__nand4_1
Xhold1727 hold387/X VGND VGND VPWR VPWR _5661_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1738 _7009_/Q VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1749 _7394_/Q VGND VGND VPWR VPWR hold150/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4035_ _6902_/Q _4007_/B _4025_/Y _4034_/X VGND VGND VPWR VPWR _4035_/X sky130_fd_sc_hd__a22o_1
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _5986_/A0 _5986_/A1 _5991_/S VGND VGND VPWR VPWR _5986_/X sky130_fd_sc_hd__mux2_1
XFILLER_169_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6395__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_820 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4937_ _4954_/A _5453_/A _4970_/C _4940_/D VGND VGND VPWR VPWR _4937_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3602__B2 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _6516_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7656_ _7656_/A VGND VGND VPWR VPWR _7656_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_31 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _4571_/Y _4646_/A _5387_/B _4617_/Y _4860_/B VGND VGND VPWR VPWR _5213_/C
+ sky130_fd_sc_hd__o311a_2
XANTENNA_42 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4158__A2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ _7357_/Q _6413_/C _6459_/C _6408_/B _7381_/Q VGND VGND VPWR VPWR _6607_/X
+ sky130_fd_sc_hd__a32o_1
X_3819_ _7497_/Q hold41/A _3812_/X _3813_/X _3818_/X VGND VGND VPWR VPWR _3819_/Y
+ sky130_fd_sc_hd__a2111oi_1
XANTENNA_75 _3526_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6552__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7587_ _7587_/CLK _7587_/D _6873_/A VGND VGND VPWR VPWR _7587_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_86 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4799_ _5107_/C _4807_/B _4799_/C VGND VGND VPWR VPWR _4800_/B sky130_fd_sc_hd__and3_1
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3905__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6538_ _7330_/Q _4105_/B _6561_/A2 _6420_/B _7306_/Q VGND VGND VPWR VPWR _6538_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6469_ _7367_/Q _6459_/B _6769_/A3 _6468_/X _7407_/Q VGND VGND VPWR VPWR _6469_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput171 _4175_/X VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_121_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput182 _3429_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 _3419_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6419__A _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2940 _7063_/Q VGND VGND VPWR VPWR hold2940/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2951 hold2951/A VGND VGND VPWR VPWR _4530_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2962 hold2962/A VGND VGND VPWR VPWR _4367_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_153_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2973 hold2973/A VGND VGND VPWR VPWR hold2973/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2984 _7519_/Q VGND VGND VPWR VPWR hold2984/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2995 _6999_/Q VGND VGND VPWR VPWR _4320_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3841__A1 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3841__B2 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3497__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5594__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6791__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5346__A1 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6543__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5932__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__C1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4609__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4085__A1 _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5840_ _5840_/A0 _5876_/A1 _5847_/S VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _5771_/A0 _5969_/A1 _5775_/S VGND VGND VPWR VPWR _5771_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7510_ _7525_/CLK hold98/X fanout745/X VGND VGND VPWR VPWR _7510_/Q sky130_fd_sc_hd__dfrtp_4
X_4722_ _5399_/A _5399_/B VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__6129__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7441_ _7561_/CLK _7441_/D fanout741/X VGND VGND VPWR VPWR _7441_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6534__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4653_ _4644_/Y _4646_/Y _4833_/A VGND VGND VPWR VPWR _5248_/A sky130_fd_sc_hd__o21a_4
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__buf_2
X_3604_ _7429_/Q hold32/A _5965_/B _3562_/X _7301_/Q VGND VGND VPWR VPWR _3604_/X
+ sky130_fd_sc_hd__a32o_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
X_7372_ _7421_/CLK _7372_/D fanout715/X VGND VGND VPWR VPWR _7372_/Q sky130_fd_sc_hd__dfrtp_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR _3859_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4584_ _4675_/A _4675_/B _4643_/C _4823_/D VGND VGND VPWR VPWR _4593_/A sky130_fd_sc_hd__nand4_4
Xhold802 hold802/A VGND VGND VPWR VPWR _7284_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR _4134_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap521 _4721_/Y VGND VGND VPWR VPWR _4807_/B sky130_fd_sc_hd__clkbuf_4
Xhold813 hold813/A VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_4
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_2
Xhold824 hold824/A VGND VGND VPWR VPWR _7373_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6323_ _7133_/Q _6091_/X _6082_/C _6322_/X VGND VGND VPWR VPWR _6323_/X sky130_fd_sc_hd__a31o_1
Xhold835 hold835/A VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3535_ _5938_/A _5938_/C _4509_/C VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__and3_4
Xhold846 hold846/A VGND VGND VPWR VPWR _7119_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold857 hold857/A VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold868 hold868/A VGND VGND VPWR VPWR _7057_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold879 hold879/A VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6254_ _7405_/Q _6091_/X _6119_/D _7469_/Q _6087_/X VGND VGND VPWR VPWR _6254_/X
+ sky130_fd_sc_hd__a32o_1
X_3466_ hold340/X _4025_/A _4181_/S VGND VGND VPWR VPWR _3466_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__6301__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2203 _4351_/X VGND VGND VPWR VPWR hold544/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5205_ wire375/X _5059_/A _5061_/B _4969_/Y VGND VGND VPWR VPWR _5205_/X sky130_fd_sc_hd__a31o_1
Xhold2214 _5676_/X VGND VGND VPWR VPWR hold560/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6185_ _7458_/Q _6075_/A _6079_/X _6094_/X _7506_/Q VGND VGND VPWR VPWR _6185_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2225 hold635/X VGND VGND VPWR VPWR _5689_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2236 _5720_/X VGND VGND VPWR VPWR hold672/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1502 _7468_/Q VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2247 _5761_/X VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5136_ _4687_/Y _5135_/Y _5134_/X VGND VGND VPWR VPWR _5139_/B sky130_fd_sc_hd__o21ba_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2258 hold587/X VGND VGND VPWR VPWR _5628_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1513 hold177/X VGND VGND VPWR VPWR _7545_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2269 hold641/X VGND VGND VPWR VPWR _5960_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1524 _7564_/Q VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1535 hold200/X VGND VGND VPWR VPWR _5962_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_123_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1546 hold228/X VGND VGND VPWR VPWR _5944_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1557 _7669_/A VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5067_ _5091_/C _5260_/C _5067_/C VGND VGND VPWR VPWR _5067_/X sky130_fd_sc_hd__and3_1
Xhold1568 _5976_/A0 VGND VGND VPWR VPWR _5985_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1579 hold222/X VGND VGND VPWR VPWR _5908_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5273__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4018_ hold44/A _6905_/Q _6904_/Q _4025_/B _3451_/Y VGND VGND VPWR VPWR _4018_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_84_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3823__A1 _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3598__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3823__B2 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6405__C _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6368__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5969_ _5969_/A0 _5969_/A1 _5973_/S VGND VGND VPWR VPWR _5969_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7639_ _7641_/CLK _7639_/D fanout751/X VGND VGND VPWR VPWR _7639_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6525__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6421__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input165_A wb_sel_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4854__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input26_A mask_rev_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2770 hold953/X VGND VGND VPWR VPWR _4374_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2781 _7150_/Q VGND VGND VPWR VPWR hold971/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2792 hold785/X VGND VGND VPWR VPWR _4205_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3814__B2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4116__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7180__RESET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3593__A3 _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3674__C _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold109 hold109/A VGND VGND VPWR VPWR _7286_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6531__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_max_cap430_A _5012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_50_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5255__B1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6941_ _7330_/CLK _6941_/D fanout711/X VGND VGND VPWR VPWR _6941_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2597_A _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5270__A3 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6872_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6872_/X sky130_fd_sc_hd__and2_1
XFILLER_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5823_ _5823_/A0 _5994_/A1 hold33/X VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5558__A1 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6755__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5558__B2 _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5837__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5754_ _5754_/A0 _5952_/A1 _5757_/S VGND VGND VPWR VPWR _5754_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3865__B _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4705_ _4825_/A _5115_/A _5089_/B VGND VGND VPWR VPWR _4705_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__6507__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5685_ _5685_/A0 _5955_/A1 _5685_/S VGND VGND VPWR VPWR _5685_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2931_A _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7424_ _7472_/CLK _7424_/D fanout719/X VGND VGND VPWR VPWR _7424_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_190_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4636_ _4814_/C _5494_/B2 _4772_/A VGND VGND VPWR VPWR _4636_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_190_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold610 hold610/A VGND VGND VPWR VPWR _7563_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5730__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold621 hold621/A VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7355_ _7563_/CLK _7355_/D fanout739/X VGND VGND VPWR VPWR _7355_/Q sky130_fd_sc_hd__dfrtp_4
X_4567_ _4909_/D _4772_/B VGND VGND VPWR VPWR _4667_/A sky130_fd_sc_hd__nand2_8
Xhold632 _5739_/X VGND VGND VPWR VPWR _7350_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6306_ _6009_/B _7609_/Q _6304_/X _6305_/X VGND VGND VPWR VPWR _6306_/X sky130_fd_sc_hd__a22o_1
Xhold654 hold654/A VGND VGND VPWR VPWR _7213_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold665 hold665/A VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3518_ hold47/A _5938_/A _4455_/A VGND VGND VPWR VPWR _5758_/A sky130_fd_sc_hd__and3_4
X_7286_ _7309_/CLK _7286_/D fanout710/X VGND VGND VPWR VPWR _7286_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold676 hold676/A VGND VGND VPWR VPWR _7386_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4498_ _5912_/A1 _4498_/A1 _4502_/S VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__mux2_1
Xhold687 hold687/A VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6286__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold698 hold698/A VGND VGND VPWR VPWR _7005_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6237_ _6649_/S _6237_/A2 _6573_/S _6236_/X VGND VGND VPWR VPWR _6237_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout582_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2000 _5743_/X VGND VGND VPWR VPWR hold418/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3449_ _3449_/A0 hold122/X _4181_/S VGND VGND VPWR VPWR _3449_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4297__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2011 hold455/X VGND VGND VPWR VPWR _5788_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2022 hold419/X VGND VGND VPWR VPWR _5977_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2033 hold497/X VGND VGND VPWR VPWR _5697_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2044 hold330/X VGND VGND VPWR VPWR _5826_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6168_ _6036_/Y _7281_/Q _6167_/X _6157_/Y _6067_/A VGND VGND VPWR VPWR _6168_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _5750_/X VGND VGND VPWR VPWR _7359_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2055 hold479/X VGND VGND VPWR VPWR _4499_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1321 hold3180/X VGND VGND VPWR VPWR hold3181/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2066 _5778_/X VGND VGND VPWR VPWR hold502/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2077 hold517/X VGND VGND VPWR VPWR _5877_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1332 hold3161/X VGND VGND VPWR VPWR _7167_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1343 hold3205/X VGND VGND VPWR VPWR hold3206/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5119_ _5059_/B _5115_/X _5118_/X _5117_/Y VGND VGND VPWR VPWR _5119_/X sky130_fd_sc_hd__a211o_1
Xhold2088 hold22/X VGND VGND VPWR VPWR _5856_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1354 _4296_/B VGND VGND VPWR VPWR hold2981/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6099_ _6332_/B _6081_/C _6112_/B _6099_/D VGND VGND VPWR VPWR _6099_/X sky130_fd_sc_hd__and4bb_4
Xhold2099 _7438_/Q VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6589__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1365 _4288_/A1 VGND VGND VPWR VPWR hold2975/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1376 _6781_/B VGND VGND VPWR VPWR hold3064/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1387 hold2149/X VGND VGND VPWR VPWR hold2150/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1398 hold1422/X VGND VGND VPWR VPWR hold1423/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_41_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6746__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5747__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6210__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4221__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3494__C _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6277__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3290 _6284_/X VGND VGND VPWR VPWR _7609_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5788__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3669__C _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4460__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6737__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6201__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3566__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5960__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5470_ _4605_/Y _5563_/A1 _4971_/X _5265_/A _5469_/Y VGND VGND VPWR VPWR _5564_/B
+ sky130_fd_sc_hd__o311a_2
X_4421_ _4421_/A0 _4420_/X _4423_/S VGND VGND VPWR VPWR _4421_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3723__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7140_ _7185_/CLK _7140_/D fanout737/X VGND VGND VPWR VPWR _7140_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4352_ _4352_/A _4352_/B _4533_/B VGND VGND VPWR VPWR _4357_/S sky130_fd_sc_hd__and3_2
Xfanout408 hold124/X VGND VGND VPWR VPWR _3598_/B sky130_fd_sc_hd__buf_4
XANTENNA__6268__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7071_ _7075_/CLK _7071_/D _6861_/X VGND VGND VPWR VPWR _7071_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_98_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4283_ _4289_/S _4283_/B VGND VGND VPWR VPWR _4283_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4279__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6022_ _7588_/Q _7589_/Q VGND VGND VPWR VPWR _6022_/X sky130_fd_sc_hd__and2b_2
XFILLER_113_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3487__C1 _3479_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6924_ _7264_/CLK _6924_/D fanout688/X VGND VGND VPWR VPWR _6924_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6440__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4451__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6855_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5806_ _5806_/A0 _5950_/A1 _5811_/S VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__mux2_1
X_6786_ _6792_/S _6786_/B VGND VGND VPWR VPWR _6786_/Y sky130_fd_sc_hd__nand2_1
X_3998_ _4058_/B _7073_/Q VGND VGND VPWR VPWR _3998_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5951__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5737_ _5737_/A0 _5953_/A1 _5739_/S VGND VGND VPWR VPWR _5737_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3962__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5668_ _5668_/A _5947_/C VGND VGND VPWR VPWR _5676_/S sky130_fd_sc_hd__nand2_8
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4203__C _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7407_ _7497_/CLK _7407_/D fanout707/X VGND VGND VPWR VPWR _7407_/Q sky130_fd_sc_hd__dfstp_2
X_4619_ _4570_/Y _4608_/Y _4618_/Y VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5703__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5599_ _5599_/A0 _5815_/A1 _5602_/S VGND VGND VPWR VPWR _5599_/X sky130_fd_sc_hd__mux2_1
Xhold440 _5972_/X VGND VGND VPWR VPWR _7557_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7338_ _7576_/CLK hold14/X fanout717/X VGND VGND VPWR VPWR _7338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold451 hold451/A VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold462 hold462/A VGND VGND VPWR VPWR _7123_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold473 hold473/A VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold484 hold484/A VGND VGND VPWR VPWR _7083_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6259__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold495 hold495/A VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7269_ _7522_/CLK _7269_/D fanout744/X VGND VGND VPWR VPWR _7269_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6427__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1140 hold3121/X VGND VGND VPWR VPWR _7197_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 hold1151/A VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XTAP_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1162 hold3023/X VGND VGND VPWR VPWR hold1162/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1173 hold2884/X VGND VGND VPWR VPWR hold2885/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input128_A wb_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1184 hold1184/A VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1195 hold3156/X VGND VGND VPWR VPWR hold3157/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1981_A _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5234__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6719__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__B2 _7315_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input93_A trap VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3953__B1 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5170__A2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3720__A3 _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6670__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6903__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4970_ _5248_/A _5248_/B _4970_/C VGND VGND VPWR VPWR _5052_/A sky130_fd_sc_hd__and3_1
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3921_ _3897_/X _3904_/X _3921_/C _3921_/D VGND VGND VPWR VPWR _3922_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__3787__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6640_ _7446_/Q _6574_/B _6574_/C _6434_/X _7470_/Q VGND VGND VPWR VPWR _6640_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6186__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3852_ input37/X _4231_/S _4467_/A _7129_/Q _3851_/X VGND VGND VPWR VPWR _3852_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__6186__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6571_ _7283_/Q _6431_/Y _6623_/B1 VGND VGND VPWR VPWR _6571_/X sky130_fd_sc_hd__o21a_1
X_3783_ _6914_/Q _5619_/A _5947_/A _3617_/X _7232_/Q VGND VGND VPWR VPWR _3792_/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_164_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3944__B1 _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5522_ _4668_/C _4827_/X _5107_/X _5110_/X VGND VGND VPWR VPWR _5559_/C sky130_fd_sc_hd__a211o_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6489__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5453_ _5453_/A _5453_/B _5453_/C VGND VGND VPWR VPWR _5453_/X sky130_fd_sc_hd__and3_1
XFILLER_173_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3862__C _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4404_ _4404_/A0 _5647_/A0 _4405_/S VGND VGND VPWR VPWR _4404_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_42_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7579_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_126_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5384_ _5384_/A _5384_/B _5384_/C VGND VGND VPWR VPWR _5390_/A sky130_fd_sc_hd__and3_1
XANTENNA__5161__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7123_ _7186_/CLK _7123_/D fanout725/X VGND VGND VPWR VPWR _7123_/Q sky130_fd_sc_hd__dfrtp_4
X_4335_ _4335_/A0 _5894_/A0 _4339_/S VGND VGND VPWR VPWR _4335_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5850__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7212_/CLK _7054_/D fanout721/X VGND VGND VPWR VPWR _7054_/Q sky130_fd_sc_hd__dfrtp_4
X_4266_ _4266_/A0 _5582_/A0 _4270_/S VGND VGND VPWR VPWR _4266_/X sky130_fd_sc_hd__mux2_1
X_6005_ _7584_/Q _6006_/A VGND VGND VPWR VPWR _6005_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_57_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7334_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6661__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4197_ _4197_/A0 _7642_/Q _4429_/B VGND VGND VPWR VPWR _4197_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout545_A _4447_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _7075_/CLK _6907_/D _6857_/X VGND VGND VPWR VPWR _6907_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3778__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6838_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6838_/X sky130_fd_sc_hd__and2_1
XANTENNA__6177__A1 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6177__B2 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6413__C _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6716__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6769_ _7040_/Q _6459_/B _6769_/A3 _6421_/X _7010_/Q VGND VGND VPWR VPWR _6769_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3935__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5137__C1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5688__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3950__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5152__A2 _4758_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold270 hold270/A VGND VGND VPWR VPWR _7290_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5045__B _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold281 hold281/A VGND VGND VPWR VPWR _7170_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5760__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout750 input75/X VGND VGND VPWR VPWR fanout750/X sky130_fd_sc_hd__buf_12
Xfanout761 input126/X VGND VGND VPWR VPWR _4831_/C sky130_fd_sc_hd__buf_8
Xfanout772 _5004_/A1 VGND VGND VPWR VPWR _4825_/A sky130_fd_sc_hd__buf_8
XANTENNA__6652__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_804 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5860__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4663__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5061__A _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6168__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6707__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output297_A _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5935__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3926__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5391__A2 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4778__C _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4140__A _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6340__B2 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4120_ _6882_/Q _4058_/A _4123_/B _4120_/B1 VGND VGND VPWR VPWR _4120_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1909 _7251_/Q VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6643__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4051_ _3998_/Y _4062_/A _4120_/B1 _4051_/B1 VGND VGND VPWR VPWR _6896_/D sky130_fd_sc_hd__a31o_1
XANTENNA__6067__A _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__C1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5851__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4406__A1 _5650_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4953_ _4954_/A _5248_/A _4954_/C VGND VGND VPWR VPWR _4953_/X sky130_fd_sc_hd__and3_4
XANTENNA_clkbuf_3_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3904_ _7062_/Q _4394_/A _3899_/X _3901_/X _3903_/X VGND VGND VPWR VPWR _3904_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_178_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7672_ _7672_/A VGND VGND VPWR VPWR _7672_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4315__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4884_ _5065_/A _4884_/B _4907_/B _4970_/C VGND VGND VPWR VPWR _5448_/D sky130_fd_sc_hd__nand4_2
X_6623_ _7285_/Q _6431_/Y _6623_/B1 VGND VGND VPWR VPWR _6623_/X sky130_fd_sc_hd__o21a_1
X_3835_ _7058_/Q _4539_/C _5623_/B _3834_/X VGND VGND VPWR VPWR _3835_/X sky130_fd_sc_hd__a31o_1
XFILLER_193_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3917__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6554_ _7403_/Q _6409_/X _6549_/X _6553_/X _6430_/X VGND VGND VPWR VPWR _6554_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3766_ _7458_/Q _4431_/A _5866_/B _3537_/X _7426_/Q VGND VGND VPWR VPWR _3766_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5505_ _5203_/A _5089_/D _5549_/A3 _5504_/Y VGND VGND VPWR VPWR _5505_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4135__A_N _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3932__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6485_ _7480_/Q _6451_/X _6480_/X _6482_/X _6484_/X VGND VGND VPWR VPWR _6485_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3697_ _7136_/Q _4473_/A _5619_/B _3661_/X _7035_/Q VGND VGND VPWR VPWR _3697_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5436_ _5339_/D _5339_/C _5425_/X _5170_/X VGND VGND VPWR VPWR _5436_/X sky130_fd_sc_hd__a31o_1
Xoutput320 hold1086/X VGND VGND VPWR VPWR hold1087/A sky130_fd_sc_hd__buf_6
XFILLER_145_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput331 hold1162/X VGND VGND VPWR VPWR hold1163/A sky130_fd_sc_hd__buf_6
Xoutput342 hold2973/X VGND VGND VPWR VPWR hold1085/A sky130_fd_sc_hd__buf_6
XANTENNA__4342__A0 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6676__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5367_ _5545_/B _5367_/B _5367_/C _5367_/D VGND VGND VPWR VPWR _5367_/Y sky130_fd_sc_hd__nor4_2
XFILLER_113_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7106_ _7111_/CLK _7106_/D fanout751/X VGND VGND VPWR VPWR _7106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4318_ _4321_/S _3734_/B _4317_/Y VGND VGND VPWR VPWR _6997_/D sky130_fd_sc_hd__o21ai_2
XFILLER_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5298_ _4583_/B _4821_/Y _4735_/Y _4687_/Y VGND VGND VPWR VPWR _5298_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6095__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7037_ _7164_/CLK _7037_/D fanout698/X VGND VGND VPWR VPWR _7037_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6634__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4249_ _4249_/A0 _4248_/X _4249_/S VGND VGND VPWR VPWR _4249_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6408__C _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4660__A4 _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__B2 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3620__A2 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5373__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire469 _4632_/Y VGND VGND VPWR VPWR _4753_/C sky130_fd_sc_hd__buf_2
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3060_A _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6322__A1 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A mgmt_gpio_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3687__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout580 hold1567/X VGND VGND VPWR VPWR _4553_/A0 sky130_fd_sc_hd__buf_6
XANTENNA__4636__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout591 hold2518/X VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__buf_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6389__A1 _7030_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3611__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3620_ _5659_/B _5623_/B _3619_/X _3558_/X _7284_/Q VGND VGND VPWR VPWR _3620_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4789__B _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3551_ input51/X _3637_/C _3738_/B _5920_/A hold52/A VGND VGND VPWR VPWR _3551_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3914__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6270_ _7414_/Q _6144_/C _6089_/C _6270_/C1 VGND VGND VPWR VPWR _6270_/X sky130_fd_sc_hd__o211a_1
X_3482_ _5803_/A _5640_/A _5722_/B VGND VGND VPWR VPWR _5794_/A sky130_fd_sc_hd__and3_4
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4324__A0 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5221_ _5065_/A _5220_/X _5219_/Y VGND VGND VPWR VPWR _5223_/B sky130_fd_sc_hd__a21oi_1
Xhold3108 _7112_/Q VGND VGND VPWR VPWR hold3108/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3119 _7197_/Q VGND VGND VPWR VPWR hold3119/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3678__A2 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2407 _5816_/X VGND VGND VPWR VPWR hold682/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2418 hold655/X VGND VGND VPWR VPWR _5916_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5152_ _4794_/A _4758_/X _5410_/B _5096_/A _5152_/B2 VGND VGND VPWR VPWR _5153_/C
+ sky130_fd_sc_hd__a32oi_4
Xhold2429 _7365_/Q VGND VGND VPWR VPWR hold799/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6077__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1706 hold271/X VGND VGND VPWR VPWR _5904_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4103_ _6441_/D _6433_/D VGND VGND VPWR VPWR _6455_/B sky130_fd_sc_hd__and2b_4
XANTENNA__6616__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1717 hold335/X VGND VGND VPWR VPWR _7544_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5083_ _5563_/A1 _4720_/Y _5516_/A3 _4748_/Y _4717_/Y VGND VGND VPWR VPWR _5083_/X
+ sky130_fd_sc_hd__o32a_1
Xhold1728 _5661_/X VGND VGND VPWR VPWR hold388/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1739 hold232/X VGND VGND VPWR VPWR _4332_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4627__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4034_ _6902_/Q _6901_/Q _6900_/Q _6903_/Q VGND VGND VPWR VPWR _4034_/X sky130_fd_sc_hd__a31o_1
XFILLER_65_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3850__A2 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5985_ _5985_/A0 _5985_/A1 _5991_/S VGND VGND VPWR VPWR _5985_/X sky130_fd_sc_hd__mux2_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4936_ _4954_/A _4940_/D VGND VGND VPWR VPWR _4936_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3602__A2 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_10 _3902_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7655_ _7655_/A VGND VGND VPWR VPWR _7655_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_21 _6585_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4947_/C _4942_/A _4948_/C VGND VGND VPWR VPWR _4933_/B sky130_fd_sc_hd__and3_4
XANTENNA_32 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_54 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ _7309_/Q _6420_/B _6425_/X _7341_/Q _6605_/X VGND VGND VPWR VPWR _6606_/X
+ sky130_fd_sc_hd__a221o_1
X_3818_ _7003_/Q _4322_/A _3799_/X _3815_/X _3817_/X VGND VGND VPWR VPWR _3818_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout410_A _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4158__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7586_ _7601_/CLK _7586_/D _6873_/A VGND VGND VPWR VPWR _7586_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_65 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _3583_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4699__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ _5107_/C _4799_/C VGND VGND VPWR VPWR _4798_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_fanout508_A _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _7002_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6537_ _7362_/Q _6462_/X _6468_/X _7410_/Q _6536_/X VGND VGND VPWR VPWR _6544_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3905__A3 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3749_ _7115_/Q _3658_/X _3661_/X _7034_/Q _3748_/X VGND VGND VPWR VPWR _3749_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6468_ _6574_/B _6600_/B _6468_/C VGND VGND VPWR VPWR _6468_/X sky130_fd_sc_hd__and3_4
X_5419_ _5419_/A _5419_/B _5491_/A VGND VGND VPWR VPWR _5419_/X sky130_fd_sc_hd__and3_1
X_6399_ _6961_/Q _6036_/Y _6067_/A VGND VGND VPWR VPWR _6399_/X sky130_fd_sc_hd__o21a_1
Xoutput172 _7648_/X VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
Xoutput183 _3428_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
XFILLER_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput194 _3418_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_102_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold288_A _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2930 hold2930/A VGND VGND VPWR VPWR _4506_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2941 hold2941/A VGND VGND VPWR VPWR _4397_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6607__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2952 _4530_/X VGND VGND VPWR VPWR hold2952/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4618__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2963 _6979_/Q VGND VGND VPWR VPWR _4289_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2974 _6978_/Q VGND VGND VPWR VPWR _4288_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2985 hold2985/A VGND VGND VPWR VPWR _5930_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2996 hold2996/A VGND VGND VPWR VPWR hold2996/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6083__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5291__A1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input110_A wb_adr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3497__C _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6543__A1 _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6543__B2 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4554__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__B1 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4609__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4085__A2 _4085_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5019__D1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3832__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ hold214/X _5986_/A1 _5775_/S VGND VGND VPWR VPWR _5770_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6782__A1 _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _5058_/D _4856_/A _5073_/A VGND VGND VPWR VPWR _4721_/Y sky130_fd_sc_hd__nor3_2
XFILLER_159_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7440_ _7522_/CLK _7440_/D fanout743/X VGND VGND VPWR VPWR _7440_/Q sky130_fd_sc_hd__dfstp_4
X_4652_ _4648_/A _4591_/Y _5005_/A _4726_/B VGND VGND VPWR VPWR _5222_/C sky130_fd_sc_hd__o211a_4
XANTENNA__6534__A1 _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3603_ _7445_/Q _3520_/X _5920_/A _7517_/Q _3602_/X VGND VGND VPWR VPWR _3606_/C
+ sky130_fd_sc_hd__a221o_1
X_7371_ _7574_/CLK _7371_/D fanout729/X VGND VGND VPWR VPWR _7371_/Q sky130_fd_sc_hd__dfrtp_4
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4583_ _4646_/A _4583_/B VGND VGND VPWR VPWR _4586_/C sky130_fd_sc_hd__nor2_2
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR _4174_/A sky130_fd_sc_hd__buf_8
Xhold803 hold803/A VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR _4135_/B sky130_fd_sc_hd__buf_4
X_6322_ _7143_/Q _6082_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6322_/X sky130_fd_sc_hd__o211a_1
Xhold814 _5772_/X VGND VGND VPWR VPWR _7379_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_4
Xhold825 hold825/A VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3534_ _7534_/Q _3529_/X _5857_/A _7462_/Q _3533_/X VGND VGND VPWR VPWR _3534_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__buf_4
XFILLER_115_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold836 _5882_/X VGND VGND VPWR VPWR _7477_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6298__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold858 hold858/A VGND VGND VPWR VPWR _7125_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6253_ _7461_/Q _6112_/C _6079_/X _6094_/X _7509_/Q VGND VGND VPWR VPWR _6253_/X
+ sky130_fd_sc_hd__a32o_1
Xhold869 hold869/A VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3465_ _4076_/B _4025_/A VGND VGND VPWR VPWR _3465_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_88_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4966__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5204_ _5495_/C1 _4679_/Y _4880_/Y _5203_/Y VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__o31a_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2204 _6926_/Q VGND VGND VPWR VPWR hold523/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6184_ _7418_/Q _6072_/X _6144_/X _7290_/Q _6183_/X VGND VGND VPWR VPWR _6184_/X
+ sky130_fd_sc_hd__a221o_1
Xhold2215 _7334_/Q VGND VGND VPWR VPWR hold563/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2226 _5689_/X VGND VGND VPWR VPWR hold636/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2237 _7281_/Q VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5135_ _4807_/B _5077_/B _5297_/B _5029_/A VGND VGND VPWR VPWR _5135_/Y sky130_fd_sc_hd__a22oi_2
Xhold1503 hold259/X VGND VGND VPWR VPWR _5872_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2248 _7378_/Q VGND VGND VPWR VPWR hold619/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2259 _7354_/Q VGND VGND VPWR VPWR hold613/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1514 _7572_/Q VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1525 hold255/X VGND VGND VPWR VPWR _5980_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1536 _5962_/X VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1547 _5944_/X VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1558 hold316/X VGND VGND VPWR VPWR _4437_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5066_ _5096_/A _5453_/C VGND VGND VPWR VPWR _5444_/B sky130_fd_sc_hd__nand2_2
Xhold1569 _4252_/X VGND VGND VPWR VPWR hold262/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6470__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4017_ hold44/A _4017_/B VGND VGND VPWR VPWR _4017_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout360_A _3549_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout458_A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3598__B _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6758__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6222__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5968_ _5968_/A0 _5968_/A1 _5973_/S VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _4919_/A _5573_/C _4919_/C VGND VGND VPWR VPWR _4922_/C sky130_fd_sc_hd__nand3_1
X_5899_ _5998_/A1 _5899_/A1 _5901_/S VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6702__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4503__A _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7638_ _7641_/CLK _7638_/D fanout751/X VGND VGND VPWR VPWR _7638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6525__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__B2 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4536__A0 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_806 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7569_ _7573_/CLK _7569_/D fanout733/X VGND VGND VPWR VPWR _7569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6828__A2 _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input158_A wb_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2760 _5696_/X VGND VGND VPWR VPWR hold542/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2771 _4374_/X VGND VGND VPWR VPWR hold954/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2782 hold971/X VGND VGND VPWR VPWR _4495_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2793 _7049_/Q VGND VGND VPWR VPWR hold889/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4384__S _4387_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input19_A mask_rev_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3814__A2 _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5016__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6764__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3750__A1 _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3463__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4786__C _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5255__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ _7578_/CLK _6940_/D fanout747/X VGND VGND VPWR VPWR _6940_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3805__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6871_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6871_/X sky130_fd_sc_hd__and2_1
XANTENNA__6204__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5822_ _5822_/A0 _5876_/A1 hold33/X VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5753_ _5753_/A0 _5951_/A1 _5757_/S VGND VGND VPWR VPWR _5753_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4704_ _4825_/A _5071_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4704_/Y sky130_fd_sc_hd__nor4_2
XANTENNA__3865__C _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5684_ _5684_/A0 _5972_/A1 _5685_/S VGND VGND VPWR VPWR _5684_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7423_ _7475_/CLK _7423_/D fanout730/X VGND VGND VPWR VPWR _7423_/Q sky130_fd_sc_hd__dfstp_1
X_4635_ _4747_/B _4574_/X _4733_/B VGND VGND VPWR VPWR _4730_/C sky130_fd_sc_hd__a21boi_4
XANTENNA__5853__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold600 hold600/A VGND VGND VPWR VPWR _6942_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7354_ _7575_/CLK _7354_/D fanout735/X VGND VGND VPWR VPWR _7354_/Q sky130_fd_sc_hd__dfrtp_4
X_4566_ _4909_/D _4772_/B VGND VGND VPWR VPWR _5100_/A sky130_fd_sc_hd__and2_4
Xhold611 hold611/A VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold622 hold622/A VGND VGND VPWR VPWR _7355_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6305_ _6957_/Q _6036_/Y _6067_/A VGND VGND VPWR VPWR _6305_/X sky130_fd_sc_hd__o21a_1
Xhold644 hold644/A VGND VGND VPWR VPWR _7281_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3741__A1 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3517_ _7242_/Q _3515_/X _5974_/A _7566_/Q _3513_/X VGND VGND VPWR VPWR _3524_/C
+ sky130_fd_sc_hd__a221o_1
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7285_ _7309_/CLK _7285_/D fanout710/X VGND VGND VPWR VPWR _7285_/Q sky130_fd_sc_hd__dfrtp_4
Xhold666 _5825_/X VGND VGND VPWR VPWR _7426_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4497_ _4497_/A _4551_/D VGND VGND VPWR VPWR _4502_/S sky130_fd_sc_hd__nand2_4
Xhold677 hold677/A VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold688 hold688/A VGND VGND VPWR VPWR _7020_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6236_ _6224_/X _6234_/X _6235_/X VGND VGND VPWR VPWR _6236_/X sky130_fd_sc_hd__o21a_1
Xhold699 hold699/A VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3448_ _4028_/A0 _6904_/Q _4025_/A VGND VGND VPWR VPWR _3448_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6286__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2001 _7385_/Q VGND VGND VPWR VPWR hold411/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2012 _7325_/Q VGND VGND VPWR VPWR hold409/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4297__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6691__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__B2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2023 _5977_/X VGND VGND VPWR VPWR hold420/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6161_/X _6163_/X _6164_/X _6166_/X VGND VGND VPWR VPWR _6167_/X sky130_fd_sc_hd__a211o_1
Xhold2034 _5697_/X VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2045 _7042_/Q VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout575_A hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 hold3263/X VGND VGND VPWR VPWR _7535_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1311 hold3185/X VGND VGND VPWR VPWR hold3186/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2056 _7557_/Q VGND VGND VPWR VPWR hold439/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1322 hold3182/X VGND VGND VPWR VPWR _7192_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2067 _7425_/Q VGND VGND VPWR VPWR hold473/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5118_ _5118_/A _5282_/C _5282_/D VGND VGND VPWR VPWR _5118_/X sky130_fd_sc_hd__and3_1
Xhold2078 _7411_/Q VGND VGND VPWR VPWR hold469/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1333 hold3213/X VGND VGND VPWR VPWR hold3214/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1344 hold3207/X VGND VGND VPWR VPWR _7006_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6098_ _7407_/Q _6097_/B _6144_/B _6097_/X _7439_/Q VGND VGND VPWR VPWR _6098_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2089 _5856_/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1355 _4302_/A1 VGND VGND VPWR VPWR hold2977/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1366 _4300_/A1 VGND VGND VPWR VPWR hold2983/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1377 _4298_/B VGND VGND VPWR VPWR hold3091/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout742_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5049_ _5339_/D _5203_/A _5049_/C _5339_/C VGND VGND VPWR VPWR _5051_/C sky130_fd_sc_hd__nand4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 hold2128/X VGND VGND VPWR VPWR hold2129/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1399 hold1473/X VGND VGND VPWR VPWR hold1474/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1592_A _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5549__A2 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1857_A _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5763__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4887__B _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold3140_A _7137_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3280 _6785_/Y VGND VGND VPWR VPWR _7631_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3291 _7606_/Q VGND VGND VPWR VPWR _6237_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2590 _5818_/X VGND VGND VPWR VPWR hold980/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3799__A1 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6737__A1 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6201__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ _4447_/A0 _4447_/A1 _4422_/S VGND VGND VPWR VPWR _4420_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4797__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3723__A1 _6992_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4351_ _4351_/A0 _5736_/A1 _4351_/S VGND VGND VPWR VPWR _4351_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3723__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4289__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2240_A _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7070_ _7160_/CLK _7070_/D _6872_/A VGND VGND VPWR VPWR _7070_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout409 _3872_/A2 VGND VGND VPWR VPWR _5983_/A sky130_fd_sc_hd__buf_6
X_4282_ _4289_/S _3856_/B _4281_/Y VGND VGND VPWR VPWR _6974_/D sky130_fd_sc_hd__o21ai_1
XFILLER_152_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4279__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6021_ _7589_/Q _7588_/Q VGND VGND VPWR VPWR _6021_/X sky130_fd_sc_hd__and2b_1
XFILLER_86_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3487__B1 _3486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ _7255_/CLK _6923_/D fanout688/X VGND VGND VPWR VPWR _6923_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__7489__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2874_A _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6854_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6854_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5805_ _5805_/A0 hold198/X _5811_/S VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__mux2_1
X_6785_ _6789_/A1 _3856_/B _6784_/Y VGND VGND VPWR VPWR _6785_/Y sky130_fd_sc_hd__o21ai_1
X_3997_ _3997_/A1 _3996_/A _3996_/Y _3923_/S VGND VGND VPWR VPWR _7214_/D sky130_fd_sc_hd__a22o_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7216__CLK_N _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5736_ _5736_/A0 _5736_/A1 _5739_/S VGND VGND VPWR VPWR _5736_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5667_ _5667_/A0 _6000_/A1 _5667_/S VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3962__B2 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4203__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4618_ _4667_/A _4899_/A2 _4831_/A VGND VGND VPWR VPWR _4618_/Y sky130_fd_sc_hd__o21bai_4
X_7406_ _7541_/CLK _7406_/D fanout711/X VGND VGND VPWR VPWR _7406_/Q sky130_fd_sc_hd__dfrtp_4
X_5598_ _5598_/A0 _5645_/A0 _5602_/S VGND VGND VPWR VPWR _5598_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7337_ _7539_/CLK _7337_/D fanout708/X VGND VGND VPWR VPWR _7337_/Q sky130_fd_sc_hd__dfrtp_4
Xhold430 _5616_/X VGND VGND VPWR VPWR _7245_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold441 hold441/A VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4549_ _5647_/A0 _4549_/A1 _4550_/S VGND VGND VPWR VPWR _4549_/X sky130_fd_sc_hd__mux2_1
Xhold452 hold452/A VGND VGND VPWR VPWR _7042_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold463 hold463/A VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold474 _5824_/X VGND VGND VPWR VPWR _7425_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold485 hold485/A VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7268_ _7268_/CLK _7268_/D _6869_/A VGND VGND VPWR VPWR _7268_/Q sky130_fd_sc_hd__dfrtp_1
Xhold496 hold496/A VGND VGND VPWR VPWR _7456_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_145_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6219_ _7516_/Q _6112_/C _6274_/A3 _6072_/X _7420_/Q VGND VGND VPWR VPWR _6219_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7199_ _7201_/CLK _7199_/D fanout728/X VGND VGND VPWR VPWR _7199_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5612__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1130 hold1130/A VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XTAP_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1141 hold3125/X VGND VGND VPWR VPWR hold3126/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1152 hold3150/X VGND VGND VPWR VPWR hold3151/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1163 hold1163/A VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
Xhold1174 _5599_/X VGND VGND VPWR VPWR _7231_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1185 hold3154/X VGND VGND VPWR VPWR hold3155/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1196 hold3158/X VGND VGND VPWR VPWR _7046_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6719__A1 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input86_A spimemio_flash_io0_oeb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3953__A1 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold3355_A _7628_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3705__A1 _7045_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__A1 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4969__B1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5630__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3920_ _7520_/Q hold77/A _5634_/A _7260_/Q _3919_/X VGND VGND VPWR VPWR _3921_/D
+ sky130_fd_sc_hd__a221oi_4
XFILLER_189_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3851_ _7545_/Q _4479_/A _5956_/B _5643_/A _4174_/A VGND VGND VPWR VPWR _3851_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6186__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6072__B _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6570_ _6554_/X _6570_/B _6570_/C VGND VGND VPWR VPWR _6570_/Y sky130_fd_sc_hd__nand3b_4
X_3782_ _3782_/A _3782_/B _3782_/C _3782_/D VGND VGND VPWR VPWR _3793_/C sky130_fd_sc_hd__nor4_1
XANTENNA__3944__A1 _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5521_ _5521_/A _5521_/B _5562_/C _5521_/D VGND VGND VPWR VPWR _5521_/Y sky130_fd_sc_hd__nand4_2
XFILLER_117_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5452_ _5510_/B _5452_/B _5574_/A VGND VGND VPWR VPWR _5456_/C sky130_fd_sc_hd__and3_1
XFILLER_173_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5697__A1 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4403_ _4403_/A0 _4548_/A0 _4405_/S VGND VGND VPWR VPWR _4403_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5383_ _5077_/Y _5255_/X _5378_/X _5380_/X _5382_/X VGND VGND VPWR VPWR _5384_/A
+ sky130_fd_sc_hd__o2111a_1
XFILLER_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7122_ _7186_/CLK _7122_/D fanout726/X VGND VGND VPWR VPWR _7122_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4334_ _4551_/A _4515_/B _4352_/A _4551_/D VGND VGND VPWR VPWR _4339_/S sky130_fd_sc_hd__and4_4
XFILLER_99_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5449__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7053_ _7164_/CLK _7053_/D fanout698/X VGND VGND VPWR VPWR _7053_/Q sky130_fd_sc_hd__dfstp_2
X_4265_ _4352_/B _4265_/B _4533_/B VGND VGND VPWR VPWR _4270_/S sky130_fd_sc_hd__and3_4
XFILLER_113_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6004_ _6009_/B _4107_/A _6932_/Q _6006_/A VGND VGND VPWR VPWR _6018_/A sky130_fd_sc_hd__a211o_1
XFILLER_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4196_ _4196_/A0 _5736_/A1 _4202_/S VGND VGND VPWR VPWR _4196_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5621__A1 _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ _7075_/CLK _6906_/D _6856_/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfrtp_2
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout538_A _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6837_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6837_/X sky130_fd_sc_hd__and2_1
XANTENNA__4188__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6768_ _7045_/Q _6408_/B _6425_/X _7020_/Q _6767_/X VGND VGND VPWR VPWR _6773_/B
+ sky130_fd_sc_hd__a221o_1
X_5719_ _5953_/A1 _5719_/A1 _5721_/S VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold116_A _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3935__B2 _7559_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6699_ _6958_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6699_/X sky130_fd_sc_hd__o21a_1
XFILLER_108_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5137__B1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6334__C1 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3699__B1 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 hold260/A VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4360__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold282 hold282/A VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6101__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout740 fanout749/X VGND VGND VPWR VPWR fanout740/X sky130_fd_sc_hd__buf_6
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5342__A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout751 fanout753/X VGND VGND VPWR VPWR fanout751/X sky130_fd_sc_hd__buf_8
XANTENNA_input140_A wb_dat_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout762 _4805_/B VGND VGND VPWR VPWR _4772_/B sky130_fd_sc_hd__buf_12
Xfanout773 _5071_/A VGND VGND VPWR VPWR _4674_/A sky130_fd_sc_hd__buf_12
XFILLER_19_816 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5061__B _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6168__A2 _7281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3926__A1 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_user_clock_A user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5679__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6340__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4351__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6628__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ _6897_/Q _3400_/A _4050_/S VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5300__B1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6067__B _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4406__A2 hold365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4952_ _5222_/A _4952_/B VGND VGND VPWR VPWR _4958_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3614__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3903_ _7448_/Q _5848_/A _3520_/X _7440_/Q _3902_/X VGND VGND VPWR VPWR _3903_/X
+ sky130_fd_sc_hd__a221o_1
X_7671_ _7671_/A VGND VGND VPWR VPWR _7671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4883_ _5180_/A _5216_/A _5342_/B VGND VGND VPWR VPWR _4904_/A sky130_fd_sc_hd__and3_2
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6622_ _7293_/Q _6422_/X _6604_/X _6615_/X _6621_/X VGND VGND VPWR VPWR _6622_/X
+ sky130_fd_sc_hd__a2111o_2
X_3834_ _7053_/Q _3931_/B _5619_/B _3544_/X _7417_/Q VGND VGND VPWR VPWR _3834_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6553_ _7531_/Q _6058_/X _6551_/X _6552_/X VGND VGND VPWR VPWR _6553_/X sky130_fd_sc_hd__a211o_1
X_3765_ _7160_/Q _4527_/A _4352_/B _4394_/A _7064_/Q VGND VGND VPWR VPWR _3765_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5382__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5504_ _5572_/A _5504_/B _5550_/A _5550_/B VGND VGND VPWR VPWR _5504_/Y sky130_fd_sc_hd__nand4_1
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6484_ _7304_/Q _6420_/B _6454_/X _7488_/Q _6483_/X VGND VGND VPWR VPWR _6484_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3696_ _7196_/Q _4545_/A _3690_/X _3691_/X _3695_/X VGND VGND VPWR VPWR _3733_/C
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_145_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xpad_flashh_clk_buff_inst _4127_/X VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_8
X_5435_ _5499_/A _5435_/B _5501_/A _5435_/D VGND VGND VPWR VPWR _5438_/A sky130_fd_sc_hd__nor4_1
XFILLER_161_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput310 _7673_/X VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 hold1090/X VGND VGND VPWR VPWR hold1091/A sky130_fd_sc_hd__buf_6
XANTENNA__5861__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput332 hold1208/X VGND VGND VPWR VPWR hold1209/A sky130_fd_sc_hd__buf_6
Xoutput343 hold1074/X VGND VGND VPWR VPWR hold1075/A sky130_fd_sc_hd__buf_6
X_5366_ _5248_/B _5453_/A _5243_/C _5367_/D VGND VGND VPWR VPWR _5366_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4985__B _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6619__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7105_ _7646_/CLK _7105_/D fanout751/X VGND VGND VPWR VPWR _7105_/Q sky130_fd_sc_hd__dfrtp_4
X_4317_ _4321_/S _4317_/B VGND VGND VPWR VPWR _4317_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout390_A _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5297_ _5297_/A _5297_/B VGND VGND VPWR VPWR _5297_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout488_A _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6095__A1 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7036_ _7164_/CLK _7036_/D fanout699/X VGND VGND VPWR VPWR _7036_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6095__B2 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4248_ hold607/X _6000_/A1 _4248_/S VGND VGND VPWR VPWR _4248_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5842__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6408__D _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7433__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4179_ _4179_/A0 hold24/X _4429_/B VGND VGND VPWR VPWR _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_41_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3605__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1672_A _7525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3620__A3 _3619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold1937_A _7422_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6322__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5771__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3687__A3 _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input49_A mgmt_gpio_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4387__S _4387_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_790 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5072__A _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout570 _5968_/A1 VGND VGND VPWR VPWR _5995_/A1 sky130_fd_sc_hd__buf_8
XANTENNA__5833__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4636__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout581 hold1567/X VGND VGND VPWR VPWR _5976_/A0 sky130_fd_sc_hd__buf_8
Xfanout592 hold26/X VGND VGND VPWR VPWR _5640_/D sky130_fd_sc_hd__buf_8
XFILLER_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6389__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_41_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7548_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4135__B _4135_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7330_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6561__A2 _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5364__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3550_ _5992_/A _5938_/A _4376_/B VGND VGND VPWR VPWR _5920_/A sky130_fd_sc_hd__and3_4
XFILLER_143_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6777__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3481_ _5938_/A _5938_/B VGND VGND VPWR VPWR _3481_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6313__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5220_ _5213_/A _5213_/C _4918_/D _5248_/C _5077_/B VGND VGND VPWR VPWR _5220_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3109 hold3109/A VGND VGND VPWR VPWR _4450_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3678__A3 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5151_ _5561_/A1 _4722_/Y _4787_/Y _4821_/Y _4783_/Y VGND VGND VPWR VPWR _5153_/B
+ sky130_fd_sc_hd__o32a_1
Xhold2408 _7005_/Q VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2419 _5916_/X VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6077__A1 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4102_ _7597_/Q _7598_/Q VGND VGND VPWR VPWR _6427_/A sky130_fd_sc_hd__and2b_4
XFILLER_111_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1707 _5904_/X VGND VGND VPWR VPWR _7496_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5082_ _4717_/Y _4748_/Y _5516_/A3 _4727_/Y _5081_/Y VGND VGND VPWR VPWR _5084_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6616__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1718 _7360_/Q VGND VGND VPWR VPWR hold332/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1729 _7665_/A VGND VGND VPWR VPWR hold421/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5824__A1 _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4627__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4033_ _4033_/A0 _4032_/X _4040_/A VGND VGND VPWR VPWR _6904_/D sky130_fd_sc_hd__mux2_1
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4872__A_N _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _5984_/A0 _5993_/A1 _5991_/S VGND VGND VPWR VPWR _5984_/X sky130_fd_sc_hd__mux2_1
X_4935_ _4954_/A _5453_/A _4940_/D VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__and3_1
Xclkbuf_3_7_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_7_0_csclk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5856__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3602__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_11 _3921_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7654_ _7654_/A VGND VGND VPWR VPWR _7654_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_22 _6647_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _5183_/C _4933_/A _5180_/A VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__and3_1
XFILLER_193_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ _7493_/Q _6463_/A _6441_/X _6409_/X _7405_/Q VGND VGND VPWR VPWR _6605_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_55 _7224_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ _7281_/Q _3558_/X _3659_/X _7008_/Q _3816_/X VGND VGND VPWR VPWR _3817_/X
+ sky130_fd_sc_hd__a221o_1
X_7585_ _7601_/CLK _7585_/D _4128_/B VGND VGND VPWR VPWR _7585_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_66 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6552__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _5260_/A _4797_/B _5107_/C VGND VGND VPWR VPWR _4797_/X sky130_fd_sc_hd__and3_1
XANTENNA_77 _3642_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5760__A0 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 input72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ _7466_/Q _6042_/X _6771_/A3 _6446_/X _7522_/Q VGND VGND VPWR VPWR _6536_/X
+ sky130_fd_sc_hd__a32o_1
X_3748_ _7354_/Q _3506_/X _5776_/A _7386_/Q _3738_/X VGND VGND VPWR VPWR _3748_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_119_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6467_ _6467_/A _6600_/B _6468_/C VGND VGND VPWR VPWR _6467_/X sky130_fd_sc_hd__and3_4
X_3679_ _7191_/Q _4551_/A _4515_/B _4539_/C _3678_/X VGND VGND VPWR VPWR _3679_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_161_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5532_/A _5531_/D _5531_/A VGND VGND VPWR VPWR _5491_/A sky130_fd_sc_hd__and3_1
X_6398_ _6383_/X _6385_/X _6397_/Y VGND VGND VPWR VPWR _6398_/X sky130_fd_sc_hd__a21bo_4
Xoutput173 _4176_/X VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
Xoutput184 _3427_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
X_5349_ _5349_/A _5349_/B VGND VGND VPWR VPWR _5355_/A sky130_fd_sc_hd__nor2_1
Xoutput195 _3417_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4740__B_N _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2920 hold2920/A VGND VGND VPWR VPWR _5870_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3405__A _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6419__C _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2931 _7562_/Q VGND VGND VPWR VPWR hold2931/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6607__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2942 _7447_/Q VGND VGND VPWR VPWR hold2942/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2953 _7144_/Q VGND VGND VPWR VPWR hold2953/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5815__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2964 hold2964/A VGND VGND VPWR VPWR hold2964/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2975 hold2975/A VGND VGND VPWR VPWR hold2975/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7019_ _7210_/CLK _7019_/D fanout701/X VGND VGND VPWR VPWR _7019_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2986 _6975_/Q VGND VGND VPWR VPWR _4283_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2997 _6993_/Q VGND VGND VPWR VPWR _4310_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_46_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3841__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input103_A wb_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5766__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6543__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4306__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4609__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5806__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5019__C1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3832__A3 hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6231__B2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6782__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3596__A2 _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4720_ _4836_/C _5079_/B VGND VGND VPWR VPWR _4720_/Y sky130_fd_sc_hd__nand2_4
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4651_ _4591_/Y _4648_/A _4726_/B VGND VGND VPWR VPWR _4948_/B sky130_fd_sc_hd__o21ai_4
XFILLER_30_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6080__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6534__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR _3930_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3602_ _7241_/Q _5612_/B _5632_/B _5686_/A _7309_/Q VGND VGND VPWR VPWR _3602_/X
+ sky130_fd_sc_hd__a32o_4
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_9_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4582_ _4879_/D _4747_/B _4887_/B _4945_/A VGND VGND VPWR VPWR _4583_/B sky130_fd_sc_hd__nand4_4
X_7370_ _7575_/CLK _7370_/D fanout734/X VGND VGND VPWR VPWR _7370_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_128_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__buf_2
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__buf_2
Xhold804 hold804/A VGND VGND VPWR VPWR _7308_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput75 porb VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6321_ _7022_/Q _6070_/X _6110_/X _7173_/Q _6320_/X VGND VGND VPWR VPWR _6327_/B
+ sky130_fd_sc_hd__a221o_1
X_3533_ input60/X _4431_/A _5965_/A _3531_/X _7342_/Q VGND VGND VPWR VPWR _3533_/X
+ sky130_fd_sc_hd__a32o_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR _4129_/B sky130_fd_sc_hd__buf_4
Xhold815 hold815/A VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold826 _4513_/X VGND VGND VPWR VPWR _7165_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap534 _5402_/B1 VGND VGND VPWR VPWR _5580_/A2 sky130_fd_sc_hd__clkbuf_2
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__clkbuf_2
Xhold837 hold837/A VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold848 hold848/A VGND VGND VPWR VPWR _7413_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6252_ _7413_/Q _6119_/D _6116_/C _6136_/C VGND VGND VPWR VPWR _6252_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6298__B2 _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold859 hold859/A VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3464_ _3504_/B _3504_/A VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5203_ _5203_/A _5203_/B _5203_/C _5339_/D VGND VGND VPWR VPWR _5203_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__7096__RESET_B fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6183_ _7386_/Q _6109_/X _6110_/X _7434_/Q _6182_/X VGND VGND VPWR VPWR _6183_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_130_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2205 hold523/X VGND VGND VPWR VPWR _4211_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2216 hold563/X VGND VGND VPWR VPWR _5721_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5134_ _5134_/A _5260_/C _5134_/C VGND VGND VPWR VPWR _5134_/X sky130_fd_sc_hd__and3_1
Xhold2227 _7457_/Q VGND VGND VPWR VPWR hold633/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2238 hold643/X VGND VGND VPWR VPWR _5662_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1504 _5872_/X VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2249 hold619/X VGND VGND VPWR VPWR _5771_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1515 hold220/X VGND VGND VPWR VPWR _5989_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1526 _5980_/X VGND VGND VPWR VPWR hold256/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1537 hold201/X VGND VGND VPWR VPWR _7548_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5065_ _5065_/A _5453_/C VGND VGND VPWR VPWR _5065_/Y sky130_fd_sc_hd__nand2_2
Xhold1548 _7092_/Q VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3808__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1559 _4437_/X VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4016_ _6905_/Q _6904_/Q _4025_/B VGND VGND VPWR VPWR _4017_/B sky130_fd_sc_hd__and3_1
XANTENNA__6470__A1 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5273__A2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3598__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5967_ _5967_/A0 _5994_/A1 _5973_/S VGND VGND VPWR VPWR _5967_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4233__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5981__A0 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4918_ _5213_/A _4997_/B _4924_/B _4918_/D VGND VGND VPWR VPWR _4919_/C sky130_fd_sc_hd__nand4_1
X_5898_ _5997_/A1 _5898_/A1 _5901_/S VGND VGND VPWR VPWR _5898_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6702__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7637_ _7641_/CLK _7637_/D fanout751/X VGND VGND VPWR VPWR _7637_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4503__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6525__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4849_ _5203_/A _4850_/B _5029_/A VGND VGND VPWR VPWR _4849_/X sky130_fd_sc_hd__and3_1
XFILLER_138_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4768__A_N _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7568_ _7572_/CLK _7568_/D fanout733/X VGND VGND VPWR VPWR _7568_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6519_ _7457_/Q _6455_/X _6463_/X _7425_/Q _6518_/X VGND VGND VPWR VPWR _6519_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_134_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7499_ _7542_/CLK _7499_/D fanout709/X VGND VGND VPWR VPWR _7499_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6289__A1 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2750 hold965/X VGND VGND VPWR VPWR _5999_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2761 _7255_/Q VGND VGND VPWR VPWR hold779/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2772 _7155_/Q VGND VGND VPWR VPWR hold963/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2783 _7120_/Q VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2794 hold889/X VGND VGND VPWR VPWR _4380_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4472__A0 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6213__A1 _7283_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6764__A2 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6516__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3443__2 _3443__2/A VGND VGND VPWR VPWR _6823_/A3 sky130_fd_sc_hd__inv_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5255__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6075__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3805__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6790__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6870_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6870_/X sky130_fd_sc_hd__and2_1
XFILLER_90_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6204__A1 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5821_ hold32/X _5965_/B hold26/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__and3_1
XANTENNA__6755__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4215__B1 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5752_ _5752_/A0 _5815_/A1 _5757_/S VGND VGND VPWR VPWR _5752_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4910__A_N _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4604__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4703_ _5399_/B _5072_/B VGND VGND VPWR VPWR _4703_/Y sky130_fd_sc_hd__nand2_2
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3865__D _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5683_ _5683_/A0 _5953_/A1 _5685_/S VGND VGND VPWR VPWR _5683_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6507__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5715__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7422_ _7478_/CLK _7422_/D fanout714/X VGND VGND VPWR VPWR _7422_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4518__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _4879_/D _4747_/B _4887_/B _4945_/A _4805_/B VGND VGND VPWR VPWR _4733_/B
+ sky130_fd_sc_hd__a41o_4
XFILLER_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3726__C1 _3725_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4565_ _4565_/A _4565_/B VGND VGND VPWR VPWR _4585_/A sky130_fd_sc_hd__nor2_2
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7353_ _7421_/CLK _7353_/D fanout716/X VGND VGND VPWR VPWR _7353_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5191__A1 _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold612 _5624_/X VGND VGND VPWR VPWR _7250_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4977__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold623 hold623/A VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold634 hold634/A VGND VGND VPWR VPWR _7457_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6304_ _6289_/X _6291_/X _6303_/Y VGND VGND VPWR VPWR _6304_/X sky130_fd_sc_hd__a21bo_2
XFILLER_116_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3741__A2 _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3516_ _5938_/A _4455_/A _5992_/C VGND VGND VPWR VPWR _5974_/A sky130_fd_sc_hd__and3_4
Xhold656 hold656/A VGND VGND VPWR VPWR _7507_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7284_ _7309_/CLK _7284_/D fanout710/X VGND VGND VPWR VPWR _7284_/Q sky130_fd_sc_hd__dfrtp_4
X_4496_ _4496_/A0 _5853_/A0 _4496_/S VGND VGND VPWR VPWR _4496_/X sky130_fd_sc_hd__mux2_1
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold678 hold678/A VGND VGND VPWR VPWR _7040_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6235_ _7284_/Q _6036_/Y _6067_/A VGND VGND VPWR VPWR _6235_/X sky130_fd_sc_hd__o21a_1
Xhold689 hold689/A VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3447_ _6904_/Q _4025_/A VGND VGND VPWR VPWR _3447_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6140__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2002 hold411/X VGND VGND VPWR VPWR _5779_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2013 hold409/X VGND VGND VPWR VPWR _5711_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5494__A2 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2024 _7410_/Q VGND VGND VPWR VPWR hold441/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2035 _7096_/Q VGND VGND VPWR VPWR hold304/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6166_ _7345_/Q _6070_/X _6072_/X _7417_/Q _6165_/X VGND VGND VPWR VPWR _6166_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_69_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2046 hold451/X VGND VGND VPWR VPWR _4372_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1301 hold3095/X VGND VGND VPWR VPWR hold3096/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1312 hold3187/X VGND VGND VPWR VPWR _7248_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2057 hold439/X VGND VGND VPWR VPWR _5972_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 hold3196/X VGND VGND VPWR VPWR hold3197/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2068 hold473/X VGND VGND VPWR VPWR _5824_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5117_ _4826_/Y _4832_/Y _5528_/A3 _5116_/X _5112_/X VGND VGND VPWR VPWR _5117_/Y
+ sky130_fd_sc_hd__o311ai_2
Xhold2079 hold469/X VGND VGND VPWR VPWR _5808_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1334 hold3215/X VGND VGND VPWR VPWR _7177_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6097_ _6317_/B _6097_/B _6097_/C VGND VGND VPWR VPWR _6097_/X sky130_fd_sc_hd__and3_4
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1345 hold3198/X VGND VGND VPWR VPWR hold3199/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout568_A _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5246__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1356 _4315_/B VGND VGND VPWR VPWR hold3012/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5048_ _5339_/D _5183_/A _5183_/B _5049_/C VGND VGND VPWR VPWR _5051_/B sky130_fd_sc_hd__nand4_1
Xhold1367 _4287_/A1 VGND VGND VPWR VPWR hold3031/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1378 _4317_/B VGND VGND VPWR VPWR hold3116/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1389 hold2084/X VGND VGND VPWR VPWR hold2085/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6999_ _6999_/CLK _6999_/D VGND VGND VPWR VPWR _6999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6746__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4757__A1 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1752_A _7298_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5706__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input170_A wb_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6131__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input31_A mask_rev_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3270 _7214_/Q VGND VGND VPWR VPWR _3997_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_49_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3281 _7104_/Q VGND VGND VPWR VPWR _4425_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3292 _6215_/X VGND VGND VPWR VPWR _7606_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2580 hold731/X VGND VGND VPWR VPWR _4472_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2591 _7461_/Q VGND VGND VPWR VPWR hold827/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1890 hold178/X VGND VGND VPWR VPWR _5712_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3799__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6198__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6737__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5173__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6370__B1 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4350_ _4350_/A0 _5625_/A1 _4351_/S VGND VGND VPWR VPWR _4350_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4281_ _4289_/S _4281_/B VGND VGND VPWR VPWR _4281_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6673__A1 _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6020_ _6067_/B _6019_/Y _7588_/Q VGND VGND VPWR VPWR _7588_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3487__A1 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3503__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6922_ _7264_/CLK _6922_/D fanout688/X VGND VGND VPWR VPWR _6922_/Q sky130_fd_sc_hd__dfstp_4
X_6853_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6853_/X sky130_fd_sc_hd__and2_1
XFILLER_23_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6728__A2 _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5936__A0 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5804_ _5804_/A0 _5948_/A1 _5811_/S VGND VGND VPWR VPWR _5804_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4334__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6784_ _6792_/S _6784_/B VGND VGND VPWR VPWR _6784_/Y sky130_fd_sc_hd__nand2_1
X_3996_ _3996_/A _3996_/B VGND VGND VPWR VPWR _3996_/Y sky130_fd_sc_hd__nor2_1
X_5735_ _5735_/A0 _5951_/A1 _5739_/S VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5864__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3962__A2 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5666_ _5666_/A0 _5954_/A1 _5667_/S VGND VGND VPWR VPWR _5666_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_1_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7405_ _7582_/CLK _7405_/D fanout717/X VGND VGND VPWR VPWR _7405_/Q sky130_fd_sc_hd__dfrtp_4
X_4617_ _4570_/Y _4608_/Y _4767_/A VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__o21bai_4
XANTENNA__6361__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5597_ _5597_/A0 _5732_/A1 _5602_/S VGND VGND VPWR VPWR _5597_/X sky130_fd_sc_hd__mux2_1
Xhold420 hold420/A VGND VGND VPWR VPWR _7561_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7336_ _7542_/CLK _7336_/D fanout708/X VGND VGND VPWR VPWR _7336_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3714__A2 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold431 hold431/A VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4548_ _4548_/A0 _4548_/A1 _4550_/S VGND VGND VPWR VPWR _4548_/X sky130_fd_sc_hd__mux2_1
Xhold442 _5807_/X VGND VGND VPWR VPWR _7410_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold464 _4493_/X VGND VGND VPWR VPWR _7148_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6113__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold475 hold475/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7267_ _7267_/CLK _7267_/D fanout748/X VGND VGND VPWR VPWR _7670_/A sky130_fd_sc_hd__dfrtp_1
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4479_ _4479_/A _4521_/B _4551_/D VGND VGND VPWR VPWR _4484_/S sky130_fd_sc_hd__and3_4
Xhold497 hold497/A VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6664__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6218_ _7412_/Q _6119_/D _6116_/C _6136_/C VGND VGND VPWR VPWR _6218_/X sky130_fd_sc_hd__o211a_1
X_7198_ _7201_/CLK _7198_/D fanout726/X VGND VGND VPWR VPWR _7198_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5612__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ _7529_/Q _6092_/X _6120_/X _7337_/Q _6148_/X VGND VGND VPWR VPWR _6149_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4509__A _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1120 _4359_/X VGND VGND VPWR VPWR _7031_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3413__A _7538_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6427__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1131 hold3111/X VGND VGND VPWR VPWR hold3112/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 _4492_/X VGND VGND VPWR VPWR _7147_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1153 _5912_/X VGND VGND VPWR VPWR _7503_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1164 hold3168/X VGND VGND VPWR VPWR hold3169/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1175 hold2845/X VGND VGND VPWR VPWR hold2846/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _4534_/X VGND VGND VPWR VPWR _7182_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1197 hold2855/X VGND VGND VPWR VPWR hold2856/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6719__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5927__A0 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5059__B _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5774__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input79_A spi_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6104__B1 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output235_A _4147_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3641__B2 _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3850_ input22/X _3488_/X _3542_/X _6921_/Q VGND VGND VPWR VPWR _3850_/X sky130_fd_sc_hd__a22o_2
XANTENNA__6072__C _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3781_ _7410_/Q _4364_/A _3590_/C _3780_/X VGND VGND VPWR VPWR _3782_/D sky130_fd_sc_hd__a31o_1
XANTENNA__6591__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5520_ _5521_/A _5521_/B _5521_/D VGND VGND VPWR VPWR _5520_/Y sky130_fd_sc_hd__nand3_1
X_5451_ _4705_/Y _4720_/Y _5509_/A3 _5448_/D _5223_/C VGND VGND VPWR VPWR _5508_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_172_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4601__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4402_ _4402_/A0 hold198/X _4405_/S VGND VGND VPWR VPWR _4402_/X sky130_fd_sc_hd__mux2_1
X_5382_ _4605_/Y _5563_/A1 _4971_/X _5265_/A _5381_/X VGND VGND VPWR VPWR _5382_/X
+ sky130_fd_sc_hd__o311a_1
X_7121_ _7197_/CLK _7121_/D fanout742/X VGND VGND VPWR VPWR _7121_/Q sky130_fd_sc_hd__dfstp_2
X_4333_ _4333_/A0 _4544_/A1 _4333_/S VGND VGND VPWR VPWR _4333_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5713__A _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4264_ _4264_/A0 _5736_/A1 _4264_/S VGND VGND VPWR VPWR _4264_/X sky130_fd_sc_hd__mux2_1
X_7052_ _7176_/CLK _7052_/D fanout723/X VGND VGND VPWR VPWR _7052_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6003_ _6932_/Q _6009_/B _6019_/A _4117_/Y VGND VGND VPWR VPWR _6006_/A sky130_fd_sc_hd__o31ai_4
X_4195_ _4195_/A0 _5625_/A1 _4202_/S VGND VGND VPWR VPWR _4195_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5859__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2984_A _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5082__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5621__A2 _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _7075_/CLK _6905_/D _6855_/X VGND VGND VPWR VPWR _6905_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5909__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6836_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6836_/X sky130_fd_sc_hd__and2_1
XANTENNA__5385__A1 _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6582__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6767_ _7030_/Q _6459_/B _6459_/C _6462_/X _7035_/Q VGND VGND VPWR VPWR _6767_/X
+ sky130_fd_sc_hd__a32o_1
X_3979_ _7439_/Q _3520_/X _3932_/X _3977_/X _3978_/X VGND VGND VPWR VPWR _3988_/C
+ sky130_fd_sc_hd__a2111o_1
X_5718_ _5736_/A1 _5718_/A1 _5721_/S VGND VGND VPWR VPWR _5718_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3935__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ _6682_/X _6698_/B _6698_/C VGND VGND VPWR VPWR _6698_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_136_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5649_ _5980_/A0 _5649_/A1 _5649_/S VGND VGND VPWR VPWR _5649_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6334__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _3563_/C VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__buf_2
X_7319_ _7542_/CLK _7319_/D fanout708/X VGND VGND VPWR VPWR _7319_/Q sky130_fd_sc_hd__dfstp_4
Xhold261 _6950_/Q VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold272 hold272/A VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold283 hold283/A VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6637__A1 _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout730 fanout750/X VGND VGND VPWR VPWR fanout730/X sky130_fd_sc_hd__buf_6
Xfanout741 fanout749/X VGND VGND VPWR VPWR fanout741/X sky130_fd_sc_hd__buf_8
XFILLER_132_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4884__D _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5342__B _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout752 input164/X VGND VGND VPWR VPWR _6780_/B sky130_fd_sc_hd__buf_12
Xfanout763 input125/X VGND VGND VPWR VPWR _4805_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_58_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout774 _4887_/D VGND VGND VPWR VPWR _5058_/D sky130_fd_sc_hd__clkbuf_16
XANTENNA_input133_A wb_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_828 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3871__A1 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5769__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3926__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6325__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output185_A _3426_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6628__A1 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2029_A _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__buf_2
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6800__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4406__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4951_ _4853_/Y _4936_/Y _4950_/Y _4681_/Y _4949_/Y VGND VGND VPWR VPWR _4958_/A
+ sky130_fd_sc_hd__o2111a_1
X_3902_ _7255_/Q _4265_/B _4364_/B _4340_/A _7017_/Q VGND VGND VPWR VPWR _3902_/X
+ sky130_fd_sc_hd__a32o_1
X_7670_ _7670_/A VGND VGND VPWR VPWR _7670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4882_ _4997_/B _4918_/D VGND VGND VPWR VPWR _4882_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ _7469_/Q _6434_/X _6616_/X _6617_/X _6620_/X VGND VGND VPWR VPWR _6621_/X
+ sky130_fd_sc_hd__a2111o_1
X_3833_ _7537_/Q _3492_/X _5947_/B _3675_/X _7189_/Q VGND VGND VPWR VPWR _3837_/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6564__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3917__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6552_ _7427_/Q _6463_/X _6467_/X _7419_/Q VGND VGND VPWR VPWR _6552_/X sky130_fd_sc_hd__a22o_1
X_3764_ input14/X _3490_/X _3760_/X _3761_/X _3763_/X VGND VGND VPWR VPWR _3764_/X
+ sky130_fd_sc_hd__a2111o_4
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5503_ _4672_/X _4873_/X _4893_/Y _5340_/D _5438_/C VGND VGND VPWR VPWR _5550_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5119__A1 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6316__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6483_ _7352_/Q _6561_/A2 _6459_/C _6462_/X _7360_/Q VGND VGND VPWR VPWR _6483_/X
+ sky130_fd_sc_hd__a32o_1
X_3695_ _7467_/Q _3565_/X _3692_/X _3694_/X VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__a211o_1
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput300 _4173_/X VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
X_5434_ _4996_/A _5329_/X _5426_/X _5053_/C _5191_/X VGND VGND VPWR VPWR _5501_/A
+ sky130_fd_sc_hd__a221o_1
X_7599__777 VGND VGND VPWR VPWR _7599_/D _7599__777/LO sky130_fd_sc_hd__conb_1
Xoutput311 _7628_/Q VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
XFILLER_133_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput322 hold1111/X VGND VGND VPWR VPWR hold1112/A sky130_fd_sc_hd__buf_6
Xoutput333 hold1156/X VGND VGND VPWR VPWR hold1157/A sky130_fd_sc_hd__buf_6
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5365_ _4601_/Y _4947_/Y _4949_/A VGND VGND VPWR VPWR _5367_/D sky130_fd_sc_hd__o21bai_2
XFILLER_160_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR _7399_/CLK sky130_fd_sc_hd__clkbuf_8
X_7104_ _7111_/CLK _7104_/D _6780_/B VGND VGND VPWR VPWR _7104_/Q sky130_fd_sc_hd__dfrtp_4
X_4316_ _4321_/S _3795_/B _4315_/Y VGND VGND VPWR VPWR _6996_/D sky130_fd_sc_hd__o21ai_1
X_5296_ _4720_/Y _4755_/Y _4761_/Y _4692_/Y _5143_/A VGND VGND VPWR VPWR _5303_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7035_ _7035_/CLK _7035_/D fanout723/X VGND VGND VPWR VPWR _7035_/Q sky130_fd_sc_hd__dfrtp_4
X_4247_ _4247_/A0 _4246_/X _4249_/S VGND VGND VPWR VPWR _4247_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout383_A _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4178_ _4178_/A _4427_/D VGND VGND VPWR VPWR _7102_/D sky130_fd_sc_hd__and2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout550_A _4446_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6252__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3605__A1 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1498_A _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6819_ _6818_/X _6819_/A1 _6822_/S VGND VGND VPWR VPWR _7643_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6555__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3908__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4879__D _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5530__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5072__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout560 _5726_/A1 VGND VGND VPWR VPWR _5647_/A0 sky130_fd_sc_hd__buf_4
XFILLER_59_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout571 _5635_/A0 VGND VGND VPWR VPWR _5968_/A1 sky130_fd_sc_hd__buf_6
XFILLER_76_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout582 hold1567/X VGND VGND VPWR VPWR _5922_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout593 hold26/X VGND VGND VPWR VPWR _5619_/C sky130_fd_sc_hd__buf_12
XFILLER_19_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3844__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5597__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6561__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ _3504_/A hold88/X VGND VGND VPWR VPWR _3647_/A sky130_fd_sc_hd__and2_1
XANTENNA__6313__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2146_A _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5150_ _5150_/A _5150_/B _5150_/C VGND VGND VPWR VPWR _5153_/A sky130_fd_sc_hd__and3_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2409 hold697/X VGND VGND VPWR VPWR _4327_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4101_ _6429_/C _7594_/Q VGND VGND VPWR VPWR _4101_/X sky130_fd_sc_hd__and2b_4
XANTENNA__6077__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5081_ _5081_/A _5387_/D _5260_/C _5091_/A VGND VGND VPWR VPWR _5081_/Y sky130_fd_sc_hd__nand4_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1708 _7486_/Q VGND VGND VPWR VPWR hold95/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1719 hold332/X VGND VGND VPWR VPWR _5751_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4032_ _6903_/Q _4025_/A _4030_/Y _4031_/X VGND VGND VPWR VPWR _4032_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_5_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5588__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5983_ _5983_/A _5992_/C _5992_/D VGND VGND VPWR VPWR _5991_/S sky130_fd_sc_hd__and3_4
XFILLER_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3599__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4934_ _4934_/A _4934_/B _4934_/C VGND VGND VPWR VPWR _4934_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4260__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7653_ _7653_/A VGND VGND VPWR VPWR _7653_/X sky130_fd_sc_hd__buf_2
X_4865_ _5183_/A _5053_/C VGND VGND VPWR VPWR _4865_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6537__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _3961_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_23 _6665_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6604_ _7373_/Q _6413_/C _6651_/C _6603_/X VGND VGND VPWR VPWR _6604_/X sky130_fd_sc_hd__a31o_1
X_3816_ _7179_/Q _5947_/B _5619_/B _7401_/Q _5794_/A VGND VGND VPWR VPWR _3816_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_45 input91/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7584_ _7601_/CLK _7584_/D _4128_/B VGND VGND VPWR VPWR _7584_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_56 _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ _5260_/A _4797_/B VGND VGND VPWR VPWR _4796_/Y sky130_fd_sc_hd__nand2_4
XANTENNA_67 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _3642_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_89 wire350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6535_ _7298_/Q _6420_/A _6530_/X _6532_/X _6534_/X VGND VGND VPWR VPWR _6545_/B
+ sky130_fd_sc_hd__a2111oi_4
X_3747_ _7185_/Q _4533_/A _3670_/X _7135_/Q _3746_/X VGND VGND VPWR VPWR _3747_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6466_ _6466_/A _6466_/B _6466_/C _6466_/D VGND VGND VPWR VPWR _6466_/X sky130_fd_sc_hd__and4_4
XFILLER_133_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3678_ _7181_/Q _4376_/B _3738_/B _3647_/X _7171_/Q VGND VGND VPWR VPWR _3678_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5417_ _4695_/Y _4732_/Y _5317_/A VGND VGND VPWR VPWR _5532_/A sky130_fd_sc_hd__o21ba_1
X_6397_ _6397_/A _6397_/B _6397_/C _6397_/D VGND VGND VPWR VPWR _6397_/Y sky130_fd_sc_hd__nor4_1
XFILLER_133_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput174 _4177_/X VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ _5094_/A _4939_/C _4907_/B _4954_/C _5213_/B VGND VGND VPWR VPWR _5349_/B
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput185 _3426_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
XFILLER_88_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput196 _3416_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
Xhold2910 _7256_/Q VGND VGND VPWR VPWR hold2910/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6068__A2 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2921 _7361_/Q VGND VGND VPWR VPWR hold2921/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6419__D _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2932 hold2932/A VGND VGND VPWR VPWR _5978_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout765_A _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5279_ _4667_/B _4828_/Y _5278_/X VGND VGND VPWR VPWR _5279_/Y sky130_fd_sc_hd__o21ai_1
Xhold2943 hold2943/A VGND VGND VPWR VPWR _5849_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2954 hold2954/A VGND VGND VPWR VPWR _4488_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ _7164_/CLK _7018_/D fanout702/X VGND VGND VPWR VPWR _7018_/Q sky130_fd_sc_hd__dfstp_1
Xhold2965 hold2965/A VGND VGND VPWR VPWR hold2965/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2976 _6987_/Q VGND VGND VPWR VPWR _4302_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2987 hold2987/A VGND VGND VPWR VPWR hold2987/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2998 hold2998/A VGND VGND VPWR VPWR hold2998/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3421__A _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6435__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold343_A _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6776__B1 _6774_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6240__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4251__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6451__B _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5751__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5782__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3762__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input61_A mgmt_gpio_in[32] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6700__B1 _6698_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5267__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3817__A1 _7281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout390 _5632_/B VGND VGND VPWR VPWR _4352_/B sky130_fd_sc_hd__buf_8
XFILLER_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4427__A _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6767__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6231__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4242__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6519__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5990__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4650_ _4591_/Y _4648_/A _4726_/B VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__o21a_4
XANTENNA__6080__C _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3601_ _6917_/Q _3527_/X _3597_/X _3598_/X _3600_/X VGND VGND VPWR VPWR _3606_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_163_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR _3863_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5742__A1 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4581_ _4879_/D _4747_/B _4887_/B _4945_/A VGND VGND VPWR VPWR _4581_/X sky130_fd_sc_hd__and4_4
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6320_ _7037_/Q _6082_/C _6388_/A3 _6072_/X _7153_/Q VGND VGND VPWR VPWR _6320_/X
+ sky130_fd_sc_hd__a32o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR _7672_/A sky130_fd_sc_hd__buf_4
X_3532_ _5992_/A _3682_/A _5965_/A VGND VGND VPWR VPWR _3532_/X sky130_fd_sc_hd__and3_1
Xhold805 hold805/A VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 qspi_enabled VGND VGND VPWR VPWR _4142_/A sky130_fd_sc_hd__buf_12
Xhold816 _5862_/X VGND VGND VPWR VPWR _7459_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR _7671_/A sky130_fd_sc_hd__buf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__clkbuf_2
Xhold827 hold827/A VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap535 _4430_/C VGND VGND VPWR VPWR _5402_/B1 sky130_fd_sc_hd__clkbuf_2
XFILLER_171_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold838 hold838/A VGND VGND VPWR VPWR _7437_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6298__A2 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6251_ _7349_/Q _6070_/X _6112_/X _7485_/Q _6250_/X VGND VGND VPWR VPWR _6257_/C
+ sky130_fd_sc_hd__a221o_1
Xhold849 hold849/A VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3463_ _3462_/X _3463_/A1 _4181_/S VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3506__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ _5202_/A _5202_/B _5202_/C VGND VGND VPWR VPWR _5202_/X sky130_fd_sc_hd__and3_1
X_6182_ _7426_/Q _6080_/A _6074_/X _6120_/X _7338_/Q VGND VGND VPWR VPWR _6182_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2206 _7242_/Q VGND VGND VPWR VPWR hold531/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2217 _5721_/X VGND VGND VPWR VPWR hold564/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2228 hold633/X VGND VGND VPWR VPWR _5860_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5133_ _5407_/A1 _5282_/A _5091_/A _5260_/D VGND VGND VPWR VPWR _5134_/C sky130_fd_sc_hd__a31o_2
XFILLER_111_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2239 _5662_/X VGND VGND VPWR VPWR hold644/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1505 hold260/X VGND VGND VPWR VPWR _7468_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1516 _5989_/X VGND VGND VPWR VPWR hold221/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1527 _7508_/Q VGND VGND VPWR VPWR hold310/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5064_ _5064_/A _5064_/B _5064_/C VGND VGND VPWR VPWR _5064_/Y sky130_fd_sc_hd__nand3_1
Xhold1538 _7524_/Q VGND VGND VPWR VPWR hold224/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1549 hold58/X VGND VGND VPWR VPWR _4439_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4015_ _6903_/Q _6902_/Q _6901_/Q _6900_/Q VGND VGND VPWR VPWR _4025_/B sky130_fd_sc_hd__and4_2
XANTENNA__6470__A2 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4481__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5966_ _5966_/A0 _5993_/A1 _5973_/S VGND VGND VPWR VPWR _5966_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4233__A1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5430__B1 _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4917_ _5213_/A _5213_/B _4924_/B _4970_/C VGND VGND VPWR VPWR _5573_/C sky130_fd_sc_hd__nand4_2
XFILLER_178_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5897_ _5978_/A0 _5897_/A1 _5901_/S VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7636_ _7636_/CLK _7636_/D VGND VGND VPWR VPWR _7636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4848_ wire375/X _4850_/B _5203_/C _4847_/X VGND VGND VPWR VPWR _4851_/B sky130_fd_sc_hd__a31oi_1
XFILLER_178_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6525__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5733__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7567_ _7573_/CLK _7567_/D fanout733/X VGND VGND VPWR VPWR _7567_/Q sky130_fd_sc_hd__dfstp_1
X_4779_ _4700_/Y _4774_/Y _4778_/Y _4776_/Y VGND VGND VPWR VPWR _4781_/B sky130_fd_sc_hd__o211ai_1
XFILLER_119_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6518_ _7393_/Q _6420_/C _6467_/X _7417_/Q _6517_/X VGND VGND VPWR VPWR _6518_/X
+ sky130_fd_sc_hd__a221o_1
X_7498_ _7514_/CLK _7498_/D fanout743/X VGND VGND VPWR VPWR _7498_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6289__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6449_ _7311_/Q _6419_/D _6425_/X _7335_/Q _6448_/X VGND VGND VPWR VPWR _6449_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3416__A _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1530_A _7436_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7551_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5631__A _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2740 hold765/X VGND VGND VPWR VPWR _5589_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2751 _5999_/X VGND VGND VPWR VPWR hold966/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2762 hold779/X VGND VGND VPWR VPWR _5629_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2773 hold963/X VGND VGND VPWR VPWR _4501_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2784 hold977/X VGND VGND VPWR VPWR _4459_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_55_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7314_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6461__A2 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2795 _4380_/X VGND VGND VPWR VPWR hold890/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5777__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6213__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5972__A1 _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3378_A _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5724__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6401__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4710__A _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__B1 _4159_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6906__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4463__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6075__C _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6204__A2 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5820_ _5820_/A0 _6000_/A1 _5820_/S VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5751_ _5751_/A0 _5949_/A1 _5757_/S VGND VGND VPWR VPWR _5751_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5963__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4604__B _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3974__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4702_ _4910_/D _4856_/A _4888_/B _5282_/A VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__nor4_4
X_5682_ _5682_/A0 _5952_/A1 _5685_/S VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7421_ _7421_/CLK _7421_/D fanout716/X VGND VGND VPWR VPWR _7421_/Q sky130_fd_sc_hd__dfrtp_2
X_4633_ _4768_/B _4641_/A VGND VGND VPWR VPWR _4802_/A sky130_fd_sc_hd__nor2_4
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7352_ _7563_/CLK _7352_/D fanout739/X VGND VGND VPWR VPWR _7352_/Q sky130_fd_sc_hd__dfstp_4
X_4564_ _4564_/A _4564_/B _4564_/C _4564_/D VGND VGND VPWR VPWR _4565_/B sky130_fd_sc_hd__nand4_1
XANTENNA__5191__A2 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold602 hold602/A VGND VGND VPWR VPWR _7406_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold613 hold613/A VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6303_ _6303_/A _6303_/B _6303_/C _6303_/D VGND VGND VPWR VPWR _6303_/Y sky130_fd_sc_hd__nor4_1
Xhold624 _5871_/X VGND VGND VPWR VPWR _7467_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3515_ _5640_/B _3598_/B _4388_/B VGND VGND VPWR VPWR _3515_/X sky130_fd_sc_hd__and3_4
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7283_ _7309_/CLK _7283_/D fanout704/X VGND VGND VPWR VPWR _7283_/Q sky130_fd_sc_hd__dfrtp_4
Xhold646 _5878_/X VGND VGND VPWR VPWR _7473_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4495_ _4495_/A0 _4555_/A0 _4496_/S VGND VGND VPWR VPWR _4495_/X sky130_fd_sc_hd__mux2_1
Xhold657 hold657/A VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold668 hold668/A VGND VGND VPWR VPWR _6952_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap376 _4836_/A VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__clkbuf_2
X_6234_ _6228_/X _6230_/X _6231_/X _6233_/X VGND VGND VPWR VPWR _6234_/X sky130_fd_sc_hd__a211o_1
Xhold679 hold679/A VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3446_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _3856_/A sky130_fd_sc_hd__nor3_4
XANTENNA__6140__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2003 _5779_/X VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6691__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _7497_/Q _6332_/B _6388_/A3 _6100_/X _7473_/Q VGND VGND VPWR VPWR _6165_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2014 _5711_/X VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2025 hold441/X VGND VGND VPWR VPWR _5807_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2036 hold304/X VGND VGND VPWR VPWR _4444_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4993__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2047 _4372_/X VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 hold3097/X VGND VGND VPWR VPWR _7263_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1313 hold3171/X VGND VGND VPWR VPWR hold3172/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5116_ _5480_/B2 _4826_/Y _4832_/Y _4828_/Y _5480_/A1 VGND VGND VPWR VPWR _5116_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2058 _7552_/Q VGND VGND VPWR VPWR hold503/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2069 _7408_/Q VGND VGND VPWR VPWR hold2069/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1324 _4395_/X VGND VGND VPWR VPWR _7061_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6096_ _7375_/Q _6090_/X _6092_/X _7527_/Q _6095_/X VGND VGND VPWR VPWR _6102_/C
+ sky130_fd_sc_hd__a221o_1
Xhold1335 hold3230/X VGND VGND VPWR VPWR hold3231/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1346 hold3200/X VGND VGND VPWR VPWR _6962_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1357 _4310_/B VGND VGND VPWR VPWR hold2998/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5246__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5047_ _5047_/A _5047_/B _5047_/C VGND VGND VPWR VPWR _5051_/A sky130_fd_sc_hd__nor3_1
Xhold1368 _4283_/B VGND VGND VPWR VPWR hold2987/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5651__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1379 _4285_/B VGND VGND VPWR VPWR hold3220/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4454__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4206__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6998_ _6999_/CLK _6998_/D VGND VGND VPWR VPWR _6998_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout728_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6746__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5954__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5949_ _5949_/A0 _5949_/A1 _5955_/S VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7619_ _7625_/CLK _7619_/D fanout705/X VGND VGND VPWR VPWR _7619_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5048__D _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4390__A0 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4887__D _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1912_A _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input163_A wb_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6131__A1 _7408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6682__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3260 hold3260/A VGND VGND VPWR VPWR _4192_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3271 _7220_/Q VGND VGND VPWR VPWR _3609_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3282 _7106_/Q VGND VGND VPWR VPWR _4425_/C sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3293 _7623_/Q VGND VGND VPWR VPWR _6700_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2570 _4378_/X VGND VGND VPWR VPWR hold936/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input24_A mask_rev_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2581 _4472_/X VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2592 hold827/X VGND VGND VPWR VPWR _5864_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4445__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1880 _7494_/Q VGND VGND VPWR VPWR hold134/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1891 _5712_/X VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3799__A3 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6198__A1 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5945__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5173__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3723__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5970__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4280_ _3922_/Y _4280_/A1 _4289_/S VGND VGND VPWR VPWR _6973_/D sky130_fd_sc_hd__mux2_1
XFILLER_152_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4133__A0 input85/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6673__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3487__A2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3503__B _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4436__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6921_ _7255_/CLK _6921_/D fanout688/X VGND VGND VPWR VPWR _6921_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_54_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6852_ _6872_/A _6872_/B VGND VGND VPWR VPWR _6852_/X sky130_fd_sc_hd__and2_1
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6728__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5803_ _5803_/A _5947_/A _5893_/B VGND VGND VPWR VPWR _5811_/S sky130_fd_sc_hd__and3_4
X_6783_ _3922_/Y _6783_/A1 _6792_/S VGND VGND VPWR VPWR _7630_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4334__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3995_ _3926_/X _3995_/B _3995_/C _3995_/D VGND VGND VPWR VPWR _3996_/B sky130_fd_sc_hd__and4b_4
XANTENNA__3947__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5734_ _5734_/A0 _5950_/A1 _5739_/S VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5665_ _5665_/A0 _5953_/A1 _5667_/S VGND VGND VPWR VPWR _5665_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3962__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7404_ _7541_/CLK _7404_/D fanout711/X VGND VGND VPWR VPWR _7404_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4616_ _4643_/C _4645_/D VGND VGND VPWR VPWR _4616_/Y sky130_fd_sc_hd__nand2_2
XFILLER_191_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5596_ _5596_/A _5596_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5602_/S sky130_fd_sc_hd__and4_4
XANTENNA__6361__B2 _6991_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4372__A0 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold410 hold410/A VGND VGND VPWR VPWR _7325_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7335_ _7539_/CLK _7335_/D fanout707/X VGND VGND VPWR VPWR _7335_/Q sky130_fd_sc_hd__dfstp_2
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4547_ _4547_/A0 _4547_/A1 _4550_/S VGND VGND VPWR VPWR _4547_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3714__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold432 hold432/A VGND VGND VPWR VPWR _7028_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5880__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold443 hold443/A VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_5_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold454 hold454/A VGND VGND VPWR VPWR _6875_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7266_ _7266_/CLK _7266_/D _6864_/A VGND VGND VPWR VPWR _7266_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6113__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6113__B2 _7479_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4478_ _4478_/A0 _5817_/A1 _4478_/S VGND VGND VPWR VPWR _4478_/X sky130_fd_sc_hd__mux2_1
Xhold476 _4535_/X VGND VGND VPWR VPWR _7183_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold487 hold487/A VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__buf_12
XFILLER_143_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold498 hold498/A VGND VGND VPWR VPWR _7312_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6217_ _7460_/Q _6080_/X _6085_/X _7500_/Q _6216_/X VGND VGND VPWR VPWR _6217_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6664__A2 _7117_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3429_ _7410_/Q VGND VGND VPWR VPWR _3429_/Y sky130_fd_sc_hd__clkinv_2
X_7197_ _7197_/CLK _7197_/D fanout741/X VGND VGND VPWR VPWR _7197_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5612__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6148_ _7489_/Q _6112_/C _6276_/A3 _6116_/X _7313_/Q VGND VGND VPWR VPWR _6148_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_100_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1110 hold3134/X VGND VGND VPWR VPWR _7117_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1121 hold3122/X VGND VGND VPWR VPWR hold3123/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1132 _4498_/X VGND VGND VPWR VPWR _7152_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 hold3140/X VGND VGND VPWR VPWR hold3141/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ _7588_/Q _6099_/D _6081_/C _7589_/Q VGND VGND VPWR VPWR _6079_/X sky130_fd_sc_hd__and4bb_4
Xhold1154 hold3036/X VGND VGND VPWR VPWR hold1154/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1165 hold3170/X VGND VGND VPWR VPWR _7127_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1176 _4262_/X VGND VGND VPWR VPWR _6959_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1187 hold2921/X VGND VGND VPWR VPWR hold2922/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 hold2857/X VGND VGND VPWR VPWR _6946_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3953__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6352__A1 _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5155__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5790__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6104__A1 _7327_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6104__B2 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__B _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5458__A3 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5863__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3090 _6984_/Q VGND VGND VPWR VPWR _4298_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4418__A1 _4446_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4969__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3641__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5918__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3780_ _7450_/Q _5848_/A _4545_/A _7195_/Q _3779_/X VGND VGND VPWR VPWR _3780_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6591__A1 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6591__B2 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5450_ _5226_/X _5450_/B _5450_/C VGND VGND VPWR VPWR _5574_/A sky130_fd_sc_hd__and3b_1
X_4401_ _4401_/A0 _5582_/A0 _4405_/S VGND VGND VPWR VPWR _4401_/X sky130_fd_sc_hd__mux2_1
X_5381_ _4700_/Y _5563_/A1 _4720_/Y _5081_/Y VGND VGND VPWR VPWR _5381_/X sky130_fd_sc_hd__o31a_1
XFILLER_172_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7120_ _7197_/CLK _7120_/D fanout741/X VGND VGND VPWR VPWR _7120_/Q sky130_fd_sc_hd__dfstp_2
Xclkbuf_3_2_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_4332_ _4332_/A0 _5625_/A1 _4333_/S VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold32_A hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5713__B _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7051_ _7164_/CLK _7051_/D fanout698/X VGND VGND VPWR VPWR _7051_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6646__A2 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4263_ _4263_/A0 _5625_/A1 _4264_/S VGND VGND VPWR VPWR _4263_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2510_A _7201_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3514__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5854__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6002_ _6065_/C _6929_/Q _7256_/Q _6001_/Y _6002_/B2 VGND VGND VPWR VPWR _7583_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4194_ _4194_/A0 _5815_/A1 _4202_/S VGND VGND VPWR VPWR _4194_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3880__A2 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5621__A3 _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6904_ _4150_/A1 _6904_/D _6854_/X VGND VGND VPWR VPWR _6904_/Q sky130_fd_sc_hd__dfrtp_4
X_6835_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6835_/X sky130_fd_sc_hd__and2_1
X_6766_ _7171_/Q _6408_/D _6454_/X _7070_/Q _6765_/X VGND VGND VPWR VPWR _6773_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3978_ _7172_/Q _3931_/B _4364_/B _3649_/X _7066_/Q VGND VGND VPWR VPWR _3978_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_138_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5717_ _5951_/A1 _5717_/A1 _5721_/S VGND VGND VPWR VPWR _5717_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6697_ _6697_/A _6697_/B _6697_/C _6697_/D VGND VGND VPWR VPWR _6698_/C sky130_fd_sc_hd__nor4_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_1__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _7075_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5648_ _5979_/A0 _5648_/A1 _5649_/S VGND VGND VPWR VPWR _5648_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5579_ _5385_/X _5520_/Y _5564_/Y _5578_/Y _5560_/X VGND VGND VPWR VPWR _5579_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_105_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3699__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7318_ _7576_/CLK _7318_/D fanout717/X VGND VGND VPWR VPWR _7318_/Q sky130_fd_sc_hd__dfrtp_4
Xhold240 hold240/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold251 _4303_/X VGND VGND VPWR VPWR _4308_/S sky130_fd_sc_hd__buf_2
XFILLER_116_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold273 hold273/A VGND VGND VPWR VPWR _7100_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold284 hold284/A VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5623__B _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6637__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold295 hold295/A VGND VGND VPWR VPWR _7539_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7249_ _7266_/CLK _7249_/D fanout692/X VGND VGND VPWR VPWR _7648_/A sky130_fd_sc_hd__dfrtp_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout720 fanout750/X VGND VGND VPWR VPWR fanout720/X sky130_fd_sc_hd__buf_12
XANTENNA__3424__A _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout731 fanout736/X VGND VGND VPWR VPWR fanout731/X sky130_fd_sc_hd__buf_8
Xfanout742 fanout749/X VGND VGND VPWR VPWR fanout742/X sky130_fd_sc_hd__clkbuf_8
Xfanout753 input164/X VGND VGND VPWR VPWR fanout753/X sky130_fd_sc_hd__buf_4
Xfanout764 _5407_/A1 VGND VGND VPWR VPWR _4888_/B sky130_fd_sc_hd__buf_12
Xfanout775 _4887_/D VGND VGND VPWR VPWR _4910_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_92_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3871__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input126_A wb_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6454__B _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6270__B1 _6089_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5376__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input91_A spimemio_flash_io3_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3926__A3 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4702__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5086__A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6325__A1 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6325__B2 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6628__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4639__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5300__A2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4950_ _4966_/A _5222_/B _5222_/C _5094_/A VGND VGND VPWR VPWR _4950_/Y sky130_fd_sc_hd__nand4_1
XFILLER_33_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3901_ _7052_/Q _3931_/B _3738_/B _3900_/X VGND VGND VPWR VPWR _3901_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4881_ _4942_/A _4948_/C _4918_/D VGND VGND VPWR VPWR _4943_/B sky130_fd_sc_hd__and3_2
XFILLER_178_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6159__A4 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6620_ _7413_/Q _6468_/X _6618_/X _6619_/X _6430_/X VGND VGND VPWR VPWR _6620_/X
+ sky130_fd_sc_hd__a2111o_1
X_3832_ _7457_/Q _3933_/A hold32/A _3537_/X _7425_/Q VGND VGND VPWR VPWR _3837_/B
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6564__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6551_ _7331_/Q _6423_/X _6452_/X _7347_/Q _6550_/X VGND VGND VPWR VPWR _6551_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3763_ input23/X _3488_/X _3521_/X _7314_/Q _3762_/X VGND VGND VPWR VPWR _3763_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_158_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5502_ _4679_/Y _4832_/Y _5528_/A3 _5438_/B _5200_/B VGND VGND VPWR VPWR _5550_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_192_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_1_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6482_ _7392_/Q _6420_/C _6419_/A _7544_/Q _6481_/X VGND VGND VPWR VPWR _6482_/X
+ sky130_fd_sc_hd__a221o_1
X_3694_ _7020_/Q _4352_/A _5619_/B _3693_/X VGND VGND VPWR VPWR _3694_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6316__B2 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5433_ _5331_/Y _5554_/B _5433_/C VGND VGND VPWR VPWR _5435_/B sky130_fd_sc_hd__nand3b_1
XFILLER_145_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput301 _4117_/B VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 hold1080/X VGND VGND VPWR VPWR hold1081/A sky130_fd_sc_hd__buf_6
XFILLER_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput323 hold1096/X VGND VGND VPWR VPWR hold1097/A sky130_fd_sc_hd__buf_6
Xoutput334 hold1082/X VGND VGND VPWR VPWR hold1083/A sky130_fd_sc_hd__buf_6
X_5364_ _5089_/D _4856_/Y _5248_/C _4935_/X VGND VGND VPWR VPWR _5545_/B sky130_fd_sc_hd__o31a_1
XFILLER_114_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7103_ _7111_/CLK _7103_/D _6780_/B VGND VGND VPWR VPWR _7103_/Q sky130_fd_sc_hd__dfrtp_4
X_4315_ _4321_/S _4315_/B VGND VGND VPWR VPWR _4315_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6619__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5295_ _5295_/A _5295_/B _5404_/D _5295_/D VGND VGND VPWR VPWR _5422_/D sky130_fd_sc_hd__nand4_2
XFILLER_141_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7034_ _7035_/CLK _7034_/D fanout723/X VGND VGND VPWR VPWR _7034_/Q sky130_fd_sc_hd__dfrtp_4
X_4246_ _5657_/A1 _5954_/A1 _4248_/S VGND VGND VPWR VPWR _4246_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6095__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4177_ _7264_/Q _4177_/B VGND VGND VPWR VPWR _4177_/X sky130_fd_sc_hd__and2_2
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6252__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout543_A _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3605__A2 _3486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6818_ _4427_/B _6818_/A2 _6818_/B1 wire536/A _6817_/X VGND VGND VPWR VPWR _6818_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5358__A2 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6749_ _6749_/A _6749_/B _6749_/C _6749_/D VGND VGND VPWR VPWR _6749_/Y sky130_fd_sc_hd__nor4_1
XANTENNA_hold1560_A _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3419__A _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1825_A _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout550 _4446_/A1 VGND VGND VPWR VPWR _5980_/A0 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _5726_/A1 VGND VGND VPWR VPWR _5951_/A1 sky130_fd_sc_hd__buf_6
Xfanout572 _5788_/A1 VGND VGND VPWR VPWR _5914_/A1 sky130_fd_sc_hd__buf_6
XANTENNA__6491__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout583 _5894_/A0 VGND VGND VPWR VPWR _5732_/A1 sky130_fd_sc_hd__buf_6
XFILLER_65_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout594 _5893_/B VGND VGND VPWR VPWR _5947_/C sky130_fd_sc_hd__buf_12
XANTENNA__3844__A2 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output295_A _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3780__A1 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4100_ _7584_/Q _7586_/Q _4100_/A3 _4099_/D _6932_/Q VGND VGND VPWR VPWR _4100_/X
+ sky130_fd_sc_hd__o41a_1
X_5080_ _5563_/A1 _4737_/Y _5516_/A3 _5077_/Y _4748_/Y VGND VGND VPWR VPWR _5084_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1709 hold95/X VGND VGND VPWR VPWR _5892_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5285__A1 _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6482__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4031_ _6903_/Q _6902_/Q _6901_/Q _6900_/Q _6904_/Q VGND VGND VPWR VPWR _4031_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_111_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3835__A2 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6785__A1 _6789_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5982_ _5991_/A1 _5982_/A1 _5982_/S VGND VGND VPWR VPWR _5982_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4933_ _4933_/A _4933_/B _5049_/C VGND VGND VPWR VPWR _4934_/B sky130_fd_sc_hd__and3_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7652_ _7652_/A VGND VGND VPWR VPWR _7652_/X sky130_fd_sc_hd__clkbuf_2
X_4864_ _5328_/A _5328_/B _5053_/C VGND VGND VPWR VPWR _4864_/X sky130_fd_sc_hd__and3_2
XANTENNA__6537__A1 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6537__B2 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_13 _3961_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3815_ _6913_/Q _3527_/X _4340_/A _7018_/Q _3814_/X VGND VGND VPWR VPWR _3815_/X
+ sky130_fd_sc_hd__a221o_1
X_6603_ _7477_/Q _6466_/C _6441_/X _6058_/X _7533_/Q VGND VGND VPWR VPWR _6603_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_24 _6712_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7583_ _7587_/CLK _7583_/D _6864_/A VGND VGND VPWR VPWR _7583_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_35 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _4860_/A _4772_/A _4831_/A _4814_/C VGND VGND VPWR VPWR _4799_/C sky130_fd_sc_hd__and4bb_4
XANTENNA_hold2842_A _6947_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _6922_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ _7538_/Q _6408_/D _6425_/X _7338_/Q _6533_/X VGND VGND VPWR VPWR _6534_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_79 _3714_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ _7394_/Q _4473_/A _5785_/B _3665_/X _7125_/Q VGND VGND VPWR VPWR _3746_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3771__A1 _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6465_ _7303_/Q _6420_/B _6462_/X _7359_/Q _6464_/X VGND VGND VPWR VPWR _6471_/C
+ sky130_fd_sc_hd__a221o_1
X_3677_ _7539_/Q _3590_/C _5947_/B _5893_/A _7491_/Q VGND VGND VPWR VPWR _3677_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_106_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5416_ _5535_/A _5416_/B _5535_/B VGND VGND VPWR VPWR _5419_/B sky130_fd_sc_hd__and3_1
X_6396_ _7025_/Q _6070_/X _6080_/X _7201_/Q _6395_/X VGND VGND VPWR VPWR _6397_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_114_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5347_ _4947_/C _4933_/A _5346_/X _5208_/Y VGND VGND VPWR VPWR _5347_/X sky130_fd_sc_hd__a31o_1
Xoutput175 _4160_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
XFILLER_88_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput186 _4158_/X VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 _3442_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
Xhold2900 _7053_/Q VGND VGND VPWR VPWR hold2900/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2911 hold2911/A VGND VGND VPWR VPWR _5630_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2922 hold2922/A VGND VGND VPWR VPWR _5752_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5278_ _5277_/X _5278_/B _5278_/C _5278_/D VGND VGND VPWR VPWR _5278_/X sky130_fd_sc_hd__and4b_1
Xhold2933 _5978_/X VGND VGND VPWR VPWR hold2933/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2944 _5849_/X VGND VGND VPWR VPWR _7447_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2955 _7194_/Q VGND VGND VPWR VPWR hold2955/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7017_ _7212_/CLK _7017_/D fanout724/X VGND VGND VPWR VPWR _7017_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2966 _7000_/Q VGND VGND VPWR VPWR _4321_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4229_ _4257_/A0 _5990_/A1 _4231_/S VGND VGND VPWR VPWR _4229_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2977 hold2977/A VGND VGND VPWR VPWR hold2977/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout758_A _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3826__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2988 _6998_/Q VGND VGND VPWR VPWR _4319_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2999 _6986_/Q VGND VGND VPWR VPWR _4301_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6225__B1 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6240__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6528__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6451__C _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3762__A1 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3762__B2 _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A mgmt_gpio_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6464__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout380 _6872_/B VGND VGND VPWR VPWR _6869_/B sky130_fd_sc_hd__buf_4
XANTENNA__4708__A _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3817__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout391 _3514_/X VGND VGND VPWR VPWR _5632_/B sky130_fd_sc_hd__buf_12
XANTENNA__4427__B _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6216__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output308_A _4135_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6767__A1 _7030_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5973__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3600_ _7341_/Q _3531_/X _3545_/X _7349_/Q _3599_/X VGND VGND VPWR VPWR _3600_/X
+ sky130_fd_sc_hd__a221o_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4580_ _4831_/A _4767_/A _4909_/D _4772_/B VGND VGND VPWR VPWR _4646_/A sky130_fd_sc_hd__nand4_4
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__buf_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__clkbuf_2
X_3531_ hold40/A _5722_/B _5731_/B VGND VGND VPWR VPWR _3531_/X sky130_fd_sc_hd__and3_4
XANTENNA__3753__A1 input95/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR _7673_/A sky130_fd_sc_hd__buf_6
XANTENNA__3753__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput77 ser_tx VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold806 hold806/A VGND VGND VPWR VPWR _7052_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_27_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR _4131_/B sky130_fd_sc_hd__buf_4
XFILLER_6_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold828 hold828/A VGND VGND VPWR VPWR _7461_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold839 hold839/A VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6250_ _7493_/Q _6112_/C _6276_/A3 _6097_/X _7445_/Q VGND VGND VPWR VPWR _6250_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3462_ _6902_/Q _6901_/Q _4025_/A VGND VGND VPWR VPWR _3462_/X sky130_fd_sc_hd__mux2_1
X_5201_ _5203_/A _5113_/A _5055_/C _5058_/C _5158_/A VGND VGND VPWR VPWR _5202_/B
+ sky130_fd_sc_hd__a32oi_4
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3506__B _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6181_ _7530_/Q _6091_/X _6179_/X _6180_/X VGND VGND VPWR VPWR _6181_/X sky130_fd_sc_hd__a211o_1
XFILLER_143_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5132_ _4722_/Y _4727_/Y _4761_/Y _4978_/Y VGND VGND VPWR VPWR _5143_/A sky130_fd_sc_hd__o22a_1
Xhold2207 hold531/X VGND VGND VPWR VPWR _5611_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2218 _6992_/Q VGND VGND VPWR VPWR hold537/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2229 _5860_/X VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1506 _7460_/Q VGND VGND VPWR VPWR hold202/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1517 _7580_/Q VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5063_ _5203_/A _5183_/B _5183_/C _5063_/D VGND VGND VPWR VPWR _5064_/C sky130_fd_sc_hd__nand4_1
Xhold1528 hold310/X VGND VGND VPWR VPWR _5917_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3808__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1539 hold224/X VGND VGND VPWR VPWR _5935_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4014_ _4040_/D _4014_/B VGND VGND VPWR VPWR _4040_/A sky130_fd_sc_hd__nand2_4
XANTENNA__6222__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5965_ _5965_/A _5965_/B hold26/X VGND VGND VPWR VPWR _5973_/S sky130_fd_sc_hd__and3_4
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4916_ _4916_/A _4916_/B _4916_/C VGND VGND VPWR VPWR _4919_/A sky130_fd_sc_hd__nor3_1
X_5896_ _5995_/A1 _5896_/A1 _5901_/S VGND VGND VPWR VPWR _5896_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3992__A1 _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7635_ _7636_/CLK _7635_/D VGND VGND VPWR VPWR _7635_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _5059_/A _5282_/C _5453_/C VGND VGND VPWR VPWR _4847_/X sky130_fd_sc_hd__and3_2
XANTENNA__5883__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7566_ _7574_/CLK hold80/X fanout745/X VGND VGND VPWR VPWR _7566_/Q sky130_fd_sc_hd__dfrtp_4
X_4778_ _4778_/A _4778_/B _5113_/A _5410_/B VGND VGND VPWR VPWR _4778_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3744__A1 _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6517_ _7497_/Q _6466_/D _6651_/C _6452_/X _7345_/Q VGND VGND VPWR VPWR _6517_/X
+ sky130_fd_sc_hd__a32o_1
X_3729_ _7131_/Q _4455_/A _3860_/D _4479_/A _3728_/X VGND VGND VPWR VPWR _3729_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7497_ _7497_/CLK _7497_/D fanout709/X VGND VGND VPWR VPWR _7497_/Q sky130_fd_sc_hd__dfrtp_2
X_6448_ _7439_/Q _6574_/B _6574_/C _6446_/X _7519_/Q VGND VGND VPWR VPWR _6448_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6694__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6379_ _7015_/Q _6384_/A4 _6097_/C _6379_/B1 _7126_/Q VGND VGND VPWR VPWR _6379_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2730 hold743/X VGND VGND VPWR VPWR _4261_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2741 _5589_/X VGND VGND VPWR VPWR hold766/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2752 _7050_/Q VGND VGND VPWR VPWR hold807/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2763 _7491_/Q VGND VGND VPWR VPWR hold859/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6446__C _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2774 _7034_/Q VGND VGND VPWR VPWR hold853/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2785 _4459_/X VGND VGND VPWR VPWR hold978/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2796 _7135_/Q VGND VGND VPWR VPWR hold987/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1892_A _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6462__B _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3578__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__B2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3983__A1 _7343_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5793__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5094__A _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6685__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3499__B1 _3498_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output258_A _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6437__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5660__A1 hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3996__B _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4215__A2 _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5750_ _5750_/A0 _5948_/A1 _5757_/S VGND VGND VPWR VPWR _5750_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4173__A _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6091__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4888_/B _4888_/C VGND VGND VPWR VPWR _5072_/B sky130_fd_sc_hd__nor2_8
X_5681_ _5681_/A0 _5951_/A1 _5685_/S VGND VGND VPWR VPWR _5681_/X sky130_fd_sc_hd__mux2_1
X_4632_ _4767_/A _4984_/C _4628_/Y _4631_/Y VGND VGND VPWR VPWR _4632_/Y sky130_fd_sc_hd__o31ai_1
X_7420_ _7582_/CLK _7420_/D fanout717/X VGND VGND VPWR VPWR _7420_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6373__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3726__A1 _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4563_ _4563_/A _4563_/B _4563_/C _4563_/D VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__nand4_1
XANTENNA__3726__B2 _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7351_ _7563_/CLK _7351_/D fanout737/X VGND VGND VPWR VPWR _7351_/Q sky130_fd_sc_hd__dfstp_2
Xhold603 hold603/A VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5191__A3 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2540_A _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6302_ _7162_/Q _6075_/X _6099_/X _7026_/Q _6301_/X VGND VGND VPWR VPWR _6303_/D
+ sky130_fd_sc_hd__a221o_1
X_3514_ _5938_/B _3576_/B _3576_/C VGND VGND VPWR VPWR _3514_/X sky130_fd_sc_hd__and3_4
Xhold614 hold614/A VGND VGND VPWR VPWR _7354_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7282_ _7309_/CLK _7282_/D fanout704/X VGND VGND VPWR VPWR _7282_/Q sky130_fd_sc_hd__dfrtp_4
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold636 hold636/A VGND VGND VPWR VPWR _7305_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4494_ _4494_/A0 _5914_/A1 _4496_/S VGND VGND VPWR VPWR _4494_/X sky130_fd_sc_hd__mux2_1
Xhold647 hold647/A VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap355 _5658_/S VGND VGND VPWR VPWR _5657_/S sky130_fd_sc_hd__buf_2
XANTENNA__3741__A4 _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5479__A1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold658 hold658/A VGND VGND VPWR VPWR _7055_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6233_ _7340_/Q _6120_/X _6121_/X _7308_/Q _6232_/X VGND VGND VPWR VPWR _6233_/X
+ sky130_fd_sc_hd__a221o_1
X_3445_ _4772_/B VGND VGND VPWR VPWR _4814_/C sky130_fd_sc_hd__inv_16
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 hold669/A VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6140__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4151__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6121_/C _6071_/X _7289_/Q _6097_/X _7441_/Q VGND VGND VPWR VPWR _6164_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2004 _7176_/Q VGND VGND VPWR VPWR hold234/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2015 _7198_/Q VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2026 _7315_/Q VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2037 _4444_/X VGND VGND VPWR VPWR hold305/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/A _5115_/B _5115_/C VGND VGND VPWR VPWR _5115_/X sky130_fd_sc_hd__and3_2
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 hold3188/X VGND VGND VPWR VPWR hold3189/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2048 _7128_/Q VGND VGND VPWR VPWR hold471/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 hold3173/X VGND VGND VPWR VPWR _7001_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2059 hold503/X VGND VGND VPWR VPWR _5967_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6095_ _7487_/Q _6110_/A _6332_/C _6094_/X _7503_/Q VGND VGND VPWR VPWR _6095_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 hold3193/X VGND VGND VPWR VPWR hold3194/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1336 hold3232/X VGND VGND VPWR VPWR _7187_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1347 hold3191/X VGND VGND VPWR VPWR hold3192/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5046_ _5046_/A _5046_/B VGND VGND VPWR VPWR _5047_/B sky130_fd_sc_hd__nor2_1
Xhold1358 _4313_/B VGND VGND VPWR VPWR hold3025/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1369 _4278_/B VGND VGND VPWR VPWR hold3047/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5878__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6997_ _7633_/CLK _6997_/D VGND VGND VPWR VPWR _6997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5403__B2 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_A _7591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5948_ _5948_/A0 _5948_/A1 _5955_/S VGND VGND VPWR VPWR _5948_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5879_ _5879_/A0 _5978_/A0 _5883_/S VGND VGND VPWR VPWR _5879_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1473_A _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7618_ _7621_/CLK _7618_/D fanout705/X VGND VGND VPWR VPWR _7618_/Q sky130_fd_sc_hd__dfrtp_1
X_7549_ _7556_/CLK _7549_/D fanout732/X VGND VGND VPWR VPWR _7549_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold1640_A _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6667__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_150_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_823 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input156_A wb_dat_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3250 _7495_/Q VGND VGND VPWR VPWR hold3250/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6457__B _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3261 _7535_/Q VGND VGND VPWR VPWR hold3261/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3272 _7217_/Q VGND VGND VPWR VPWR _3797_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3283 _7639_/Q VGND VGND VPWR VPWR _6807_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3294 _6676_/X VGND VGND VPWR VPWR _7623_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2560 _4342_/X VGND VGND VPWR VPWR hold922/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold3119_A _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2571 _6971_/Q VGND VGND VPWR VPWR hold673/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2582 _7373_/Q VGND VGND VPWR VPWR hold823/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2593 _5864_/X VGND VGND VPWR VPWR hold828/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5788__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5642__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1870 _4489_/X VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input17_A mask_rev_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1881 hold134/X VGND VGND VPWR VPWR _5901_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1892 _7330_/Q VGND VGND VPWR VPWR hold336/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4705__B _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6198__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__B2 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3708__A1 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__B2 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5173__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4381__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6658__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4133__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6673__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5881__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6086__C _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3503__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5698__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5633__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6920_ _7255_/CLK _6920_/D fanout688/X VGND VGND VPWR VPWR _6920_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6851_ _6869_/A _6872_/B VGND VGND VPWR VPWR _6851_/X sky130_fd_sc_hd__and2_1
XANTENNA__4615__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5802_ _5955_/A1 _5802_/A1 _5802_/S VGND VGND VPWR VPWR _5802_/X sky130_fd_sc_hd__mux2_1
X_3994_ input34/X _3486_/X _3990_/X _3992_/X _3993_/X VGND VGND VPWR VPWR _3995_/D
+ sky130_fd_sc_hd__a2111oi_4
X_6782_ _6792_/S _3996_/B _6781_/Y VGND VGND VPWR VPWR _7629_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__4334__C _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5733_ _5733_/A0 _5949_/A1 _5739_/S VGND VGND VPWR VPWR _5733_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2755_A _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5664_ _5664_/A0 _5952_/A1 _5667_/S VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7403_ _7435_/CLK _7403_/D fanout736/X VGND VGND VPWR VPWR _7403_/Q sky130_fd_sc_hd__dfrtp_4
X_4615_ _4615_/A _4645_/D VGND VGND VPWR VPWR _4615_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_54_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7306_/CLK sky130_fd_sc_hd__clkbuf_16
X_5595_ _5595_/A0 _5736_/A1 _5595_/S VGND VGND VPWR VPWR _5595_/X sky130_fd_sc_hd__mux2_1
Xhold400 hold400/A VGND VGND VPWR VPWR _7002_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7334_ _7334_/CLK _7334_/D fanout711/X VGND VGND VPWR VPWR _7334_/Q sky130_fd_sc_hd__dfrtp_4
Xhold411 hold411/A VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4546_ _5582_/A0 _4546_/A1 _4550_/S VGND VGND VPWR VPWR _4546_/X sky130_fd_sc_hd__mux2_1
Xhold422 hold422/A VGND VGND VPWR VPWR _7086_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold433 hold433/A VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold444 hold444/A VGND VGND VPWR VPWR _7322_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold466 hold466/A VGND VGND VPWR VPWR _7138_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7265_ _7266_/CLK _7265_/D _6873_/A VGND VGND VPWR VPWR _7265_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6113__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4477_ _4477_/A0 _5585_/A0 _4478_/S VGND VGND VPWR VPWR _4477_/X sky130_fd_sc_hd__mux2_1
Xhold477 hold477/A VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold488 hold488/A VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3428_ _7418_/Q VGND VGND VPWR VPWR _3428_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_69_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7360_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold499 hold499/A VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6216_ _7492_/Q _6075_/A _6276_/A3 _6097_/X _7444_/Q VGND VGND VPWR VPWR _6216_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_131_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7196_ _7212_/CLK _7196_/D fanout721/X VGND VGND VPWR VPWR _7196_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6664__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6147_ _6146_/X _6145_/Y _6069_/X _6169_/A2 VGND VGND VPWR VPWR _7603_/D sky130_fd_sc_hd__o2bb2a_1
XANTENNA_input9_A mask_rev_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5612__D _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1100 hold3031/X VGND VGND VPWR VPWR hold1100/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout573_A _5635_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 hold2987/X VGND VGND VPWR VPWR hold1111/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4509__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1122 hold3124/X VGND VGND VPWR VPWR _6874_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1133 hold3127/X VGND VGND VPWR VPWR hold3128/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1144 hold3142/X VGND VGND VPWR VPWR _7137_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6078_ _6099_/D _6081_/C VGND VGND VPWR VPWR _6078_/X sky130_fd_sc_hd__and2b_1
XTAP_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 hold1155/A VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
XANTENNA__5624__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1166 hold2910/X VGND VGND VPWR VPWR hold2911/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1177 hold2863/X VGND VGND VPWR VPWR hold2864/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5029_ _5029_/A _5034_/B _5030_/C VGND VGND VPWR VPWR _5031_/A sky130_fd_sc_hd__and3_1
Xhold1188 _5752_/X VGND VGND VPWR VPWR _7361_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4806__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 hold2903/X VGND VGND VPWR VPWR hold2904/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3938__A1 _7243_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6352__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4899__C1 wire649/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4363__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6468__A _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6104__A2 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5803__C _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6655__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5091__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3080 hold3080/A VGND VGND VPWR VPWR _5921_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3091 hold3091/A VGND VGND VPWR VPWR hold3091/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2390 hold733/X VGND VGND VPWR VPWR _5725_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5615__A1 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3626__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6591__A2 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4170__B _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5146__A3 _4977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4400_ _5596_/A _4527_/A _5596_/B _5619_/C VGND VGND VPWR VPWR _4405_/S sky130_fd_sc_hd__and4_4
XANTENNA__4354__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5380_ _5255_/X _5509_/A3 _5480_/A1 _4737_/Y _5563_/A1 VGND VGND VPWR VPWR _5380_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_126_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4331_ _4331_/A0 _4548_/A0 _4333_/S VGND VGND VPWR VPWR _4331_/X sky130_fd_sc_hd__mux2_1
X_7050_ _7471_/CLK _7050_/D fanout729/X VGND VGND VPWR VPWR _7050_/Q sky130_fd_sc_hd__dfrtp_4
X_4262_ _4262_/A0 _5815_/A1 _4264_/S VGND VGND VPWR VPWR _4262_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6097__B _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6001_ _6932_/Q _6929_/Q _4100_/X VGND VGND VPWR VPWR _6001_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_140_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4193_ _4193_/A0 _5645_/A0 _4202_/S VGND VGND VPWR VPWR _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5606__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3530__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5082__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6903_ _4150_/A1 _6903_/D _6853_/X VGND VGND VPWR VPWR _6903_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6834_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6834_/X sky130_fd_sc_hd__and2_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6765_ _6992_/Q _6420_/B _6460_/X _7116_/Q VGND VGND VPWR VPWR _6765_/X sky130_fd_sc_hd__a22o_1
X_3977_ _6927_/Q hold90/A _4265_/B _3682_/X _7224_/Q VGND VGND VPWR VPWR _3977_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__6582__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5716_ _5995_/A1 _5716_/A1 _5721_/S VGND VGND VPWR VPWR _5716_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6696_ _6989_/Q _6420_/B _6422_/X _6963_/Q _6695_/X VGND VGND VPWR VPWR _6697_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _5647_/A0 _5647_/A1 _5649_/S VGND VGND VPWR VPWR _5647_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7672__A _7672_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5578_ _4707_/Y _4722_/Y _5089_/Y _5254_/X _5474_/C VGND VGND VPWR VPWR _5578_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA_clkbuf_leaf_75_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 hold230/A VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3699__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7317_ _7478_/CLK _7317_/D fanout714/X VGND VGND VPWR VPWR _7317_/Q sky130_fd_sc_hd__dfrtp_4
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold252 hold252/A VGND VGND VPWR VPWR _6991_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4529_ _4529_/A0 _4547_/A0 _4532_/S VGND VGND VPWR VPWR _4529_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold263 hold263/A VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__B2 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold285 _5754_/X VGND VGND VPWR VPWR _7363_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4300__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7248_ _7250_/CLK _7248_/D _6873_/A VGND VGND VPWR VPWR _7248_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5623__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout710 fanout711/X VGND VGND VPWR VPWR fanout710/X sky130_fd_sc_hd__buf_8
Xfanout721 fanout724/X VGND VGND VPWR VPWR fanout721/X sky130_fd_sc_hd__buf_8
XANTENNA__5845__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout732 fanout736/X VGND VGND VPWR VPWR fanout732/X sky130_fd_sc_hd__clkbuf_8
Xfanout743 fanout749/X VGND VGND VPWR VPWR fanout743/X sky130_fd_sc_hd__buf_8
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout754 _4860_/A VGND VGND VPWR VPWR _4767_/A sky130_fd_sc_hd__buf_8
X_7179_ _7179_/CLK _7179_/D fanout698/X VGND VGND VPWR VPWR _7179_/Q sky130_fd_sc_hd__dfstp_2
Xfanout765 _5407_/A1 VGND VGND VPWR VPWR _4887_/B sky130_fd_sc_hd__buf_12
XANTENNA__5920__A _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout776 _4887_/D VGND VGND VPWR VPWR _4879_/D sky130_fd_sc_hd__buf_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3440__A _7322_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6270__A1 _7414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input119_A wb_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5781__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input84_A spimemio_flash_csb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4336__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5836__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4639__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5830__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6645__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3614__A3 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3900_ _7067_/Q _3649_/X _3675_/X _7188_/Q VGND VGND VPWR VPWR _3900_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4880_ _5282_/A _5199_/C VGND VGND VPWR VPWR _4880_/Y sky130_fd_sc_hd__nand2_4
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3831_ _7409_/Q _3493_/X _3657_/X _6959_/Q _3830_/X VGND VGND VPWR VPWR _3837_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6564__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6550_ _7451_/Q _6467_/A _6771_/A3 _6446_/X _7523_/Q VGND VGND VPWR VPWR _6550_/X
+ sky130_fd_sc_hd__a32o_1
X_3762_ _7474_/Q _3494_/X _5704_/A _7322_/Q _3737_/X VGND VGND VPWR VPWR _3762_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_158_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ _5501_/A _5501_/B VGND VGND VPWR VPWR _5504_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3693_ _7347_/Q _3590_/C _4352_/A _3659_/X _7010_/Q VGND VGND VPWR VPWR _3693_/X
+ sky130_fd_sc_hd__a32o_1
X_6481_ _7456_/Q _4101_/X _6574_/C _6425_/X _7336_/Q VGND VGND VPWR VPWR _6481_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6316__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5432_ _4667_/B _4821_/Y _5174_/Y _5012_/Y VGND VGND VPWR VPWR _5433_/C sky130_fd_sc_hd__a31o_1
XFILLER_173_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput302 _3619_/X VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput313 hold1088/X VGND VGND VPWR VPWR hold1089/A sky130_fd_sc_hd__buf_6
Xoutput324 hold1183/X VGND VGND VPWR VPWR hold1184/A sky130_fd_sc_hd__buf_6
X_5363_ _5347_/X _5363_/B _5510_/A VGND VGND VPWR VPWR _5367_/C sky130_fd_sc_hd__nand3b_1
Xoutput335 hold1154/X VGND VGND VPWR VPWR hold1155/A sky130_fd_sc_hd__buf_6
XANTENNA__3525__A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7102_ _7111_/CLK _7102_/D fanout751/X VGND VGND VPWR VPWR _7102_/Q sky130_fd_sc_hd__dfrtp_4
X_4314_ _4321_/S _3856_/B _4313_/Y VGND VGND VPWR VPWR _6995_/D sky130_fd_sc_hd__o21ai_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5294_ _5294_/A _5294_/B _5294_/C VGND VGND VPWR VPWR _5294_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5827__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4245_ _4245_/A0 _4244_/X _4249_/S VGND VGND VPWR VPWR _4245_/X sky130_fd_sc_hd__mux2_1
X_7033_ _7035_/CLK _7033_/D fanout723/X VGND VGND VPWR VPWR _7033_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_141_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5740__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4176_ _7263_/Q _4176_/B VGND VGND VPWR VPWR _4176_/X sky130_fd_sc_hd__and2_2
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout369_A hold31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6817_ _4427_/D _6817_/A2 _6817_/B1 _4427_/C VGND VGND VPWR VPWR _6817_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6555__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5358__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6891__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5763__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6748_ _7024_/Q _6452_/X _6747_/X _6746_/X _6745_/X VGND VGND VPWR VPWR _6749_/D
+ sky130_fd_sc_hd__a2111o_1
XFILLER_137_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold114_A _7227_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7423__SET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6679_ _7148_/Q _6408_/A _6451_/X _6875_/Q _6678_/X VGND VGND VPWR VPWR _6679_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4318__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7411__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3435__A _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1720_A _7528_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5818__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3829__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout540 hold1494/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__clkbuf_2
Xfanout551 _5952_/A1 VGND VGND VPWR VPWR _5736_/A1 sky130_fd_sc_hd__buf_8
XANTENNA__6491__A1 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout562 _5996_/A1 VGND VGND VPWR VPWR _5585_/A0 sky130_fd_sc_hd__buf_6
Xfanout573 _5635_/A0 VGND VGND VPWR VPWR _5788_/A1 sky130_fd_sc_hd__buf_6
Xmgmt_gpio_14_buff_inst _4162_/X VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_8
Xfanout584 _5894_/A0 VGND VGND VPWR VPWR _5948_/A1 sky130_fd_sc_hd__buf_4
Xfanout595 hold26/X VGND VGND VPWR VPWR _5893_/B sky130_fd_sc_hd__buf_12
XFILLER_76_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5796__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6546__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3780__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5809__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4030_ _6904_/Q _4025_/B _4025_/A VGND VGND VPWR VPWR _4030_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6482__A1 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5285__A2 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3835__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold2201_A _7025_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5981_ _5990_/A1 _5981_/A1 _5982_/S VGND VGND VPWR VPWR _5981_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6785__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3599__A2 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4932_ _4947_/C _4997_/B _4933_/A _5260_/D VGND VGND VPWR VPWR _4932_/X sky130_fd_sc_hd__and4_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7651_ _7651_/A VGND VGND VPWR VPWR _7651_/X sky130_fd_sc_hd__clkbuf_2
X_4863_ _4805_/B _4668_/C _4660_/Y VGND VGND VPWR VPWR _5053_/C sky130_fd_sc_hd__o21a_4
XANTENNA__4623__B _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6537__A2 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ _7349_/Q _6452_/X _6463_/X _7429_/Q VGND VGND VPWR VPWR _6602_/X sky130_fd_sc_hd__a22o_1
XANTENNA_14 _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _7297_/Q _3848_/A2 _5731_/B input26/X _3503_/X VGND VGND VPWR VPWR _3814_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_25 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7582_ _7582_/CLK _7582_/D fanout718/X VGND VGND VPWR VPWR _7582_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_36 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _4794_/A _4803_/A _5410_/B VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__and3_1
XANTENNA_47 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_58 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ _7354_/Q _6561_/A2 _6428_/X _6451_/X _7482_/Q VGND VGND VPWR VPWR _6533_/X
+ sky130_fd_sc_hd__a32o_1
X_3745_ _7370_/Q _5758_/A _4370_/A _7044_/Q VGND VGND VPWR VPWR _3745_/X sky130_fd_sc_hd__a22o_1
XFILLER_192_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3771__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6464_ _7375_/Q _6408_/B _6463_/X _7423_/Q VGND VGND VPWR VPWR _6464_/X sky130_fd_sc_hd__a22o_1
X_3676_ _7060_/Q _4539_/C _4364_/B _4322_/A _7005_/Q VGND VGND VPWR VPWR _3676_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_173_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5415_ _4706_/Y _4796_/Y _4802_/Y _4759_/Y _5414_/Y VGND VGND VPWR VPWR _5535_/B
+ sky130_fd_sc_hd__o221a_1
X_6395_ _7050_/Q _6317_/B _6317_/C _6072_/X _7156_/Q VGND VGND VPWR VPWR _6395_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3523__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5346_ _5089_/D _4939_/C _4942_/A _4948_/C VGND VGND VPWR VPWR _5346_/X sky130_fd_sc_hd__o211a_4
Xoutput176 _3435_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 _3425_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
Xoutput198 _3415_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
Xhold2901 hold2901/A VGND VGND VPWR VPWR _4385_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_153_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2912 _7442_/Q VGND VGND VPWR VPWR hold2912/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2923 _6964_/Q VGND VGND VPWR VPWR hold2923/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5277_ _5222_/A _5061_/B _5399_/C _5107_/C VGND VGND VPWR VPWR _5277_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout486_A _6084_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2934 _7490_/Q VGND VGND VPWR VPWR hold2934/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2945 _7013_/Q VGND VGND VPWR VPWR hold2945/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5276__A2 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7016_ _7211_/CLK _7016_/D fanout699/X VGND VGND VPWR VPWR _7016_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2956 hold2956/A VGND VGND VPWR VPWR _4548_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4228_ _4228_/A0 _4227_/X _4232_/S VGND VGND VPWR VPWR _4228_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2967 hold2967/A VGND VGND VPWR VPWR hold2967/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2978 _6973_/Q VGND VGND VPWR VPWR _4280_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2989 hold2989/A VGND VGND VPWR VPWR hold2989/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4159_ input1/X input2/X VGND VGND VPWR VPWR _4159_/Y sky130_fd_sc_hd__nand2_4
XFILLER_83_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6225__A1 _7292_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4814__A _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6528__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4533__B _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1768_A _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5197__D1 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3762__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A mgmt_gpio_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout370 _4864_/X VGND VGND VPWR VPWR _5180_/A sky130_fd_sc_hd__buf_6
Xfanout381 _6839_/B VGND VGND VPWR VPWR _6872_/B sky130_fd_sc_hd__buf_4
XFILLER_143_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout392 _3562_/C VGND VGND VPWR VPWR _5731_/B sky130_fd_sc_hd__buf_6
XFILLER_120_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4427__C _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6216__A1 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6216__B2 _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6767__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__A0 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output203_A wire378/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6519__A2 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_2
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__buf_4
X_3530_ _5612_/A _3682_/A hold32/X VGND VGND VPWR VPWR _5857_/A sky130_fd_sc_hd__and3_4
XFILLER_116_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3753__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__buf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR _4168_/D sky130_fd_sc_hd__buf_12
Xhold807 hold807/A VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap515 wire516/X VGND VGND VPWR VPWR _5399_/D sky130_fd_sc_hd__clkbuf_2
Xinput78 spi_csb VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_4
XFILLER_171_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold818 hold818/A VGND VGND VPWR VPWR _6968_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap537 _4426_/Y VGND VGND VPWR VPWR wire536/A sky130_fd_sc_hd__clkbuf_4
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3461_ _3460_/X hold103/X _4181_/S VGND VGND VPWR VPWR _3505_/C sky130_fd_sc_hd__mux2_1
XFILLER_116_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6089__C _6089_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5200_ _5200_/A _5200_/B _5200_/C VGND VGND VPWR VPWR _5202_/A sky130_fd_sc_hd__and3_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3506__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6180_ _7466_/Q _6121_/A _6116_/A _6267_/B1 _7522_/Q VGND VGND VPWR VPWR _6180_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2208 _5611_/X VGND VGND VPWR VPWR hold532/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5131_ _5480_/A1 _5561_/A1 _4716_/Y _5028_/C VGND VGND VPWR VPWR _5145_/A sky130_fd_sc_hd__o31a_1
Xhold2219 hold537/X VGND VGND VPWR VPWR _4308_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1507 hold202/X VGND VGND VPWR VPWR _5863_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5062_ _5495_/C1 _4654_/Y _4880_/Y _4846_/Y _4744_/Y VGND VGND VPWR VPWR _5064_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_97_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1518 hold180/X VGND VGND VPWR VPWR _5998_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1529 _5917_/X VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4013_ _6892_/Q _6891_/Q _3401_/Y _4062_/A _4011_/X VGND VGND VPWR VPWR _4014_/B
+ sky130_fd_sc_hd__o311ai_4
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6833__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6758__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5964_ _5964_/A0 hold20/X _5964_/S VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__mux2_1
X_4915_ _5213_/B _5260_/D _4915_/C VGND VGND VPWR VPWR _4916_/B sky130_fd_sc_hd__and3_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5895_ _5994_/A1 _5895_/A1 _5901_/S VGND VGND VPWR VPWR _5895_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5718__A0 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7634_ _7636_/CLK _7634_/D VGND VGND VPWR VPWR _7634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ _5059_/A _5282_/C VGND VGND VPWR VPWR _4846_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__3992__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6391__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7565_ _7565_/CLK hold84/X fanout746/X VGND VGND VPWR VPWR _7565_/Q sky130_fd_sc_hd__dfrtp_4
X_4777_ _4733_/A _4733_/B _4641_/B _4768_/Y VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__a211o_1
XFILLER_147_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout401_A _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6516_ _7545_/Q _6419_/A _6512_/X _6515_/X VGND VGND VPWR VPWR _6516_/X sky130_fd_sc_hd__a211o_4
X_3728_ _7141_/Q _4479_/A _4364_/B _5974_/A _7563_/Q VGND VGND VPWR VPWR _3728_/X
+ sky130_fd_sc_hd__a32o_1
X_7496_ _7537_/CLK _7496_/D fanout707/X VGND VGND VPWR VPWR _7496_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_113_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6447_ _6455_/B _6447_/B _6447_/C VGND VGND VPWR VPWR _6447_/X sky130_fd_sc_hd__and3_4
X_3659_ _4328_/A _4388_/B _4346_/C VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__and3_4
XFILLER_162_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6694__B2 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6378_ _6377_/X _6376_/Y _6069_/X _6400_/A2 VGND VGND VPWR VPWR _7613_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_115_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout770_A _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5329_ _5011_/B _5183_/C _5049_/C _5038_/B _5339_/A VGND VGND VPWR VPWR _5329_/X
+ sky130_fd_sc_hd__o311a_2
Xhold2720 hold755/X VGND VGND VPWR VPWR _4550_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5249__A2 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2731 _7264_/Q VGND VGND VPWR VPWR hold745/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2742 _7381_/Q VGND VGND VPWR VPWR hold937/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2753 hold807/X VGND VGND VPWR VPWR _4381_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2764 hold859/X VGND VGND VPWR VPWR _5898_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2775 hold853/X VGND VGND VPWR VPWR _4362_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2786 _7523_/Q VGND VGND VPWR VPWR hold875/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2797 hold987/X VGND VGND VPWR VPWR _4477_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3680__A1 _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input101_A wb_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5709__A0 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3983__A2 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6382__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3266_A _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6134__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6685__A1 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4160__A2 input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3623__A _3623_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6437__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5260__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4215__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4700_ _4887_/B _5399_/B VGND VGND VPWR VPWR _4700_/Y sky130_fd_sc_hd__nand2b_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4604__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A0 _5995_/A1 _5685_/S VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4631_ _4570_/Y _5494_/B2 _4767_/A VGND VGND VPWR VPWR _4631_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6373__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7350_ _7365_/CLK _7350_/D fanout713/X VGND VGND VPWR VPWR _7350_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3726__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4562_ _4562_/A _4562_/B _4562_/C _4562_/D VGND VGND VPWR VPWR _4562_/Y sky130_fd_sc_hd__nand4_4
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold604 hold604/A VGND VGND VPWR VPWR _7310_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6301_ _7046_/Q _6332_/B _6317_/C _6072_/X _7152_/Q VGND VGND VPWR VPWR _6301_/X
+ sky130_fd_sc_hd__a32o_1
X_3513_ _7574_/Q _3872_/A2 _5965_/A _5686_/A _7310_/Q VGND VGND VPWR VPWR _3513_/X
+ sky130_fd_sc_hd__a32o_1
Xhold615 hold615/A VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7281_ _7329_/CLK _7281_/D fanout704/X VGND VGND VPWR VPWR _7281_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6125__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold626 hold626/A VGND VGND VPWR VPWR _7483_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4493_ _4493_/A0 _4553_/A0 _4496_/S VGND VGND VPWR VPWR _4493_/X sky130_fd_sc_hd__mux2_1
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold648 hold648/A VGND VGND VPWR VPWR _7531_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5479__A2 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold659 hold659/A VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6232_ _7436_/Q _6110_/X _6116_/X _7316_/Q VGND VGND VPWR VPWR _6232_/X sky130_fd_sc_hd__a22o_1
XFILLER_104_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3444_ _6332_/B VGND VGND VPWR VPWR _3444_/Y sky130_fd_sc_hd__inv_6
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _7449_/Q _6081_/X _6089_/X _7505_/Q _6162_/X VGND VGND VPWR VPWR _6163_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2005 hold234/X VGND VGND VPWR VPWR _4526_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2016 hold445/X VGND VGND VPWR VPWR _4553_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2027 hold397/X VGND VGND VPWR VPWR _5700_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2038 _7576_/Q VGND VGND VPWR VPWR hold499/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5114_ _5118_/A _5399_/C _5282_/C _5113_/X VGND VGND VPWR VPWR _5559_/A sky130_fd_sc_hd__a31o_1
Xhold1304 hold3190/X VGND VGND VPWR VPWR _7222_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6112_/C _6119_/A _6119_/B _6097_/B VGND VGND VPWR VPWR _6094_/X sky130_fd_sc_hd__and4_4
XFILLER_97_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2049 hold471/X VGND VGND VPWR VPWR _4469_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 hold3183/X VGND VGND VPWR VPWR hold3184/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 hold3195/X VGND VGND VPWR VPWR _7016_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1337 hold3201/X VGND VGND VPWR VPWR hold3202/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1348 _4510_/X VGND VGND VPWR VPWR _7162_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5045_ _5339_/D _5183_/C _5183_/B VGND VGND VPWR VPWR _5046_/B sky130_fd_sc_hd__nand3_1
Xhold1359 _4280_/A1 VGND VGND VPWR VPWR hold2979/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4364__A _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6996_ _6999_/CLK _6996_/D VGND VGND VPWR VPWR _6996_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout449_A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5947_ _5947_/A _5947_/B _5947_/C VGND VGND VPWR VPWR _5955_/S sky130_fd_sc_hd__and3_4
XFILLER_179_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5894__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6796__B1_N _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3965__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5878_ _5878_/A0 _5950_/A1 _5883_/S VGND VGND VPWR VPWR _5878_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout616_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7617_ _7621_/CLK _7617_/D fanout705/X VGND VGND VPWR VPWR _7617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6364__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4829_ _5089_/D _5399_/C _5282_/C VGND VGND VPWR VPWR _4830_/B sky130_fd_sc_hd__and3_1
XFILLER_166_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3717__A2 _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7548_ _7548_/CLK _7548_/D fanout734/X VGND VGND VPWR VPWR _7548_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7479_ _7562_/CLK _7479_/D fanout739/X VGND VGND VPWR VPWR _7479_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6667__A1 _7197_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4539__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3240 _7359_/Q VGND VGND VPWR VPWR hold3240/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3251 hold3251/A VGND VGND VPWR VPWR _5903_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3262 hold3262/A VGND VGND VPWR VPWR _5948_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3273 _3797_/X VGND VGND VPWR VPWR _7217_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input149_A wb_dat_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3284 _7641_/Q VGND VGND VPWR VPWR _6813_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3295 _7644_/Q VGND VGND VPWR VPWR _6822_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2550 _7449_/Q VGND VGND VPWR VPWR hold839/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2561 _7437_/Q VGND VGND VPWR VPWR hold837/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2572 hold673/X VGND VGND VPWR VPWR _4276_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2583 hold823/X VGND VGND VPWR VPWR _5765_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2594 _7129_/Q VGND VGND VPWR VPWR hold913/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1860 hold363/X VGND VGND VPWR VPWR _4476_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1871 _6991_/Q VGND VGND VPWR VPWR hold1871/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1882 _5901_/X VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1893 hold336/X VGND VGND VPWR VPWR _5717_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4721__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output270_A _6913_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6107__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4118__C1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6658__A1 _7026_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6658__B2 _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4669__B1 _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5330__B2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4168__B _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3892__A1 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3644__A1 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6850_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6850_/X sky130_fd_sc_hd__and2_1
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5801_ _5999_/A1 _5801_/A1 _5802_/S VGND VGND VPWR VPWR _5801_/X sky130_fd_sc_hd__mux2_1
X_6781_ _6792_/S _6781_/B VGND VGND VPWR VPWR _6781_/Y sky130_fd_sc_hd__nand2_1
X_3993_ _6988_/Q _5731_/B _5623_/B _5704_/A _7319_/Q VGND VGND VPWR VPWR _3993_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_16_791 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4334__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5732_ _5732_/A0 _5732_/A1 _5739_/S VGND VGND VPWR VPWR _5732_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3947__A2 _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5149__A1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5663_ _5663_/A0 _5951_/A1 _5667_/S VGND VGND VPWR VPWR _5663_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6346__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7402_ _7576_/CLK _7402_/D fanout731/X VGND VGND VPWR VPWR _7402_/Q sky130_fd_sc_hd__dfrtp_4
X_4614_ _4657_/D _4657_/C _4909_/C _4909_/A VGND VGND VPWR VPWR _4870_/A sky130_fd_sc_hd__a22oi_4
X_5594_ hold114/X _5625_/A1 _5595_/S VGND VGND VPWR VPWR _5594_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7333_ _7334_/CLK _7333_/D fanout710/X VGND VGND VPWR VPWR _7333_/Q sky130_fd_sc_hd__dfrtp_4
X_4545_ _4545_/A _4551_/D VGND VGND VPWR VPWR _4550_/S sky130_fd_sc_hd__nand2_4
XFILLER_128_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold412 hold412/A VGND VGND VPWR VPWR _7385_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold434 hold434/A VGND VGND VPWR VPWR _7448_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold445 hold445/A VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7264_ _7264_/CLK _7264_/D fanout689/X VGND VGND VPWR VPWR _7264_/Q sky130_fd_sc_hd__dfrtp_1
X_4476_ _4476_/A0 _5788_/A1 _4478_/S VGND VGND VPWR VPWR _4476_/X sky130_fd_sc_hd__mux2_1
Xhold456 _5788_/X VGND VGND VPWR VPWR _7393_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold467 hold467/A VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6113__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold478 hold478/A VGND VGND VPWR VPWR _6940_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6215_ _6214_/X _6237_/A2 _6573_/S VGND VGND VPWR VPWR _6215_/X sky130_fd_sc_hd__mux2_1
Xhold489 hold489/A VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3427_ _7426_/Q VGND VGND VPWR VPWR _3427_/Y sky130_fd_sc_hd__clkinv_2
X_7195_ _7213_/CLK _7195_/D fanout701/X VGND VGND VPWR VPWR _7195_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5321__B2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout399_A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ _6649_/S _7602_/Q _4116_/X _6067_/X VGND VGND VPWR VPWR _6146_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4078__B _4078_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 hold1101/A VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1112 hold1112/A VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
XANTENNA__4509__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1123 hold3064/X VGND VGND VPWR VPWR hold1123/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6077_ _7343_/Q _6070_/X _6072_/X _7415_/Q _6076_/X VGND VGND VPWR VPWR _6102_/A
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6574__A _7444_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1134 hold3129/X VGND VGND VPWR VPWR _7026_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout566_A _5726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1145 hold3146/X VGND VGND VPWR VPWR hold3147/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 hold3018/X VGND VGND VPWR VPWR hold1156/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1167 _5630_/X VGND VGND VPWR VPWR _5631_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1178 hold2865/X VGND VGND VPWR VPWR _7237_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5028_ _5028_/A _5028_/B _5028_/C VGND VGND VPWR VPWR _5031_/C sky130_fd_sc_hd__nand3_1
XANTENNA__3635__A1 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 hold2882/X VGND VGND VPWR VPWR hold2883/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3635__B2 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_71_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6585__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6979_ _7636_/CLK _6979_/D VGND VGND VPWR VPWR _6979_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3938__A2 _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6337__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6085__A_N _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6468__B _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5312__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold990 hold990/A VGND VGND VPWR VPWR _7276_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3070 hold3070/A VGND VGND VPWR VPWR _4389_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3081 _5921_/X VGND VGND VPWR VPWR hold3081/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5799__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3092 _7487_/Q VGND VGND VPWR VPWR hold3092/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2380 hold821/X VGND VGND VPWR VPWR _5657_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6812__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2391 _5725_/X VGND VGND VPWR VPWR hold734/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4969__A4 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1690 hold112/X VGND VGND VPWR VPWR _5874_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_32_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5379__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6576__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6343__A3 _6086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4330_ _4330_/A0 hold198/X _4333_/S VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__mux2_1
X_4261_ _4261_/A0 _5645_/A0 _4264_/S VGND VGND VPWR VPWR _4261_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6500__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6000_ _6000_/A0 _6000_/A1 _6000_/S VGND VGND VPWR VPWR _6000_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2329_A _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4192_ _4192_/A0 _5732_/A1 _4202_/S VGND VGND VPWR VPWR _4192_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6803__A1 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3530__B _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6902_ _4150_/A1 _6902_/D _6852_/X VGND VGND VPWR VPWR _6902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6833_ _6839_/A _6839_/B VGND VGND VPWR VPWR _6833_/X sky130_fd_sc_hd__and2_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6567__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6764_ _6878_/Q _6451_/X _6759_/X _6761_/X _6763_/X VGND VGND VPWR VPWR _6774_/B
+ sky130_fd_sc_hd__a2111oi_4
X_3976_ _7583_/Q _5659_/B _4364_/B _3973_/X _3975_/X VGND VGND VPWR VPWR _3988_/B
+ sky130_fd_sc_hd__a311o_1
X_5715_ _5949_/A1 _5715_/A1 _5721_/S VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5790__A1 _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6695_ _7138_/Q _6419_/C _6446_/X _7188_/Q VGND VGND VPWR VPWR _6695_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ _5986_/A1 _5646_/A1 _5649_/S VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5577_ _5533_/Y _5569_/X _5576_/X VGND VGND VPWR VPWR _5577_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_191_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7316_ _7478_/CLK _7316_/D fanout713/X VGND VGND VPWR VPWR _7316_/Q sky130_fd_sc_hd__dfrtp_4
Xhold231 hold231/A VGND VGND VPWR VPWR _7521_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4528_ _4528_/A0 _5582_/A0 _4532_/S VGND VGND VPWR VPWR _4528_/X sky130_fd_sc_hd__mux2_1
Xhold242 hold242/A VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold253 hold253/A VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold264 hold264/A VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6098__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold275 hold275/A VGND VGND VPWR VPWR _7538_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7247_ _7334_/CLK _7247_/D fanout710/X VGND VGND VPWR VPWR _7247_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout683_A _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4459_ _4459_/A0 _4555_/A0 _4460_/S VGND VGND VPWR VPWR _4459_/X sky130_fd_sc_hd__mux2_1
Xhold286 hold286/A VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout700 fanout702/X VGND VGND VPWR VPWR fanout700/X sky130_fd_sc_hd__buf_8
Xhold297 hold297/A VGND VGND VPWR VPWR _7160_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout711 fanout720/X VGND VGND VPWR VPWR fanout711/X sky130_fd_sc_hd__buf_8
Xfanout722 fanout724/X VGND VGND VPWR VPWR fanout722/X sky130_fd_sc_hd__buf_8
XFILLER_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout733 fanout736/X VGND VGND VPWR VPWR fanout733/X sky130_fd_sc_hd__buf_8
Xfanout744 fanout749/X VGND VGND VPWR VPWR fanout744/X sky130_fd_sc_hd__buf_4
X_7178_ _7181_/CLK _7178_/D fanout721/X VGND VGND VPWR VPWR _7178_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout755 input128/X VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__clkbuf_16
Xfanout766 _5407_/A1 VGND VGND VPWR VPWR _4748_/A sky130_fd_sc_hd__buf_4
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _7448_/Q _6144_/A _6116_/A _6379_/B1 _7520_/Q VGND VGND VPWR VPWR _6129_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_100_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A1 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1965_A _7028_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4271__B _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6325__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input77_A ser_tx VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6730__B1 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3847__A1 _7246_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5830__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6645__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_csclk _7399_/CLK VGND VGND VPWR VPWR _7478_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6261__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4272__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6549__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3830_ _6964_/Q _5632_/B _5659_/B _3829_/X VGND VGND VPWR VPWR _3830_/X sky130_fd_sc_hd__a31o_1
XFILLER_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_68_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7537_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ input6/X _5695_/A _5612_/B _3542_/X _6922_/Q VGND VGND VPWR VPWR _3761_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5772__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2181_A _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5500_ _5053_/C _5329_/X _5426_/X _5203_/B _5171_/X VGND VGND VPWR VPWR _5501_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3783__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6480_ _7432_/Q _6747_/B _6747_/C _6421_/X _7320_/Q VGND VGND VPWR VPWR _6480_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4980__C1 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3692_ _7055_/Q _3931_/B _5619_/B _3649_/X _7070_/Q VGND VGND VPWR VPWR _3692_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ _5342_/B _4956_/Y _5180_/A _4876_/Y VGND VGND VPWR VPWR _5499_/A sky130_fd_sc_hd__o211a_1
XFILLER_146_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6721__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput303 _3578_/X VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
Xoutput314 hold1076/X VGND VGND VPWR VPWR hold1077/A sky130_fd_sc_hd__buf_6
XFILLER_114_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5362_ _4954_/C _4933_/A _5346_/X _5233_/X VGND VGND VPWR VPWR _5510_/A sky130_fd_sc_hd__a31oi_2
Xoutput325 hold1100/X VGND VGND VPWR VPWR hold1101/A sky130_fd_sc_hd__buf_6
Xoutput336 hold1147/X VGND VGND VPWR VPWR hold1148/A sky130_fd_sc_hd__buf_6
X_7101_ _7646_/CLK _7101_/D fanout751/X VGND VGND VPWR VPWR _7101_/Q sky130_fd_sc_hd__dfstp_2
X_4313_ _4321_/S _4313_/B VGND VGND VPWR VPWR _4313_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3525__B _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5293_ _5168_/X _5206_/Y _5292_/Y _4428_/Y hold37/A VGND VGND VPWR VPWR _7203_/D
+ sky130_fd_sc_hd__o32a_1
XFILLER_114_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7032_ _7186_/CLK _7032_/D fanout723/X VGND VGND VPWR VPWR _7032_/Q sky130_fd_sc_hd__dfrtp_4
X_4244_ _5656_/A1 _5881_/A1 _4248_/S VGND VGND VPWR VPWR _4244_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3838__A1 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6836__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3838__B2 _7114_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5740__B _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4175_ _4175_/A input1/X VGND VGND VPWR VPWR _4175_/X sky130_fd_sc_hd__and2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3541__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6852__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4263__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6816_ _6815_/X _6816_/A1 _6822_/S VGND VGND VPWR VPWR _7642_/D sky130_fd_sc_hd__mux2_1
XFILLER_168_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6555__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6747_ _7175_/Q _6747_/B _6747_/C VGND VGND VPWR VPWR _6747_/X sky130_fd_sc_hd__and3_1
X_3959_ _7503_/Q _5983_/A _5938_/C _3955_/X _3958_/X VGND VGND VPWR VPWR _3959_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_149_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6678_ _7037_/Q _6459_/B _6769_/A3 _6423_/X _7012_/Q VGND VGND VPWR VPWR _6678_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5629_ _5629_/A0 _5645_/A0 _5629_/S VGND VGND VPWR VPWR _5629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6712__B1 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout530 _4997_/A VGND VGND VPWR VPWR _5158_/A sky130_fd_sc_hd__buf_12
Xfanout541 hold1494/X VGND VGND VPWR VPWR _4422_/A1 sky130_fd_sc_hd__buf_6
Xfanout552 _5952_/A1 VGND VGND VPWR VPWR _4544_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout563 _5996_/A1 VGND VGND VPWR VPWR _4555_/A0 sky130_fd_sc_hd__clkbuf_4
XANTENNA__6491__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout574 _5635_/A0 VGND VGND VPWR VPWR _5986_/A1 sky130_fd_sc_hd__buf_8
XFILLER_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout585 _5894_/A0 VGND VGND VPWR VPWR _5582_/A0 sky130_fd_sc_hd__buf_6
Xfanout596 _4551_/D VGND VGND VPWR VPWR _4533_/B sky130_fd_sc_hd__buf_8
XANTENNA_input131_A wb_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6243__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_9__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X VGND VGND VPWR VPWR _7633_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4254__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5754__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3765__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6701__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6703__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3517__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4221__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6909__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6482__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5690__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4493__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4176__B _4176_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6094__D _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5980_ _5980_/A0 _5980_/A1 _5982_/S VGND VGND VPWR VPWR _5980_/X sky130_fd_sc_hd__mux2_1
X_4931_ _4939_/C _4933_/A _4933_/B VGND VGND VPWR VPWR _4934_/A sky130_fd_sc_hd__and3_1
XANTENNA__5993__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7650_ _7650_/A VGND VGND VPWR VPWR _7650_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold2396_A _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4862_ _4831_/C _4574_/X _4797_/B _4669_/X _4974_/B VGND VGND VPWR VPWR _4862_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6601_ _7517_/Q _6435_/X _6446_/X _7525_/Q VGND VGND VPWR VPWR _6601_/X sky130_fd_sc_hd__a22o_1
XFILLER_178_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3813_ _7473_/Q _3931_/B _5947_/A _3617_/X _7231_/Q VGND VGND VPWR VPWR _3813_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_15 _6150_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7581_ _7581_/CLK _7581_/D fanout717/X VGND VGND VPWR VPWR _7581_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5745__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _7411_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4794_/A _5410_/B VGND VGND VPWR VPWR _4793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_37 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6532_ _7290_/Q _6422_/X _6443_/X _7450_/Q _6531_/X VGND VGND VPWR VPWR _6532_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__3756__B1 _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 _3854_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3744_ _7546_/Q _3637_/C hold90/A _3741_/X _3743_/X VGND VGND VPWR VPWR _3744_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_21_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6463_ _6463_/A _6466_/D _6468_/C VGND VGND VPWR VPWR _6463_/X sky130_fd_sc_hd__and3_4
X_3675_ _5612_/A _5596_/A _4539_/C VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__and3_4
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5414_ _5113_/A _5404_/D _5404_/C _4802_/A _5410_/A VGND VGND VPWR VPWR _5414_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_161_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6394_ _7055_/Q _6087_/X _6119_/X _7136_/Q _6393_/X VGND VGND VPWR VPWR _6397_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4181__A0 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5345_ _5343_/Y _5506_/C _4969_/Y VGND VGND VPWR VPWR _5345_/Y sky130_fd_sc_hd__a21oi_1
Xoutput177 _3434_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 _3424_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
Xhold2902 _4385_/X VGND VGND VPWR VPWR hold2902/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xoutput199 _3414_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
Xhold2913 hold2913/A VGND VGND VPWR VPWR _5843_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5276_ _5561_/A1 _5480_/B2 _4814_/Y _5102_/Y VGND VGND VPWR VPWR _5278_/B sky130_fd_sc_hd__o31a_1
XFILLER_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2924 hold2924/A VGND VGND VPWR VPWR _4268_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7015_ _7181_/CLK _7015_/D fanout721/X VGND VGND VPWR VPWR _7015_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2935 hold2935/A VGND VGND VPWR VPWR _5897_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2946 hold2946/A VGND VGND VPWR VPWR _4337_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4227_ _4256_/A0 _5998_/A1 _4231_/S VGND VGND VPWR VPWR _4227_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5276__A3 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2957 _4548_/X VGND VGND VPWR VPWR hold2957/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout381_A _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4484__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2968 _7068_/Q VGND VGND VPWR VPWR hold2968/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout479_A _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2979 hold2979/A VGND VGND VPWR VPWR hold2979/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4158_ _7257_/Q _7306_/Q _4168_/D _6881_/Q _4157_/Y VGND VGND VPWR VPWR _4158_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5897__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6225__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4089_ input118/X input119/X _4089_/C _4089_/D VGND VGND VPWR VPWR _4093_/C sky130_fd_sc_hd__and4bb_1
XANTENNA__4236__A1 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5984__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4888__A_N _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5736__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1928_A _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold3044_A _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6464__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout360 _3549_/X VGND VGND VPWR VPWR _4422_/S sky130_fd_sc_hd__buf_12
Xfanout371 _4725_/X VGND VGND VPWR VPWR _5065_/A sky130_fd_sc_hd__buf_8
XANTENNA__5672__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4475__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout382 _4078_/Y VGND VGND VPWR VPWR _6839_/B sky130_fd_sc_hd__buf_12
XFILLER_59_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout393 _4346_/C VGND VGND VPWR VPWR _3562_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA_hold3309_A _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4427__D _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4227__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__B1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6767__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5727__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__buf_4
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__buf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__buf_2
XANTENNA__3753__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR _4173_/A sky130_fd_sc_hd__buf_4
Xhold808 hold808/A VGND VGND VPWR VPWR _7050_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 spi_enabled VGND VGND VPWR VPWR _4174_/B sky130_fd_sc_hd__buf_6
Xmax_cap527 _4667_/Y VGND VGND VPWR VPWR _5024_/A1 sky130_fd_sc_hd__clkbuf_8
Xhold819 hold819/A VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6152__A1 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3460_ hold246/X _6902_/Q _4025_/A VGND VGND VPWR VPWR _3460_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5130_ _5480_/A1 _4707_/Y _4783_/Y _4625_/Y VGND VGND VPWR VPWR _5150_/A sky130_fd_sc_hd__o22a_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2209 _7329_/Q VGND VGND VPWR VPWR hold627/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5258__A3 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1508 _5863_/X VGND VGND VPWR VPWR hold203/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5061_ _5134_/A _5061_/B _5282_/C VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__and3_1
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1519 _5998_/X VGND VGND VPWR VPWR hold181/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4466__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4012_ _6892_/Q _6891_/Q VGND VGND VPWR VPWR _4123_/C sky130_fd_sc_hd__nor2_1
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ _5963_/A0 _5990_/A1 _5964_/S VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5966__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4914_ _5213_/B _5183_/C _4933_/A _4940_/D VGND VGND VPWR VPWR _4916_/A sky130_fd_sc_hd__and4_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5894_ _5894_/A0 _5894_/A1 _5901_/S VGND VGND VPWR VPWR _5894_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7633_ _7633_/CLK _7633_/D VGND VGND VPWR VPWR _7633_/Q sky130_fd_sc_hd__dfxtp_1
X_4845_ _5115_/A _5115_/B _5059_/A VGND VGND VPWR VPWR _4845_/X sky130_fd_sc_hd__and3_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7564_ _7565_/CLK _7564_/D fanout746/X VGND VGND VPWR VPWR _7564_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4776_ _4776_/A _4776_/B VGND VGND VPWR VPWR _4776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_193_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6515_ _7561_/Q _6419_/C _6443_/X _7449_/Q _6514_/X VGND VGND VPWR VPWR _6515_/X
+ sky130_fd_sc_hd__a221o_1
X_3727_ _7315_/Q _3521_/X _3723_/X _3724_/X _3726_/X VGND VGND VPWR VPWR _3727_/X
+ sky130_fd_sc_hd__a2111o_4
X_7495_ _7537_/CLK _7495_/D fanout709/X VGND VGND VPWR VPWR _7495_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__3744__A3 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6446_ _6466_/A _6466_/B _6463_/A _6466_/D VGND VGND VPWR VPWR _6446_/X sky130_fd_sc_hd__and4_4
X_3658_ _4473_/A _4455_/A _4388_/B VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__and3_2
XANTENNA__6694__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6377_ _6930_/Q _7612_/Q _4116_/X _6067_/X VGND VGND VPWR VPWR _6377_/X sky130_fd_sc_hd__o2bb2a_1
X_3589_ _7581_/Q _3501_/X _5776_/A _7389_/Q _3588_/X VGND VGND VPWR VPWR _3589_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout596_A _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5328_ _5328_/A _5328_/B _5339_/B VGND VGND VPWR VPWR _5328_/X sky130_fd_sc_hd__and3_4
XFILLER_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2710 _6877_/Q VGND VGND VPWR VPWR hold831/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2721 _4550_/X VGND VGND VPWR VPWR hold756/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2732 hold745/X VGND VGND VPWR VPWR _5642_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5259_ _4605_/Y _5563_/A1 _4744_/Y _5072_/Y VGND VGND VPWR VPWR _5265_/A sky130_fd_sc_hd__o31a_1
XANTENNA__4457__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5654__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2743 hold937/X VGND VGND VPWR VPWR _5774_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2754 _4381_/X VGND VGND VPWR VPWR hold808/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2765 _6928_/Q VGND VGND VPWR VPWR hold783/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2776 _7029_/Q VGND VGND VPWR VPWR hold851/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2787 hold875/X VGND VGND VPWR VPWR _5934_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2798 _6966_/Q VGND VGND VPWR VPWR hold865/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5406__B1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3680__A2 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5957__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1780_A _7446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3968__B1 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5421__A3 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6382__B2 _7045_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4393__A0 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6134__A1 _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6134__B2 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6685__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3499__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6437__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4448__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5645__A0 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5948__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4630_ _4570_/Y _5494_/B2 _4627_/Y VGND VGND VPWR VPWR _4767_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5176__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4384__A0 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4561_ _4562_/A _4562_/B _4562_/C _4562_/D VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__and4_4
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6300_ _7006_/Q _6082_/X _6111_/X _7036_/Q _6299_/X VGND VGND VPWR VPWR _6303_/C
+ sky130_fd_sc_hd__a221o_1
X_3512_ _5640_/A _4328_/A _3562_/C VGND VGND VPWR VPWR _5686_/A sky130_fd_sc_hd__and3_4
X_7280_ _7329_/CLK _7280_/D fanout704/X VGND VGND VPWR VPWR _7280_/Q sky130_fd_sc_hd__dfstp_4
Xhold605 hold605/A VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6125__A1 _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4492_ _4492_/A0 _5912_/A1 _4496_/S VGND VGND VPWR VPWR _4492_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6125__B2 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold616 hold616/A VGND VGND VPWR VPWR _7370_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold627 hold627/A VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold638 hold638/A VGND VGND VPWR VPWR _7345_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6231_ _7404_/Q _6091_/X _6119_/D _7356_/Q _6099_/X VGND VGND VPWR VPWR _6231_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5479__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _7521_/Q _6119_/A _6119_/B _6136_/B _6121_/C VGND VGND VPWR VPWR _6162_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2006 _4526_/X VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2017 _4553_/X VGND VGND VPWR VPWR hold446/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/A _5282_/C _5282_/D VGND VGND VPWR VPWR _5113_/X sky130_fd_sc_hd__and3_1
Xhold2028 _5700_/X VGND VGND VPWR VPWR hold398/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _7588_/Q _6081_/C _6099_/D _7589_/Q VGND VGND VPWR VPWR _6093_/X sky130_fd_sc_hd__and4bb_4
Xhold2039 hold499/X VGND VGND VPWR VPWR _5994_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4439__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1305 hold3259/X VGND VGND VPWR VPWR hold3260/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5636__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _4486_/X VGND VGND VPWR VPWR _7142_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1327 hold3216/X VGND VGND VPWR VPWR hold3217/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B _5044_/C VGND VGND VPWR VPWR _5047_/C sky130_fd_sc_hd__nand3_1
Xhold1338 _4504_/X VGND VGND VPWR VPWR _7157_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1349 _4321_/A1 VGND VGND VPWR VPWR hold2967/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5939__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4364__B _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6995_ _6999_/CLK _6995_/D VGND VGND VPWR VPWR _6995_/Q sky130_fd_sc_hd__dfxtp_1
X_5946_ _5946_/A0 hold20/X _5946_/S VGND VGND VPWR VPWR _5946_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4611__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ _5877_/A0 _5994_/A1 _5883_/S VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3965__A3 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7616_ _7621_/CLK _7616_/D fanout708/X VGND VGND VPWR VPWR _7616_/Q sky130_fd_sc_hd__dfrtp_1
X_4828_ _5399_/C _5399_/D VGND VGND VPWR VPWR _4828_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout511_A _4857_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4375__A0 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4759_ _5158_/A _5183_/A VGND VGND VPWR VPWR _4759_/Y sky130_fd_sc_hd__nand2_8
X_7547_ _7579_/CLK _7547_/D fanout732/X VGND VGND VPWR VPWR _7547_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_181_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7478_ _7478_/CLK _7478_/D fanout713/X VGND VGND VPWR VPWR _7478_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4127__A0 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6667__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6429_ _6466_/B _6441_/D _6429_/C _7594_/Q VGND VGND VPWR VPWR _6429_/X sky130_fd_sc_hd__and4b_4
XANTENNA__4539__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3230 _7187_/Q VGND VGND VPWR VPWR hold3230/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3241 hold3241/A VGND VGND VPWR VPWR _5750_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3252 _5903_/X VGND VGND VPWR VPWR hold3252/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3263 _5948_/X VGND VGND VPWR VPWR hold3263/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3274 _7215_/Q VGND VGND VPWR VPWR _3924_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2540 _7467_/Q VGND VGND VPWR VPWR hold623/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3285 _7618_/Q VGND VGND VPWR VPWR _6572_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2551 hold839/X VGND VGND VPWR VPWR _5851_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3296 _7611_/Q VGND VGND VPWR VPWR _6354_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2562 hold837/X VGND VGND VPWR VPWR _5837_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2573 _4276_/X VGND VGND VPWR VPWR hold674/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2584 _5765_/X VGND VGND VPWR VPWR hold824/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1850 _5652_/X VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2595 hold913/X VGND VGND VPWR VPWR _4470_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1861 _4476_/X VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1872 hold1872/A VGND VGND VPWR VPWR _4307_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1883 _7290_/Q VGND VGND VPWR VPWR hold269/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1894 _5717_/X VGND VGND VPWR VPWR hold337/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3956__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__A3 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6107__A1 _7295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6107__B2 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output263_A _7227_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4669__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5330__A2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3892__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__C _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__buf_6
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6291__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5995__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5800_ _5953_/A1 _5800_/A1 _5802_/S VGND VGND VPWR VPWR _5800_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6780_ _7102_/Q _6780_/B VGND VGND VPWR VPWR _6792_/S sky130_fd_sc_hd__nand2_8
XANTENNA__6594__A1 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3992_ _7367_/Q _5758_/A _5634_/A _7262_/Q _3991_/X VGND VGND VPWR VPWR _3992_/X
+ sky130_fd_sc_hd__a221o_4
X_5731_ _5731_/A _5731_/B _5947_/C VGND VGND VPWR VPWR _5739_/S sky130_fd_sc_hd__and3_4
XANTENNA__3947__A3 _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5662_ _5662_/A0 _5995_/A1 _5667_/S VGND VGND VPWR VPWR _5662_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6346__B2 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4613_ _4909_/A _4909_/C VGND VGND VPWR VPWR _4657_/B sky130_fd_sc_hd__nand2_2
X_7401_ _7542_/CLK _7401_/D fanout719/X VGND VGND VPWR VPWR _7401_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5593_ _5593_/A0 _5815_/A1 _5595_/S VGND VGND VPWR VPWR _5593_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2643_A _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7332_ _7365_/CLK _7332_/D fanout720/X VGND VGND VPWR VPWR _7332_/Q sky130_fd_sc_hd__dfrtp_4
X_4544_ _4544_/A0 _4544_/A1 _4544_/S VGND VGND VPWR VPWR _4544_/X sky130_fd_sc_hd__mux2_1
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6839__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold413 hold413/A VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold424 _4361_/X VGND VGND VPWR VPWR _7033_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold435 hold435/A VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__B2 _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7263_ _7263_/CLK _7263_/D fanout689/X VGND VGND VPWR VPWR _7263_/Q sky130_fd_sc_hd__dfrtp_1
Xhold446 hold446/A VGND VGND VPWR VPWR _7198_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4475_ _4475_/A0 _4553_/A0 _4478_/S VGND VGND VPWR VPWR _4475_/X sky130_fd_sc_hd__mux2_1
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2810_A _7140_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold468 hold468/A VGND VGND VPWR VPWR _7118_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3544__A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6214_ _6213_/Y _6212_/Y _7605_/Q _6649_/S VGND VGND VPWR VPWR _6214_/X sky130_fd_sc_hd__a2bb2o_1
X_3426_ _7434_/Q VGND VGND VPWR VPWR _3426_/Y sky130_fd_sc_hd__inv_2
Xhold479 hold479/A VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7194_ _7211_/CLK _7194_/D fanout699/X VGND VGND VPWR VPWR _7194_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5321__A2 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _6036_/Y _7280_/Q _6143_/X _6133_/X _6067_/A VGND VGND VPWR VPWR _6145_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_98_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6855__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3883__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4078__C _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 hold2983/X VGND VGND VPWR VPWR hold1102/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 hold3117/X VGND VGND VPWR VPWR hold3118/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _7511_/Q _6110_/A _6317_/C _6075_/X _7423_/Q VGND VGND VPWR VPWR _6076_/X
+ sky130_fd_sc_hd__a32o_1
Xhold1124 hold1124/A VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
Xhold1135 hold3135/X VGND VGND VPWR VPWR hold3136/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6574__B _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__A1 _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1146 _5876_/X VGND VGND VPWR VPWR _7471_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5339_/A _5203_/C _5034_/B _5339_/C VGND VGND VPWR VPWR _5028_/B sky130_fd_sc_hd__nand4_1
Xhold1157 hold1157/A VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold1168 _5631_/X VGND VGND VPWR VPWR _7256_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1179 hold2866/X VGND VGND VPWR VPWR hold2867/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3635__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_A _5726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_14_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6585__A1 _7316_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ _7636_/CLK _6978_/D VGND VGND VPWR VPWR _6978_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7476__RESET_B fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__A3 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5929_ hold77/X _5956_/C VGND VGND VPWR VPWR _5937_/S sky130_fd_sc_hd__nand2_8
XANTENNA__6337__B2 _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4899__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input161_A wb_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5312__A2 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold980 hold980/A VGND VGND VPWR VPWR _7420_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold991 hold991/A VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3060 _7243_/Q VGND VGND VPWR VPWR hold3060/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3874__A2 _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3071 _4389_/X VGND VGND VPWR VPWR hold3071/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3082 _7527_/Q VGND VGND VPWR VPWR hold3082/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3093 hold3093/A VGND VGND VPWR VPWR _5894_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2370 _7350_/Q VGND VGND VPWR VPWR hold631/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2381 _5657_/X VGND VGND VPWR VPWR hold822/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input22_A mask_rev_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2392 hold734/X VGND VGND VPWR VPWR _7337_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4285__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3626__A2 hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1680 _4253_/X VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1691 _5874_/X VGND VGND VPWR VPWR hold113/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5379__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6733__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4260_ _4260_/A0 _5732_/A1 _4264_/S VGND VGND VPWR VPWR _4260_/X sky130_fd_sc_hd__mux2_1
X_4191_ _5619_/A _5947_/A _5640_/D VGND VGND VPWR VPWR _4191_/X sky130_fd_sc_hd__and3_4
XFILLER_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6264__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6901_ _4150_/A1 _6901_/D _6851_/X VGND VGND VPWR VPWR _6901_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6832_/X sky130_fd_sc_hd__and2_1
XFILLER_23_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3975_ _7407_/Q _3493_/X _4322_/A _7001_/Q _3974_/X VGND VGND VPWR VPWR _3975_/X
+ sky130_fd_sc_hd__a221o_1
X_6763_ _7151_/Q _6408_/A _6435_/X _7050_/Q _6762_/X VGND VGND VPWR VPWR _6763_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2858_A _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5714_ _5948_/A1 _5714_/A1 _5721_/S VGND VGND VPWR VPWR _5714_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6319__A1 _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6694_ _7047_/Q _6435_/X _6452_/X _7022_/Q _6693_/X VGND VGND VPWR VPWR _6697_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_148_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5645_ _5645_/A0 _5645_/A1 _5649_/S VGND VGND VPWR VPWR _5645_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5576_ _5543_/X _5575_/Y _5550_/Y _5572_/X VGND VGND VPWR VPWR _5576_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5542__A2 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold210 hold210/A VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7315_ _7478_/CLK _7315_/D fanout714/X VGND VGND VPWR VPWR _7315_/Q sky130_fd_sc_hd__dfrtp_4
X_4527_ _4527_/A _5619_/B _5619_/C VGND VGND VPWR VPWR _4532_/S sky130_fd_sc_hd__and3_4
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold221 hold221/A VGND VGND VPWR VPWR _7572_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold232 hold232/A VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold243 hold243/A VGND VGND VPWR VPWR _6960_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold254 hold254/A VGND VGND VPWR VPWR _7190_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6098__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4458_ _4458_/A0 _5914_/A1 _4460_/S VGND VGND VPWR VPWR _4458_/X sky130_fd_sc_hd__mux2_1
Xhold276 hold276/A VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7246_ _7330_/CLK _7246_/D fanout711/X VGND VGND VPWR VPWR _7246_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold287 hold287/A VGND VGND VPWR VPWR _7268_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout701 fanout702/X VGND VGND VPWR VPWR fanout701/X sky130_fd_sc_hd__buf_4
XFILLER_120_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout712 fanout714/X VGND VGND VPWR VPWR _4079_/A sky130_fd_sc_hd__buf_8
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4502__A0 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3409_ _7256_/Q VGND VGND VPWR VPWR _3409_/Y sky130_fd_sc_hd__inv_2
Xfanout723 fanout724/X VGND VGND VPWR VPWR fanout723/X sky130_fd_sc_hd__buf_8
X_7177_ _7268_/CLK _7177_/D fanout699/X VGND VGND VPWR VPWR _7177_/Q sky130_fd_sc_hd__dfrtp_4
X_4389_ _5894_/A0 _4389_/A1 _4393_/S VGND VGND VPWR VPWR _4389_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout734 fanout736/X VGND VGND VPWR VPWR fanout734/X sky130_fd_sc_hd__buf_8
Xfanout745 fanout747/X VGND VGND VPWR VPWR fanout745/X sky130_fd_sc_hd__buf_8
Xfanout756 input127/X VGND VGND VPWR VPWR _4831_/A sky130_fd_sc_hd__buf_12
Xfanout767 input124/X VGND VGND VPWR VPWR _5407_/A1 sky130_fd_sc_hd__buf_8
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _7424_/Q _6075_/X _6121_/X _7304_/Q _6127_/X VGND VGND VPWR VPWR _6128_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6050_/Y _7598_/Q _6427_/A _6058_/X VGND VGND VPWR VPWR _6059_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_4_8__f_wb_clk_i clkbuf_3_4_0_wb_clk_i/X VGND VGND VPWR VPWR _7000_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1693_A _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A1 _7443_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4271__C _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3847__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5830__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6246__B1 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4219__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6797__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6797__B2 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6214__A2_N _6212_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5839__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3760_ _6991_/Q _4346_/C _5623_/B _3667_/X _7024_/Q VGND VGND VPWR VPWR _3760_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _7299_/Q _5965_/B _4352_/A _5794_/A _7403_/Q VGND VGND VPWR VPWR _3691_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_187_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5430_ _5429_/X _5216_/X _4997_/B VGND VGND VPWR VPWR _5554_/B sky130_fd_sc_hd__o21ai_1
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput304 _4167_/X VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
X_5361_ _5361_/A _5361_/B _5573_/B _5444_/A VGND VGND VPWR VPWR _5363_/B sky130_fd_sc_hd__and4_1
XFILLER_160_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput315 hold1150/X VGND VGND VPWR VPWR hold1151/A sky130_fd_sc_hd__buf_6
XFILLER_126_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput326 hold1098/X VGND VGND VPWR VPWR hold1099/A sky130_fd_sc_hd__buf_6
Xoutput337 hold1078/X VGND VGND VPWR VPWR hold1079/A sky130_fd_sc_hd__buf_6
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7100_ _7519_/CLK _7100_/D fanout742/X VGND VGND VPWR VPWR _7100_/Q sky130_fd_sc_hd__dfrtp_1
X_4312_ _3922_/Y _4312_/A1 _4321_/S VGND VGND VPWR VPWR _6994_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3525__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5292_ _4969_/Y _5506_/B _5288_/Y _4428_/Y _5290_/X VGND VGND VPWR VPWR _5292_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_113_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7031_ _7035_/CLK _7031_/D fanout723/X VGND VGND VPWR VPWR _7031_/Q sky130_fd_sc_hd__dfrtp_4
X_4243_ _4243_/A0 _4242_/X _4249_/S VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3838__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2606_A _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4174_ _4174_/A _4174_/B VGND VGND VPWR VPWR _4174_/X sky130_fd_sc_hd__and2_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4637__B _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3541__B _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5749__A _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6815_ _4427_/C _6815_/A2 _6815_/B1 wire536/A _6814_/X VGND VGND VPWR VPWR _6815_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6746_ _7039_/Q _6459_/B _6769_/A3 _6463_/X _7165_/Q VGND VGND VPWR VPWR _6746_/X
+ sky130_fd_sc_hd__a32o_1
X_3958_ _7519_/Q _5785_/B _4376_/B _3957_/X VGND VGND VPWR VPWR _3958_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3889_ _7245_/Q _5731_/A _5614_/B _5713_/A _7328_/Q VGND VGND VPWR VPWR _3889_/X
+ sky130_fd_sc_hd__a32o_4
X_6677_ _7178_/Q _6058_/X _6409_/X _7133_/Q VGND VGND VPWR VPWR _6677_/X sky130_fd_sc_hd__a22o_1
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5628_ _5628_/A0 _5954_/A1 _5629_/S VGND VGND VPWR VPWR _5628_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6173__C1 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6712__B2 _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5559_ _5559_/A _5559_/B _5559_/C _5559_/D VGND VGND VPWR VPWR _5560_/C sky130_fd_sc_hd__nor4_1
XFILLER_117_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7229_ _7232_/CLK _7229_/D fanout689/X VGND VGND VPWR VPWR _7229_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout520 _4721_/Y VGND VGND VPWR VPWR _5059_/B sky130_fd_sc_hd__buf_8
XANTENNA__3829__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout531 _4605_/Y VGND VGND VPWR VPWR _5495_/C1 sky130_fd_sc_hd__buf_6
Xfanout542 _5972_/A1 VGND VGND VPWR VPWR _5954_/A1 sky130_fd_sc_hd__buf_8
Xfanout553 _5673_/A0 VGND VGND VPWR VPWR _5952_/A1 sky130_fd_sc_hd__buf_8
Xfanout564 _5969_/A1 VGND VGND VPWR VPWR _5978_/A0 sky130_fd_sc_hd__clkbuf_8
Xfanout575 hold198/X VGND VGND VPWR VPWR _5645_/A0 sky130_fd_sc_hd__buf_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout586 hold487/X VGND VGND VPWR VPWR _5894_/A0 sky130_fd_sc_hd__buf_12
Xfanout597 hold26/X VGND VGND VPWR VPWR _4551_/D sky130_fd_sc_hd__buf_12
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7491__RESET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input124_A wb_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__A _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6400__B1 _6398_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6703__A1 _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3517__A1 _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4190__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6219__B1 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5690__A1 hold365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4930_ _4930_/A _4930_/B _4930_/C VGND VGND VPWR VPWR _4934_/C sky130_fd_sc_hd__nand3_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _4861_/A _4861_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _4861_/X sky130_fd_sc_hd__and4_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6600_ _7501_/Q _6600_/B _6651_/C VGND VGND VPWR VPWR _6600_/X sky130_fd_sc_hd__and3_1
XFILLER_177_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3812_ _7489_/Q _5893_/A _3669_/X _6969_/Q _3811_/X VGND VGND VPWR VPWR _3812_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_16 _6283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7580_ _7580_/CLK _7580_/D fanout735/X VGND VGND VPWR VPWR _7580_/Q sky130_fd_sc_hd__dfrtp_4
X_4792_ _4700_/Y _4789_/Y _4791_/Y VGND VGND VPWR VPWR _4800_/C sky130_fd_sc_hd__o21ai_1
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_27 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_38 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3756__A1 _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _4093_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ _7434_/Q _6747_/B _6747_/C _6447_/X _7442_/Q VGND VGND VPWR VPWR _6531_/X
+ sky130_fd_sc_hd__a32o_1
X_3743_ _7562_/Q _5974_/A _4231_/S input38/X _3742_/X VGND VGND VPWR VPWR _3743_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3756__B2 input46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4412__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6462_ _6466_/B _6463_/A _6462_/C _6466_/A VGND VGND VPWR VPWR _6462_/X sky130_fd_sc_hd__and4b_4
X_3674_ _5830_/C _4515_/B _4539_/C VGND VGND VPWR VPWR _5581_/A sky130_fd_sc_hd__and3_4
XFILLER_118_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5413_ _5538_/B _5569_/A _5568_/A _5488_/B VGND VGND VPWR VPWR _5416_/B sky130_fd_sc_hd__and4_1
X_6393_ _7213_/Q _6317_/B _6089_/X _6092_/X _7181_/Q VGND VGND VPWR VPWR _6393_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6170__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5344_ _5058_/D _5073_/A _4846_/Y _5204_/X VGND VGND VPWR VPWR _5506_/C sky130_fd_sc_hd__o31a_1
XFILLER_142_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6458__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput178 _3433_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 _3423_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ _5561_/A1 _4806_/Y _5255_/X _5274_/X VGND VGND VPWR VPWR _5278_/C sky130_fd_sc_hd__o31a_1
XFILLER_153_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2903 _7648_/A VGND VGND VPWR VPWR hold2903/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2914 _7522_/Q VGND VGND VPWR VPWR hold2914/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3552__A _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2925 _4268_/X VGND VGND VPWR VPWR hold2925/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7014_ _7212_/CLK _7014_/D fanout723/X VGND VGND VPWR VPWR _7014_/Q sky130_fd_sc_hd__dfrtp_4
X_4226_ _4226_/A0 _4225_/X _4232_/S VGND VGND VPWR VPWR _4226_/X sky130_fd_sc_hd__mux2_1
Xhold2936 _5897_/X VGND VGND VPWR VPWR hold2936/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6473__A3 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2947 _4337_/X VGND VGND VPWR VPWR hold2947/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2958 _7058_/Q VGND VGND VPWR VPWR hold2958/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5681__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2969 hold2969/A VGND VGND VPWR VPWR _4403_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4157_ _7257_/Q _7306_/Q _4168_/D _7290_/Q VGND VGND VPWR VPWR _4157_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6225__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4088_ _4825_/A _4674_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4088_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_102_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout541_A hold1494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4814__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3747__A1 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6729_ _7014_/Q _4105_/B _6459_/B _6422_/X _6965_/Q VGND VGND VPWR VPWR _6729_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_csclk _7399_/CLK VGND VGND VPWR VPWR _7421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6161__A2 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6449__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7497_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout361 _4527_/A VGND VGND VPWR VPWR _4539_/C sky130_fd_sc_hd__buf_8
Xfanout372 _5453_/A VGND VGND VPWR VPWR _5213_/B sky130_fd_sc_hd__buf_2
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout383 _4364_/B VGND VGND VPWR VPWR _5623_/B sky130_fd_sc_hd__clkbuf_16
Xfanout394 hold250/X VGND VGND VPWR VPWR _4346_/C sky130_fd_sc_hd__buf_8
XFILLER_59_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6216__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5424__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_62_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3637__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR _4175_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_168_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_4
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR _4076_/B sky130_fd_sc_hd__buf_12
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold809 hold809/A VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap528 _4730_/C VGND VGND VPWR VPWR _4801_/B sky130_fd_sc_hd__buf_4
XANTENNA__6152__A2 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3910__A1 _7496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5060_ _5060_/A _5060_/B _5060_/C VGND VGND VPWR VPWR _5064_/A sky130_fd_sc_hd__nor3_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 hold203/X VGND VGND VPWR VPWR _7460_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5998__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5663__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4011_ _6910_/Q _6909_/Q _6908_/Q _7073_/Q VGND VGND VPWR VPWR _4011_/X sky130_fd_sc_hd__and4_2
XFILLER_93_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4915__B _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5415__B2 _4759_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5962_ _5962_/A0 _5998_/A1 _5964_/S VGND VGND VPWR VPWR _5962_/X sky130_fd_sc_hd__mux2_1
X_4913_ _4913_/A _4913_/B _4913_/C VGND VGND VPWR VPWR _4916_/C sky130_fd_sc_hd__nand3_1
X_5893_ _5893_/A _5893_/B VGND VGND VPWR VPWR _5901_/S sky130_fd_sc_hd__nand2_8
X_7632_ _7636_/CLK _7632_/D VGND VGND VPWR VPWR _7632_/Q sky130_fd_sc_hd__dfxtp_1
X_4844_ _4748_/A _4844_/B _5091_/A VGND VGND VPWR VPWR _4844_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__6376__C1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7563_ _7563_/CLK _7563_/D fanout739/X VGND VGND VPWR VPWR _7563_/Q sky130_fd_sc_hd__dfrtp_2
X_4775_ _5107_/C _5059_/B _4775_/C VGND VGND VPWR VPWR _4776_/A sky130_fd_sc_hd__and3_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6514_ _7441_/Q _6574_/B _6771_/A3 _6513_/X VGND VGND VPWR VPWR _6514_/X sky130_fd_sc_hd__a31o_1
X_3726_ _7307_/Q _5686_/A _3667_/X _7025_/Q _3725_/X VGND VGND VPWR VPWR _3726_/X
+ sky130_fd_sc_hd__a221o_1
X_7494_ _7576_/CLK _7494_/D fanout718/X VGND VGND VPWR VPWR _7494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6679__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6445_ _7535_/Q _6408_/D _6420_/A _7295_/Q _6444_/X VGND VGND VPWR VPWR _6445_/X
+ sky130_fd_sc_hd__a221o_1
X_3657_ _5640_/B _5596_/A _5640_/C VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__and3_4
XFILLER_134_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4154__A1 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5351__B1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6376_ _6960_/Q _6036_/Y _6362_/Y _6375_/X _6067_/A VGND VGND VPWR VPWR _6376_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3588_ _7541_/Q _3590_/C _4527_/A _3544_/X _7421_/Q VGND VGND VPWR VPWR _3588_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5327_ _5058_/D _5072_/B _5203_/C _5049_/C VGND VGND VPWR VPWR _5339_/B sky130_fd_sc_hd__a211o_4
XANTENNA_fanout491_A _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2700 _7054_/Q VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout589_A hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2711 hold831/X VGND VGND VPWR VPWR _4188_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2722 _7175_/Q VGND VGND VPWR VPWR hold763/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5258_ _5260_/C _5387_/D _5061_/B _5257_/X VGND VGND VPWR VPWR _5266_/A sky130_fd_sc_hd__a31o_1
Xhold2733 _5642_/X VGND VGND VPWR VPWR hold746/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2744 _7230_/Q VGND VGND VPWR VPWR hold793/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2755 _7200_/Q VGND VGND VPWR VPWR hold951/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4209_ _4209_/A0 _5627_/A1 _4211_/S VGND VGND VPWR VPWR _4209_/X sky130_fd_sc_hd__mux2_1
Xhold2766 hold783/X VGND VGND VPWR VPWR _4214_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5189_ _4924_/B _5180_/B _5034_/C _5031_/B VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__a31o_1
Xhold2777 hold851/X VGND VGND VPWR VPWR _4356_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5701__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2788 _7115_/Q VGND VGND VPWR VPWR hold969/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2799 hold865/X VGND VGND VPWR VPWR _4270_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6603__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3968__A1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6382__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6134__A2 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4145__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3154_A _7182_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input52_A mgmt_gpio_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_605 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4227__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3959__A1 _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6373__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5176__A3 _4971_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4560_ _4825_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4788_/C sky130_fd_sc_hd__nor3_4
X_3511_ _3511_/A hold46/X _3511_/C VGND VGND VPWR VPWR _3563_/C sky130_fd_sc_hd__and3_4
XFILLER_144_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 hold606/A VGND VGND VPWR VPWR _7060_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4491_ _4515_/B _5965_/A _4491_/C _4551_/D VGND VGND VPWR VPWR _4496_/S sky130_fd_sc_hd__and4_4
XFILLER_156_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold617 hold617/A VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold628 hold628/A VGND VGND VPWR VPWR _7329_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold639 hold639/A VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3442_ _7298_/Q VGND VGND VPWR VPWR _3442_/Y sky130_fd_sc_hd__inv_2
X_6230_ _7476_/Q _6032_/Y _6081_/X _7452_/Q _6229_/X VGND VGND VPWR VPWR _6230_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_170_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ _7361_/Q _6332_/C _6158_/X _6160_/X VGND VGND VPWR VPWR _6161_/X sky130_fd_sc_hd__a211o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__B1 _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2007 _7456_/Q VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _4828_/Y _5528_/A3 _5200_/C _4840_/D _5111_/Y VGND VGND VPWR VPWR _5112_/X
+ sky130_fd_sc_hd__o221a_1
Xhold2018 _7113_/Q VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2029 _7322_/Q VGND VGND VPWR VPWR hold443/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6092_ _6112_/C _6119_/A _6119_/B _6121_/A VGND VGND VPWR VPWR _6092_/X sky130_fd_sc_hd__and4_4
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 _4192_/X VGND VGND VPWR VPWR _6911_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1317 hold3152/X VGND VGND VPWR VPWR hold3153/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5043_ _4984_/B _4984_/A _4672_/X _4660_/Y _4759_/Y VGND VGND VPWR VPWR _5044_/B
+ sky130_fd_sc_hd__a2111o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 hold3218/X VGND VGND VPWR VPWR _7051_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1339 hold3208/X VGND VGND VPWR VPWR hold3209/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4926__A _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_wbbd_sck _7645_/Q VGND VGND VPWR VPWR clkbuf_0_wbbd_sck/X sky130_fd_sc_hd__clkbuf_16
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6994_ _6999_/CLK _6994_/D VGND VGND VPWR VPWR _6994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5945_ _5945_/A0 _5990_/A1 _5946_/S VGND VGND VPWR VPWR _5945_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5876_ _5876_/A0 _5876_/A1 _5883_/S VGND VGND VPWR VPWR _5876_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7615_ _7621_/CLK _7615_/D fanout707/X VGND VGND VPWR VPWR _7615_/Q sky130_fd_sc_hd__dfrtp_1
X_4827_ _5115_/A _5115_/B _4983_/C VGND VGND VPWR VPWR _4827_/X sky130_fd_sc_hd__and3_1
XANTENNA__6364__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7546_ _7573_/CLK _7546_/D fanout734/X VGND VGND VPWR VPWR _7546_/Q sky130_fd_sc_hd__dfrtp_4
X_4758_ _5158_/A _5012_/A _5328_/B VGND VGND VPWR VPWR _4758_/X sky130_fd_sc_hd__and3_4
XFILLER_119_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ _7151_/Q _3652_/X _3654_/X _7121_/Q _3655_/X VGND VGND VPWR VPWR _3709_/X
+ sky130_fd_sc_hd__a221o_1
X_7477_ _7478_/CLK _7477_/D fanout720/X VGND VGND VPWR VPWR _7477_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_10_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4689_ _4679_/C _4679_/A _5328_/B VGND VGND VPWR VPWR _4689_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__4127__A1 _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ _7594_/Q _6433_/D _6441_/D _6429_/C VGND VGND VPWR VPWR _6428_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__6667__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6100__B _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6359_ _7155_/Q _6072_/X _6099_/X _7029_/Q _6358_/X VGND VGND VPWR VPWR _6362_/B
+ sky130_fd_sc_hd__a221oi_4
Xhold3220 hold3220/A VGND VGND VPWR VPWR hold3220/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4539__C _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3231 hold3231/A VGND VGND VPWR VPWR _4540_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold1521_A _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3242 _7407_/Q VGND VGND VPWR VPWR hold3242/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3253 _7235_/Q VGND VGND VPWR VPWR hold3253/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3264 _7633_/Q VGND VGND VPWR VPWR _6788_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2530 hold841/X VGND VGND VPWR VPWR _5842_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3275 _7216_/Q VGND VGND VPWR VPWR _3858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2541 hold623/X VGND VGND VPWR VPWR _5871_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3286 _6548_/X VGND VGND VPWR VPWR _7618_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2552 _5851_/X VGND VGND VPWR VPWR hold840/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3297 _7624_/Q VGND VGND VPWR VPWR _6726_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2563 _5837_/X VGND VGND VPWR VPWR hold838/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2574 _7141_/Q VGND VGND VPWR VPWR hold737/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__B1 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1840 _7064_/Q VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2585 _7413_/Q VGND VGND VPWR VPWR hold847/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2596 _4470_/X VGND VGND VPWR VPWR hold914/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1851 _7352_/Q VGND VGND VPWR VPWR hold357/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1862 _7499_/Q VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1873 _4307_/X VGND VGND VPWR VPWR hold252/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1884 hold269/X VGND VGND VPWR VPWR _5672_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1895 _7392_/Q VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5089__D _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4571__A _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6355__A2 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4366__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6107__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6658__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output256_A _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__B1 _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5618__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4168__D _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3892__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3629__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3650__A _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6594__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3991_ _7375_/Q _5740_/A _5983_/A _3658_/X _7112_/Q VGND VGND VPWR VPWR _3991_/X
+ sky130_fd_sc_hd__a32o_1
X_5730_ _5730_/A0 hold20/X _5730_/S VGND VGND VPWR VPWR _5730_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3801__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5661_ _5661_/A0 _5949_/A1 _5667_/S VGND VGND VPWR VPWR _5661_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6346__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5149__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7400_ _7542_/CLK _7400_/D fanout709/X VGND VGND VPWR VPWR _7400_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4357__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4612_ _4571_/Y _5387_/B _4814_/C VGND VGND VPWR VPWR _4909_/C sky130_fd_sc_hd__o21ai_4
XANTENNA_hold2469_A _6876_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5592_ _5592_/A0 _5645_/A0 _5595_/S VGND VGND VPWR VPWR _5592_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7331_ _7360_/CLK _7331_/D fanout703/X VGND VGND VPWR VPWR _7331_/Q sky130_fd_sc_hd__dfrtp_4
X_4543_ _4543_/A0 _5647_/A0 _4544_/S VGND VGND VPWR VPWR _4543_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold403 hold403/A VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold414 hold414/A VGND VGND VPWR VPWR _7272_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4109__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4420__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold425 hold425/A VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold436 hold436/A VGND VGND VPWR VPWR _7480_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3580__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7262_ _7578_/CLK _7262_/D fanout747/X VGND VGND VPWR VPWR _7262_/Q sky130_fd_sc_hd__dfrtp_4
X_4474_ _4474_/A0 _5876_/A1 _4478_/S VGND VGND VPWR VPWR _4474_/X sky130_fd_sc_hd__mux2_1
Xhold447 hold447/A VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3544__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold458 _5787_/X VGND VGND VPWR VPWR _7392_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6213_ _7283_/Q _6036_/Y _6623_/B1 VGND VGND VPWR VPWR _6213_/Y sky130_fd_sc_hd__o21ai_1
Xhold469 hold469/A VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3425_ _7442_/Q VGND VGND VPWR VPWR _3425_/Y sky130_fd_sc_hd__inv_2
X_7193_ _7212_/CLK _7193_/D fanout721/X VGND VGND VPWR VPWR _7193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3868__B1 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _6144_/A _6144_/B _6144_/C VGND VGND VPWR VPWR _6144_/X sky130_fd_sc_hd__and3_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 hold1103/A VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
XANTENNA__3883__A3 _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1114 _4272_/X VGND VGND VPWR VPWR _6967_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6136_/B _6144_/B VGND VGND VPWR VPWR _6075_/X sky130_fd_sc_hd__and3_4
XFILLER_112_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X VGND VGND VPWR VPWR _7610_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 hold3108/X VGND VGND VPWR VPWR hold3109/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1136 hold3137/X VGND VGND VPWR VPWR _7122_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6574__C _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1147 hold3029/X VGND VGND VPWR VPWR hold1147/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5026_ _5026_/A _5026_/B _5026_/C VGND VGND VPWR VPWR _5028_/A sky130_fd_sc_hd__nor3_1
Xhold1158 hold3148/X VGND VGND VPWR VPWR hold3149/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1169 hold3116/X VGND VGND VPWR VPWR hold1169/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4293__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3635__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6871__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7636_/CLK _6977_/D VGND VGND VPWR VPWR _6977_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6585__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5928_ _5991_/A1 hold52/X _5928_/S VGND VGND VPWR VPWR _5928_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6894__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout719_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__A4 _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4822__C _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6337__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5859_ _5994_/A1 _5859_/A1 _5865_/S VGND VGND VPWR VPWR _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4348__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7529_ _7563_/CLK _7529_/D fanout740/X VGND VGND VPWR VPWR _7529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold970 hold970/A VGND VGND VPWR VPWR _7115_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold981 hold981/A VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1903_A _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold992 hold992/A VGND VGND VPWR VPWR _7130_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input154_A wb_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4520__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3050 _5639_/X VGND VGND VPWR VPWR hold3050/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3061 hold3061/A VGND VGND VPWR VPWR _5613_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3874__A3 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3072 _7011_/Q VGND VGND VPWR VPWR hold3072/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3083 hold3083/A VGND VGND VPWR VPWR _5939_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3094 _5894_/X VGND VGND VPWR VPWR hold3094/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2360 _4255_/X VGND VGND VPWR VPWR hold546/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2371 hold631/X VGND VGND VPWR VPWR _5739_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2382 _7555_/Q VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2393 _7371_/Q VGND VGND VPWR VPWR hold583/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1670 _5869_/X VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input15_A mask_rev_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3626__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1681 _7202_/Q VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6781__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1692 hold113/X VGND VGND VPWR VPWR _7470_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6025__A1 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6576__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5784__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4339__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4240__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4511__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4190_ _4190_/A0 _5853_/A0 _4190_/S VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4907__C _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6264__A1 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6264__B2 _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6900_ _4127_/A1 _6900_/D _6850_/X VGND VGND VPWR VPWR _6900_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6831_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6831_/X sky130_fd_sc_hd__and2_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6567__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4415__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6762_ _7186_/Q _6574_/B _6771_/A3 _6468_/X _7146_/Q VGND VGND VPWR VPWR _6762_/X
+ sky130_fd_sc_hd__a32o_1
X_3974_ _6957_/Q _3657_/X _4485_/A _7142_/Q VGND VGND VPWR VPWR _3974_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5100__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5713_ _5713_/A _5947_/C VGND VGND VPWR VPWR _5721_/S sky130_fd_sc_hd__nand2_8
XFILLER_188_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6693_ _7067_/Q _4101_/X _6441_/X _6466_/X _7210_/Q VGND VGND VPWR VPWR _6693_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6319__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ _5732_/A1 _5644_/A1 _5649_/S VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5575_ _5575_/A _5575_/B _5575_/C VGND VGND VPWR VPWR _5575_/Y sky130_fd_sc_hd__nand3_2
XFILLER_163_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5542__A3 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold200 hold200/A VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3555__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7314_ _7314_/CLK _7314_/D _4079_/A VGND VGND VPWR VPWR _7314_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4150__S _6898_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold211 hold211/A VGND VGND VPWR VPWR _7481_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4526_ _4526_/A0 _5826_/A1 _4526_/S VGND VGND VPWR VPWR _4526_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold244 hold244/A VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7245_ _7330_/CLK _7245_/D fanout711/X VGND VGND VPWR VPWR _7245_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_171_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4457_ _4457_/A0 _4553_/A0 _4460_/S VGND VGND VPWR VPWR _4457_/X sky130_fd_sc_hd__mux2_1
Xhold266 hold266/A VGND VGND VPWR VPWR _7275_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold277 hold277/A VGND VGND VPWR VPWR _7298_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold288 _7247_/Q VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout702 fanout750/X VGND VGND VPWR VPWR fanout702/X sky130_fd_sc_hd__buf_6
Xhold299 _4538_/X VGND VGND VPWR VPWR _7186_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3408_ _6009_/B VGND VGND VPWR VPWR _3408_/Y sky130_fd_sc_hd__clkinv_2
Xfanout713 fanout720/X VGND VGND VPWR VPWR fanout713/X sky130_fd_sc_hd__buf_8
XFILLER_172_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout724 fanout728/X VGND VGND VPWR VPWR fanout724/X sky130_fd_sc_hd__buf_8
X_7176_ _7176_/CLK _7176_/D fanout722/X VGND VGND VPWR VPWR _7176_/Q sky130_fd_sc_hd__dfrtp_4
X_4388_ _4527_/A _4388_/B _5596_/B _5619_/C VGND VGND VPWR VPWR _4393_/S sky130_fd_sc_hd__nand4_4
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout735 fanout736/X VGND VGND VPWR VPWR fanout735/X sky130_fd_sc_hd__clkbuf_8
Xfanout746 fanout747/X VGND VGND VPWR VPWR fanout746/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout757 input127/X VGND VGND VPWR VPWR _4786_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA_input7_A mask_rev_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _7496_/Q _6075_/A _6084_/X _6120_/X _7336_/Q VGND VGND VPWR VPWR _6127_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A _5635_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout768 _4844_/B VGND VGND VPWR VPWR _4888_/C sky130_fd_sc_hd__buf_12
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6441_/D _6433_/D _6747_/B VGND VGND VPWR VPWR _6058_/X sky130_fd_sc_hd__and3_4
XTAP_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4596__A_N _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5009_ _5024_/A1 _4669_/X _4996_/A _4974_/B VGND VGND VPWR VPWR _5013_/C sky130_fd_sc_hd__o211a_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1686_A _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5766__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6106__A _7591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__A2 _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7072__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4271__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6730__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3067_A _7295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_760 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6479__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3847__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4296__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6246__A1 _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2190 _7497_/Q VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5839__B _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4743__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6549__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4235__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3783__A2 _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3690_ _7331_/Q _5785_/B _4352_/A _3666_/X _7015_/Q VGND VGND VPWR VPWR _3690_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6182__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5360_ _5213_/A _4924_/B _5346_/X _5231_/C VGND VGND VPWR VPWR _5444_/A sky130_fd_sc_hd__a31oi_2
Xoutput305 _4166_/X VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput316 hold1102/X VGND VGND VPWR VPWR hold1103/A sky130_fd_sc_hd__buf_6
XFILLER_160_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput327 hold2965/X VGND VGND VPWR VPWR hold1093/A sky130_fd_sc_hd__buf_6
X_4311_ _4321_/S _3996_/B _4310_/Y VGND VGND VPWR VPWR _6993_/D sky130_fd_sc_hd__o21ai_1
Xoutput338 hold1169/X VGND VGND VPWR VPWR hold1170/A sky130_fd_sc_hd__buf_6
X_5291_ _4821_/Y _4858_/Y _4672_/X _4873_/X _4679_/Y VGND VGND VPWR VPWR _5506_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5590__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6485__A1 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7030_ _7035_/CLK _7030_/D fanout723/X VGND VGND VPWR VPWR _7030_/Q sky130_fd_sc_hd__dfrtp_4
X_4242_ _5655_/A1 _5952_/A1 _4248_/S VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4918__B _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3838__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4173_ _4173_/A _4173_/B VGND VGND VPWR VPWR _4173_/X sky130_fd_sc_hd__and2_1
XANTENNA__6625__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5460__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6814_ _4427_/D _6814_/A2 _6814_/B1 _4427_/B VGND VGND VPWR VPWR _6814_/X sky130_fd_sc_hd__a22o_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ _7212_/Q _6466_/X _6467_/X _7155_/Q _6744_/X VGND VGND VPWR VPWR _6745_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3957_ _7479_/Q _3535_/X _3673_/X _7197_/Q _3956_/X VGND VGND VPWR VPWR _3957_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4971__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3774__A2 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6676_ _6675_/X _6700_/A2 _6777_/S VGND VGND VPWR VPWR _6676_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout417_A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3888_ _7512_/Q _5920_/A _3881_/X _3884_/X _3887_/X VGND VGND VPWR VPWR _3888_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_5627_ _5627_/A0 _5627_/A1 _5629_/S VGND VGND VPWR VPWR _5627_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6173__B1 _6089_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6712__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5558_ _5061_/B _4827_/X _5115_/X _4645_/D _5324_/A VGND VGND VPWR VPWR _5559_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_132_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4509_ _4551_/B _4515_/B _4509_/C _4533_/B VGND VGND VPWR VPWR _4514_/S sky130_fd_sc_hd__and4_4
XFILLER_117_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5489_ _5038_/A _5127_/A _4831_/Y _5164_/A VGND VGND VPWR VPWR _5489_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6476__A1 _7520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7228_ _7232_/CLK _7228_/D _4128_/B VGND VGND VPWR VPWR _7228_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6476__B2 _7440_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__A0 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout510 _4857_/X VGND VGND VPWR VPWR _5183_/C sky130_fd_sc_hd__buf_8
XFILLER_104_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout532 _4600_/Y VGND VGND VPWR VPWR _5222_/A sky130_fd_sc_hd__buf_8
XFILLER_59_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout543 _5972_/A1 VGND VGND VPWR VPWR _5999_/A1 sky130_fd_sc_hd__clkbuf_8
X_7159_ _7268_/CLK _7159_/D _6861_/A VGND VGND VPWR VPWR _7159_/Q sky130_fd_sc_hd__dfstp_2
Xfanout554 _5826_/A1 VGND VGND VPWR VPWR _5817_/A1 sky130_fd_sc_hd__buf_6
Xfanout565 _5996_/A1 VGND VGND VPWR VPWR _5969_/A1 sky130_fd_sc_hd__buf_8
XANTENNA_hold1601_A _7517_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout576 hold1567/X VGND VGND VPWR VPWR hold198/A sky130_fd_sc_hd__buf_6
Xfanout587 hold487/X VGND VGND VPWR VPWR _5876_/A1 sky130_fd_sc_hd__buf_8
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout598 _5992_/D VGND VGND VPWR VPWR _5956_/C sky130_fd_sc_hd__buf_12
XFILLER_46_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__B _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input117_A wb_adr_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7217__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3765__A2 _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input82_A spi_sdoenb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6164__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3517__A2 _3515_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4761__A_N _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_795 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6219__A1 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4473__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4860_ _4860_/A _4860_/B VGND VGND VPWR VPWR _4860_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _7289_/Q hold90/A _4346_/C _3666_/X _7013_/Q VGND VGND VPWR VPWR _3811_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_60_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4791_ _4791_/A _4791_/B VGND VGND VPWR VPWR _4791_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 _6440_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _7671_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6530_ _7554_/Q _6408_/A _6463_/X _7426_/Q VGND VGND VPWR VPWR _6530_/X sky130_fd_sc_hd__a22o_1
X_3742_ _7140_/Q _5965_/A _4364_/B _3531_/X _7338_/Q VGND VGND VPWR VPWR _3742_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3756__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4920__C _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6155__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6461_ _7383_/Q _6460_/X _6459_/X _6458_/X _6456_/X VGND VGND VPWR VPWR _6471_/B
+ sky130_fd_sc_hd__a2111o_1
X_3673_ _4551_/A _4551_/B _4551_/C VGND VGND VPWR VPWR _3673_/X sky130_fd_sc_hd__and3_2
XFILLER_146_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5412_ _5406_/Y _4783_/Y _5150_/A _5311_/B VGND VGND VPWR VPWR _5488_/B sky130_fd_sc_hd__o211a_1
X_6392_ _7186_/Q _6097_/X _6110_/X _7176_/Q _6391_/X VGND VGND VPWR VPWR _6397_/B
+ sky130_fd_sc_hd__a221o_1
X_5343_ _5343_/A _5343_/B _5343_/C VGND VGND VPWR VPWR _5343_/Y sky130_fd_sc_hd__nor3_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput179 _3432_/Y VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
XANTENNA__4469__A0 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5274_ _5255_/X _4798_/Y _5476_/A _5272_/X VGND VGND VPWR VPWR _5274_/X sky130_fd_sc_hd__o211a_1
Xhold2904 hold2904/A VGND VGND VPWR VPWR _5621_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_99_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2915 hold2915/A VGND VGND VPWR VPWR _5933_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3552__B _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7013_ _7179_/CLK _7013_/D fanout698/X VGND VGND VPWR VPWR _7013_/Q sky130_fd_sc_hd__dfstp_2
Xhold2926 _6990_/Q VGND VGND VPWR VPWR hold2926/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4225_ _4255_/A0 _5997_/A1 _4231_/S VGND VGND VPWR VPWR _4225_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5130__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2937 _7018_/Q VGND VGND VPWR VPWR hold2937/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2948 _7164_/Q VGND VGND VPWR VPWR hold2948/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2959 hold2959/A VGND VGND VPWR VPWR _4391_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4156_ _6941_/Q input3/X input1/X VGND VGND VPWR VPWR _4156_/X sky130_fd_sc_hd__mux2_4
XFILLER_55_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4087_ _5071_/B _5071_/C VGND VGND VPWR VPWR _5115_/A sky130_fd_sc_hd__nor2_8
XFILLER_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout367_A hold31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6394__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4989_ _5029_/A _5038_/B _5038_/C VGND VGND VPWR VPWR _5039_/A sky130_fd_sc_hd__and3_1
X_6728_ _7593_/Q _7120_/Q _6408_/C _6409_/X _7135_/Q VGND VGND VPWR VPWR _6728_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_183_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6146__B1 _4116_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6659_ _7011_/Q _6423_/X _6462_/X _7031_/Q _6658_/X VGND VGND VPWR VPWR _6659_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_5 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6449__A1 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout362 _4527_/A VGND VGND VPWR VPWR _5947_/B sky130_fd_sc_hd__buf_8
Xfanout373 _4725_/X VGND VGND VPWR VPWR _5453_/A sky130_fd_sc_hd__clkbuf_8
Xfanout384 _3576_/X VGND VGND VPWR VPWR _4364_/B sky130_fd_sc_hd__buf_12
XFILLER_101_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout395 hold250/X VGND VGND VPWR VPWR _4352_/A sky130_fd_sc_hd__buf_8
XFILLER_74_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6621__A1 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5424__A2 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4740__C _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_2
XFILLER_7_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3637__B _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__buf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3653__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3910__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5112__B2 _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4010_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _4010_/Y sky130_fd_sc_hd__nand3_1
XFILLER_96_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6612__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5961_ _5961_/A0 _5997_/A1 _5964_/S VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__mux2_1
X_4912_ _4943_/B _4915_/C VGND VGND VPWR VPWR _4913_/C sky130_fd_sc_hd__nand2_1
XANTENNA_hold2499_A _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3977__A2 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5892_ _5892_/A0 _5991_/A1 hold91/X VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold90_A hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7631_ _7636_/CLK _7631_/D VGND VGND VPWR VPWR _7631_/Q sky130_fd_sc_hd__dfxtp_1
X_4843_ _4843_/A _5073_/B VGND VGND VPWR VPWR _5067_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4423__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3729__A2 _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7562_ _7562_/CLK _7562_/D fanout740/X VGND VGND VPWR VPWR _7562_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_159_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4774_ _4778_/B _4775_/C VGND VGND VPWR VPWR _4774_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__6391__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6513_ _7465_/Q _6434_/B _6771_/A3 _6466_/X _7505_/Q VGND VGND VPWR VPWR _6513_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6128__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3725_ _7259_/Q _3738_/B _4265_/B _4497_/A _7156_/Q VGND VGND VPWR VPWR _3725_/X
+ sky130_fd_sc_hd__a32o_4
X_7493_ _7582_/CLK _7493_/D fanout717/X VGND VGND VPWR VPWR _7493_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_hold2833_A _7367_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6444_ _7447_/Q _6467_/A _6574_/C _6423_/X _7327_/Q VGND VGND VPWR VPWR _6444_/X
+ sky130_fd_sc_hd__a32o_1
X_3656_ _4473_/A _4455_/A _4515_/B VGND VGND VPWR VPWR _4370_/A sky130_fd_sc_hd__and3_4
XFILLER_161_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5351__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6375_ _6317_/B _6365_/X _6370_/X _6374_/X VGND VGND VPWR VPWR _6375_/X sky130_fd_sc_hd__a211o_4
X_3587_ _3587_/A _3587_/B _3587_/C _3587_/D VGND VGND VPWR VPWR _3607_/B sky130_fd_sc_hd__nor4_2
XANTENNA__3563__A _7302_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5326_ _4672_/X _4980_/X _5174_/Y _5325_/X VGND VGND VPWR VPWR _5423_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3901__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2701 hold849/X VGND VGND VPWR VPWR _4386_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2712 _4188_/X VGND VGND VPWR VPWR hold832/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5257_ _5255_/X _5077_/Y _4765_/B _4803_/A VGND VGND VPWR VPWR _5257_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_57_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2723 hold763/X VGND VGND VPWR VPWR _4525_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2734 _7379_/Q VGND VGND VPWR VPWR hold813/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2745 hold793/X VGND VGND VPWR VPWR _5598_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2756 hold951/X VGND VGND VPWR VPWR _4555_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4208_ _4208_/A0 _5736_/A1 _4211_/S VGND VGND VPWR VPWR _4208_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2767 _4214_/X VGND VGND VPWR VPWR hold784/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5188_ _5203_/C _5183_/C _5038_/B VGND VGND VPWR VPWR _5188_/X sky130_fd_sc_hd__o21a_2
Xhold2778 _4356_/X VGND VGND VPWR VPWR hold852/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2789 hold969/X VGND VGND VPWR VPWR _4453_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4139_ _7269_/Q input89/X _4142_/A VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__mux2_2
XFILLER_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4394__A _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout651_A _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6603__B2 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3968__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6367__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4569__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input45_A mgmt_gpio_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6784__A _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3959__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4081__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4243__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4908__A1 wire649/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _7582_/Q _3501_/X _3503_/X input33/X _3509_/X VGND VGND VPWR VPWR _3524_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_128_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4490_ _4544_/A1 _4490_/A1 _4490_/S VGND VGND VPWR VPWR _4490_/X sky130_fd_sc_hd__mux2_1
Xhold607 hold607/A VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6125__A3 _6086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold618 _4436_/X VGND VGND VPWR VPWR _7089_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3441_ _7314_/Q VGND VGND VPWR VPWR _3441_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6530__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ _7297_/Q _6074_/X _6079_/X _7329_/Q _6159_/X VGND VGND VPWR VPWR _6160_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5111_ _5111_/A _5111_/B _5111_/C VGND VGND VPWR VPWR _5111_/Y sky130_fd_sc_hd__nor3_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2008 hold495/X VGND VGND VPWR VPWR _5859_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6119_/A _6119_/B _6121_/A VGND VGND VPWR VPWR _6091_/X sky130_fd_sc_hd__and3_4
Xhold2019 hold459/X VGND VGND VPWR VPWR _4451_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5802__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1307 hold3256/X VGND VGND VPWR VPWR hold3257/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_4_6__f_wb_clk_i clkbuf_3_3_0_wb_clk_i/X VGND VGND VPWR VPWR _7627_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1318 _5644_/X VGND VGND VPWR VPWR _7265_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5042_ _5042_/A _5042_/B VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__nor2_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 hold3211/X VGND VGND VPWR VPWR hold3212/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4418__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6993_ _6999_/CLK _6993_/D VGND VGND VPWR VPWR _6993_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_51_csclk _7399_/CLK VGND VGND VPWR VPWR _7581_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold2783_A _7120_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5944_ _5944_/A0 _5998_/A1 _5946_/S VGND VGND VPWR VPWR _5944_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5875_ hold32/X _5947_/A _5893_/B VGND VGND VPWR VPWR _5883_/S sky130_fd_sc_hd__and3_4
XFILLER_179_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3558__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4153__S _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7614_ _7627_/CLK _7614_/D fanout691/X VGND VGND VPWR VPWR _7614_/Q sky130_fd_sc_hd__dfrtp_1
X_4826_ _5115_/A _5115_/B VGND VGND VPWR VPWR _4826_/Y sky130_fd_sc_hd__nand2_8
X_7545_ _7573_/CLK _7545_/D fanout736/X VGND VGND VPWR VPWR _7545_/Q sky130_fd_sc_hd__dfrtp_4
X_4757_ _4692_/Y _4730_/Y _4741_/Y _4755_/Y VGND VGND VPWR VPWR _4760_/C sky130_fd_sc_hd__o22a_1
XFILLER_119_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3583__B1 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3708_ input7/X _3872_/A2 _3485_/X _3532_/X input56/X VGND VGND VPWR VPWR _3708_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7476_ _7542_/CLK _7476_/D fanout720/X VGND VGND VPWR VPWR _7476_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4688_ _4088_/Y _4558_/X _4591_/Y VGND VGND VPWR VPWR _5328_/B sky130_fd_sc_hd__o21a_4
X_6427_ _6427_/A _6455_/B _6467_/A VGND VGND VPWR VPWR _6427_/X sky130_fd_sc_hd__and3_4
XANTENNA__6521__B1 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3639_ _7580_/Q _3501_/X _5643_/A _7673_/A _3638_/X VGND VGND VPWR VPWR _3642_/C
+ sky130_fd_sc_hd__a221o_4
XFILLER_150_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6358_ _7200_/Q _6317_/B _6079_/X _6120_/X _7019_/Q VGND VGND VPWR VPWR _6358_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3210 _4401_/X VGND VGND VPWR VPWR hold3210/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3886__A1 _7480_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3221 _7021_/Q VGND VGND VPWR VPWR hold3221/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3232 _4540_/X VGND VGND VPWR VPWR hold3232/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3886__B2 _7198_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5309_ _4698_/Y _4755_/Y _4777_/X _4692_/Y _5150_/C VGND VGND VPWR VPWR _5311_/B
+ sky130_fd_sc_hd__o221a_1
Xhold3243 hold3243/A VGND VGND VPWR VPWR _5804_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3254 hold3254/A VGND VGND VPWR VPWR _5604_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6289_ _7041_/Q _6089_/X _6285_/X _6286_/X _6288_/X VGND VGND VPWR VPWR _6289_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold2520 hold488/X VGND VGND VPWR VPWR _7287_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5712__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3265 hold3265/A VGND VGND VPWR VPWR hold3265/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3276 _7108_/Q VGND VGND VPWR VPWR _7105_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2531 _7124_/Q VGND VGND VPWR VPWR hold887/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3287 _7610_/Q VGND VGND VPWR VPWR _6330_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2542 _7563_/Q VGND VGND VPWR VPWR hold609/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3298 _7612_/Q VGND VGND VPWR VPWR _6355_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2553 _7477_/Q VGND VGND VPWR VPWR hold835/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2564 _7396_/Q VGND VGND VPWR VPWR hold975/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3638__B2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2575 hold737/X VGND VGND VPWR VPWR _4484_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1830 _4549_/X VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2586 hold847/X VGND VGND VPWR VPWR _5810_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1841 hold236/X VGND VGND VPWR VPWR _4398_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2597 _7119_/Q VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1852 hold357/X VGND VGND VPWR VPWR _5742_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1863 hold204/X VGND VGND VPWR VPWR _5907_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6109__A _7591_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1874 _7190_/Q VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5013__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1885 _5672_/X VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1896 hold457/X VGND VGND VPWR VPWR _5787_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_19_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7519_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6588__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6052__A2 _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1883_A _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6760__B1 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3574__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6107__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5315__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6512__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3877__A1 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3877__B2 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__D _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6815__A1 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3650__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4238__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6291__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6579__B1 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3990_ input11/X _3490_/X _5686_/A _7303_/Q _3989_/X VGND VGND VPWR VPWR _3990_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_90_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3801__A1 _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5660_ _5660_/A0 hold487/X _5667_/S VGND VGND VPWR VPWR _5660_/X sky130_fd_sc_hd__mux2_1
X_4611_ _4814_/C _4899_/A2 _4909_/D VGND VGND VPWR VPWR _4657_/C sky130_fd_sc_hd__o21bai_4
XFILLER_176_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5591_ _5591_/A0 _5732_/A1 _5595_/S VGND VGND VPWR VPWR _5591_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7330_ _7330_/CLK _7330_/D fanout711/X VGND VGND VPWR VPWR _7330_/Q sky130_fd_sc_hd__dfrtp_4
X_4542_ _4542_/A0 _4548_/A0 _4544_/S VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold404 hold404/A VGND VGND VPWR VPWR _7169_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7261_ _7525_/CLK _7261_/D fanout745/X VGND VGND VPWR VPWR _7261_/Q sky130_fd_sc_hd__dfrtp_4
Xhold426 hold426/A VGND VGND VPWR VPWR _7344_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6503__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4473_ _4473_/A _5619_/B _4533_/B VGND VGND VPWR VPWR _4478_/S sky130_fd_sc_hd__and3_2
Xhold437 hold437/A VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold448 _5841_/X VGND VGND VPWR VPWR _7440_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2531_A _7124_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6212_ _6212_/A _6212_/B _6212_/C VGND VGND VPWR VPWR _6212_/Y sky130_fd_sc_hd__nor3_4
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3424_ _7450_/Q VGND VGND VPWR VPWR _3424_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3544__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7192_ _7210_/CLK _7192_/D fanout700/X VGND VGND VPWR VPWR _7192_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_171_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6119_/D _6138_/X _6140_/X _6142_/X VGND VGND VPWR VPWR _6143_/X sky130_fd_sc_hd__a211o_2
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6806__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1104 hold2984/X VGND VGND VPWR VPWR hold2985/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _7588_/Q _6121_/B _7589_/Q VGND VGND VPWR VPWR _6074_/X sky130_fd_sc_hd__and3b_4
XFILLER_58_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3883__A4 _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_736 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1115 hold3054/X VGND VGND VPWR VPWR hold1115/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 hold3110/X VGND VGND VPWR VPWR _7112_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1137 hold3162/X VGND VGND VPWR VPWR hold3163/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6282__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5025_ _5025_/A _5185_/B _5025_/C _5025_/D VGND VGND VPWR VPWR _5026_/C sky130_fd_sc_hd__nand4_2
XFILLER_100_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1148 hold1148/A VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold1159 _5822_/X VGND VGND VPWR VPWR _7423_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6976_ _7633_/CLK _6976_/D VGND VGND VPWR VPWR _6976_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5388__A4 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5927_ _5990_/A1 _5927_/A1 _5928_/S VGND VGND VPWR VPWR _5927_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5793__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5858_ _5993_/A1 _5858_/A1 _5865_/S VGND VGND VPWR VPWR _5858_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6337__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4809_ _4809_/A _4809_/B _4809_/C VGND VGND VPWR VPWR _4812_/A sky130_fd_sc_hd__nor3_1
XANTENNA__6742__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5789_ _5789_/A0 _5996_/A1 hold48/X VGND VGND VPWR VPWR _5789_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5707__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7528_ _7528_/CLK _7528_/D fanout730/X VGND VGND VPWR VPWR _7528_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7459_ _7475_/CLK _7459_/D fanout729/X VGND VGND VPWR VPWR _7459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold960 hold960/A VGND VGND VPWR VPWR _7180_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold971 hold971/A VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold982 hold982/A VGND VGND VPWR VPWR _7433_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold993 hold993/A VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3040 hold3040/A VGND VGND VPWR VPWR _7575_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_135_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3051 _7093_/Q VGND VGND VPWR VPWR hold3051/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3062 _5613_/X VGND VGND VPWR VPWR hold3062/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3073 hold3073/A VGND VGND VPWR VPWR _4335_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input147_A wb_dat_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3084 _5939_/X VGND VGND VPWR VPWR hold3084/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3095 _7263_/Q VGND VGND VPWR VPWR hold3095/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2350 _7040_/Q VGND VGND VPWR VPWR hold677/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2361 _7541_/Q VGND VGND VPWR VPWR hold769/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_95_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2372 _7213_/Q VGND VGND VPWR VPWR hold653/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2383 hold549/X VGND VGND VPWR VPWR _5970_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4284__A1 _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2394 hold583/X VGND VGND VPWR VPWR _5763_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1660 hold194/X VGND VGND VPWR VPWR _5797_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1671 hold209/X VGND VGND VPWR VPWR _7465_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1682 hold74/X VGND VGND VPWR VPWR _3468_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1693 _7481_/Q VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6025__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4582__A _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5536__A1 _4997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3547__B1 _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6500__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3661__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6264__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4275__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6830_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6830_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_53_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6567__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6761_ _7191_/Q _6446_/X _6452_/X _7025_/Q _6760_/X VGND VGND VPWR VPWR _6761_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5775__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3973_ _7535_/Q _5947_/A _4539_/C _3972_/X VGND VGND VPWR VPWR _3973_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4642__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5712_ _6000_/A1 _5712_/A1 _5712_/S VGND VGND VPWR VPWR _5712_/X sky130_fd_sc_hd__mux2_1
X_6692_ _7123_/Q _6420_/C _6419_/A _7158_/Q _6691_/X VGND VGND VPWR VPWR _6697_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_188_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _5643_/A _5992_/D VGND VGND VPWR VPWR _5649_/S sky130_fd_sc_hd__nand2_8
XFILLER_191_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5574_ _5574_/A _5574_/B VGND VGND VPWR VPWR _5575_/C sky130_fd_sc_hd__and2_1
XFILLER_117_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7313_ _7581_/CLK _7313_/D fanout715/X VGND VGND VPWR VPWR _7313_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3555__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold201 hold201/A VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4525_ _4525_/A0 _5585_/A0 _4526_/S VGND VGND VPWR VPWR _4525_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold212 hold212/A VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold223 hold223/A VGND VGND VPWR VPWR _7500_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold234 hold234/A VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7244_ _7330_/CLK _7244_/D fanout711/X VGND VGND VPWR VPWR _7244_/Q sky130_fd_sc_hd__dfrtp_4
Xhold245 hold245/A VGND VGND VPWR VPWR _7358_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4456_ _4456_/A0 _5876_/A1 _4460_/S VGND VGND VPWR VPWR _4456_/X sky130_fd_sc_hd__mux2_1
Xhold256 hold256/A VGND VGND VPWR VPWR _7564_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold267 hold267/A VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold278 hold278/A VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3407_ _6932_/Q VGND VGND VPWR VPWR _6065_/C sky130_fd_sc_hd__inv_2
Xfanout703 fanout706/X VGND VGND VPWR VPWR fanout703/X sky130_fd_sc_hd__buf_6
Xhold289 hold289/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout714 fanout720/X VGND VGND VPWR VPWR fanout714/X sky130_fd_sc_hd__buf_4
XANTENNA__4667__A _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7175_ _7176_/CLK _7175_/D fanout722/X VGND VGND VPWR VPWR _7175_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4387_ _5817_/A1 _4387_/A1 _4387_/S VGND VGND VPWR VPWR _4387_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout725 _6839_/A VGND VGND VPWR VPWR fanout725/X sky130_fd_sc_hd__buf_8
Xfanout736 fanout750/X VGND VGND VPWR VPWR fanout736/X sky130_fd_sc_hd__buf_8
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _7528_/Q _6092_/X _6112_/X _7480_/Q _6125_/X VGND VGND VPWR VPWR _6126_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3710__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout747 fanout749/X VGND VGND VPWR VPWR fanout747/X sky130_fd_sc_hd__buf_6
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout758 _4831_/C VGND VGND VPWR VPWR _4984_/B sky130_fd_sc_hd__clkbuf_16
Xfanout769 _4844_/B VGND VGND VPWR VPWR _5282_/A sky130_fd_sc_hd__buf_8
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6255__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6057_ _7594_/Q _6429_/C _6466_/D VGND VGND VPWR VPWR _6747_/B sky130_fd_sc_hd__and3_4
XTAP_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout564_A _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5008_ _5113_/A _5180_/B _5049_/C _5059_/A VGND VGND VPWR VPWR _5008_/X sky130_fd_sc_hd__o31a_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6558__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4833__C _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold142_A _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ _7238_/CLK _6959_/D fanout691/X VGND VGND VPWR VPWR _6959_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6106__B _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_789 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_772 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4577__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold790 hold790/A VGND VGND VPWR VPWR _7404_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3481__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3701__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2180 _4415_/X VGND VGND VPWR VPWR hold510/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5900__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4257__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2191 hold585/X VGND VGND VPWR VPWR _5905_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1490 _5945_/X VGND VGND VPWR VPWR hold107/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5757__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_0__f_mgmt_gpio_in[4] clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR VPWR _4127_/A1
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_842 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5509__A1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3783__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6706__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6721__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput306 _4174_/X VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
Xoutput317 hold1068/X VGND VGND VPWR VPWR hold1069/A sky130_fd_sc_hd__buf_6
X_4310_ _4321_/S _4310_/B VGND VGND VPWR VPWR _4310_/Y sky130_fd_sc_hd__nand2_1
Xoutput328 hold1123/X VGND VGND VPWR VPWR hold1124/A sky130_fd_sc_hd__buf_6
XANTENNA_hold2062_A _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3940__B1 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput339 hold1066/X VGND VGND VPWR VPWR hold1067/A sky130_fd_sc_hd__buf_6
X_5290_ _5252_/Y _5461_/B _4854_/X VGND VGND VPWR VPWR _5290_/X sky130_fd_sc_hd__a21bo_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5590__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4241_ _4241_/A0 _4240_/X _4249_/S VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6485__A2 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5693__A0 _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4496__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4918__C _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4172_ _4178_/A _4427_/C VGND VGND VPWR VPWR _7103_/D sky130_fd_sc_hd__and2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4248__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5810__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5996__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2696_A _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5749__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6813_ _6812_/X _6813_/A1 _6822_/S VGND VGND VPWR VPWR _7641_/D sky130_fd_sc_hd__mux2_1
XFILLER_169_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5748__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5212__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6744_ _7200_/Q _4101_/X _6771_/A3 _6419_/C _7140_/Q VGND VGND VPWR VPWR _6744_/X
+ sky130_fd_sc_hd__a32o_1
X_3956_ input98/X _5785_/B _4265_/B _4370_/A _7041_/Q VGND VGND VPWR VPWR _3956_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4420__A1 _4447_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6675_ _6751_/S _7622_/Q _6673_/X _6674_/X VGND VGND VPWR VPWR _6675_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3774__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3887_ _7133_/Q _3670_/X _4497_/A _7153_/Q _3886_/X VGND VGND VPWR VPWR _3887_/X
+ sky130_fd_sc_hd__a221o_1
X_5626_ _5626_/A0 _5815_/A1 _5629_/S VGND VGND VPWR VPWR _5626_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6173__A1 _7410_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5557_ _5543_/X _5548_/Y _5556_/Y VGND VGND VPWR VPWR _5557_/X sky130_fd_sc_hd__a21o_1
X_4508_ _4508_/A0 _4544_/A1 _4508_/S VGND VGND VPWR VPWR _4508_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5488_ _5488_/A _5488_/B _5488_/C VGND VGND VPWR VPWR _5488_/Y sky130_fd_sc_hd__nand3_1
XFILLER_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6476__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4439_ _4439_/A0 _5991_/A1 _4439_/S VGND VGND VPWR VPWR _4439_/X sky130_fd_sc_hd__mux2_1
X_7227_ _7232_/CLK _7227_/D fanout689/X VGND VGND VPWR VPWR _7227_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout500 _6035_/Y VGND VGND VPWR VPWR _6136_/C sky130_fd_sc_hd__buf_6
XFILLER_132_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout511 _4857_/X VGND VGND VPWR VPWR _4939_/C sky130_fd_sc_hd__clkbuf_4
Xfanout522 _4709_/Y VGND VGND VPWR VPWR _5480_/B2 sky130_fd_sc_hd__buf_8
Xfanout533 _4585_/A VGND VGND VPWR VPWR _4675_/B sky130_fd_sc_hd__buf_12
XANTENNA_hold1427_A hold16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7158_ _7268_/CLK _7158_/D _6861_/A VGND VGND VPWR VPWR _7158_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout544 _4447_/A1 VGND VGND VPWR VPWR _5972_/A1 sky130_fd_sc_hd__buf_6
XFILLER_58_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout555 _5826_/A1 VGND VGND VPWR VPWR _5853_/A0 sky130_fd_sc_hd__buf_6
XFILLER_59_745 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout566 _5726_/A1 VGND VGND VPWR VPWR _5996_/A1 sky130_fd_sc_hd__buf_6
Xfanout577 hold1567/X VGND VGND VPWR VPWR _5949_/A1 sky130_fd_sc_hd__buf_6
XANTENNA__6228__A2 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6109_ _7591_/Q _7590_/Q _6144_/A _6144_/C VGND VGND VPWR VPWR _6109_/X sky130_fd_sc_hd__and4_1
Xfanout588 hold487/X VGND VGND VPWR VPWR _5912_/A1 sky130_fd_sc_hd__buf_4
XFILLER_100_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7089_ _7514_/CLK _7089_/D fanout744/X VGND VGND VPWR VPWR _7668_/A sky130_fd_sc_hd__dfrtp_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout599 hold26/X VGND VGND VPWR VPWR _5992_/D sky130_fd_sc_hd__buf_12
XFILLER_46_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5987__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4844__B _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5659__C _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4860__A _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3765__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6164__B2 _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6703__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input75_A porb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5675__A0 _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4478__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4246__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5442__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4473__C _4533_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5866__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _7553_/Q _3508_/X _3800_/X _3802_/X _3809_/X VGND VGND VPWR VPWR _3810_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_82_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4790_ _5107_/C _4807_/B _4790_/C VGND VGND VPWR VPWR _4791_/A sky130_fd_sc_hd__and3_1
XANTENNA__4402__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _6447_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_29 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ _7120_/Q _4455_/A _3637_/C _4455_/C _3740_/X VGND VGND VPWR VPWR _3741_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_119_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4920__D _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6460_ _6466_/A _6466_/B _6467_/A _6651_/B VGND VGND VPWR VPWR _6460_/X sky130_fd_sc_hd__and4_4
X_3672_ _4473_/A _5938_/B _4455_/C VGND VGND VPWR VPWR _4497_/A sky130_fd_sc_hd__and3_4
XFILLER_173_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5411_ _5408_/Y _4769_/Y _5145_/A _5306_/B VGND VGND VPWR VPWR _5568_/A sky130_fd_sc_hd__o211a_1
X_6391_ _7070_/Q _6317_/B _6332_/C _6075_/X _7166_/Q VGND VGND VPWR VPWR _6391_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5805__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5342_ _5342_/A _5342_/B _5342_/C VGND VGND VPWR VPWR _5343_/A sky130_fd_sc_hd__and3_2
XFILLER_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4929__B _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6458__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5273_ _5561_/A1 _5480_/B2 _4806_/Y _5516_/A3 _4798_/Y VGND VGND VPWR VPWR _5476_/A
+ sky130_fd_sc_hd__o32a_1
Xhold2905 _5621_/X VGND VGND VPWR VPWR hold2905/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_7012_ _7181_/CLK _7012_/D fanout721/X VGND VGND VPWR VPWR _7012_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3552__C _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2916 _7008_/Q VGND VGND VPWR VPWR hold2916/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4224_ _4224_/A0 _4223_/X _4232_/S VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__mux2_1
Xhold2927 hold2927/A VGND VGND VPWR VPWR _4306_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_99_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2938 hold2938/A VGND VGND VPWR VPWR _4343_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2949 hold2949/A VGND VGND VPWR VPWR _4512_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4155_ _4154_/X _4135_/B _6896_/Q VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__mux2_2
XANTENNA__3692__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ _4825_/A _4674_/A VGND VGND VPWR VPWR _4086_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5969__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4156__S input1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6630__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5776__A _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4680__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5197__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4988_ _5339_/D _5183_/A _5203_/C _5339_/C VGND VGND VPWR VPWR _5041_/D sky130_fd_sc_hd__nand4_1
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6727_ _6726_/X _6751_/A1 _6777_/S VGND VGND VPWR VPWR _7625_/D sky130_fd_sc_hd__mux2_1
X_3939_ _7137_/Q _4479_/A _3576_/X _4467_/A _7127_/Q VGND VGND VPWR VPWR _3939_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6658_ _7026_/Q _6651_/B _6459_/C _6408_/B _7041_/Q VGND VGND VPWR VPWR _6658_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4157__B1 _7290_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5609_ _5609_/A0 _5627_/A1 _5611_/S VGND VGND VPWR VPWR _5609_/X sky130_fd_sc_hd__mux2_1
X_6589_ _7500_/Q _6600_/B _6651_/C _6468_/X _7412_/Q VGND VGND VPWR VPWR _6589_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6449__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5657__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1809_A _7520_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout363 hold1254/X VGND VGND VPWR VPWR _4527_/A sky130_fd_sc_hd__buf_8
Xfanout374 _5404_/A VGND VGND VPWR VPWR _5410_/A sky130_fd_sc_hd__buf_6
Xfanout385 _5659_/B VGND VGND VPWR VPWR _5640_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__3683__A2 _3848_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout396 _3848_/A2 VGND VGND VPWR VPWR _5965_/B sky130_fd_sc_hd__buf_8
XFILLER_100_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6621__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5686__A _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5188__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4396__A0 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__6137__A1 _7288_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_4
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_4
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6688__A2 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5896__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5360__A2 _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3653__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5648__A0 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_5__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X VGND VGND VPWR VPWR _7621_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5112__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4320__A0 _3607_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5960_ _5960_/A0 _5969_/A1 _5964_/S VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4911_ _5065_/A _4933_/A _4970_/C _4940_/D VGND VGND VPWR VPWR _4913_/B sky130_fd_sc_hd__nand4_2
X_5891_ _5891_/A0 _5990_/A1 hold91/X VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3977__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5596__A _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7630_ _7630_/CLK _7630_/D VGND VGND VPWR VPWR _7630_/Q sky130_fd_sc_hd__dfxtp_1
X_4842_ _4748_/A _5091_/A VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__4387__A0 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4773_ _5100_/A _4797_/B _5260_/C VGND VGND VPWR VPWR _5086_/B sky130_fd_sc_hd__and3_2
XANTENNA__3729__A3 _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7561_ _7561_/CLK _7561_/D fanout737/X VGND VGND VPWR VPWR _7561_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3724_ _6923_/Q _3542_/X _5704_/A _7323_/Q VGND VGND VPWR VPWR _3724_/X sky130_fd_sc_hd__a22o_1
X_6512_ _7513_/Q _6435_/X _6446_/X _7521_/Q VGND VGND VPWR VPWR _6512_/X sky130_fd_sc_hd__a22o_1
XFILLER_158_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7492_ _7579_/CLK _7492_/D fanout732/X VGND VGND VPWR VPWR _7492_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6679__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6443_ _6455_/B _6443_/B _6466_/D VGND VGND VPWR VPWR _6443_/X sky130_fd_sc_hd__and3_4
X_3655_ _7672_/A _5992_/A _3860_/D _4479_/A VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__and4_1
XFILLER_173_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6374_ _6877_/Q _6112_/X _6371_/X _6373_/X _6372_/X VGND VGND VPWR VPWR _6374_/X
+ sky130_fd_sc_hd__a2111o_1
X_3586_ _7357_/Q _3506_/X _5758_/A _7373_/Q _3585_/X VGND VGND VPWR VPWR _3587_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5351__A2 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4659__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3563__B _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5325_ _5295_/B _4977_/X _5046_/A _5007_/Y VGND VGND VPWR VPWR _5325_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3901__A3 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5639__A0 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5256_ _4601_/Y _4744_/Y _4716_/Y _5563_/A1 VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__a211o_1
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2702 _4386_/X VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2713 _7419_/Q VGND VGND VPWR VPWR hold787/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2724 _7125_/Q VGND VGND VPWR VPWR hold857/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2735 hold813/X VGND VGND VPWR VPWR _5772_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4207_ hold120/X _5625_/A1 _4207_/S VGND VGND VPWR VPWR _4207_/X sky130_fd_sc_hd__mux2_1
Xhold2746 _7236_/Q VGND VGND VPWR VPWR hold761/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_180_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2757 _4555_/X VGND VGND VPWR VPWR hold952/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5187_ _5178_/X _5038_/C _5186_/X _5185_/Y VGND VGND VPWR VPWR _5187_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6793__B1_N _7107_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2768 hold784/X VGND VGND VPWR VPWR _6928_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4862__A1 _4831_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2779 _7459_/Q VGND VGND VPWR VPWR hold815/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4138_ _7270_/Q input91/X _4142_/A VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__mux2_2
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6603__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4069_ hold18/A hold9/A _4074_/S VGND VGND VPWR VPWR _6889_/D sky130_fd_sc_hd__mux2_1
XFILLER_43_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5024__D1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3738__B _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5327__C1 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4550__A0 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__B _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4302__A0 _3570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input38_A mgmt_gpio_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5802__A0 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3959__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__A1 _7200_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3664__A _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold608 hold608/A VGND VGND VPWR VPWR _7278_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6040__A _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3440_ _7322_/Q VGND VGND VPWR VPWR _3440_/Y sky130_fd_sc_hd__inv_2
Xhold619 hold619/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6530__A1 _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5110_ _5282_/B _5453_/B _5282_/C VGND VGND VPWR VPWR _5110_/X sky130_fd_sc_hd__and3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6090_ _6119_/A _6119_/B _6097_/B _6144_/C VGND VGND VPWR VPWR _6090_/X sky130_fd_sc_hd__and4_4
Xhold2009 _5859_/X VGND VGND VPWR VPWR hold496/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__B1 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5041_/A _5041_/B _5041_/C _5041_/D VGND VGND VPWR VPWR _5042_/B sky130_fd_sc_hd__nand4_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1308 hold3258/X VGND VGND VPWR VPWR _7343_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1319 hold3174/X VGND VGND VPWR VPWR hold3175/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4645__D _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6992_ _7497_/CLK _6992_/D fanout693/X VGND VGND VPWR VPWR _6992_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__7532__RESET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5943_ _5943_/A0 _5979_/A0 _5946_/S VGND VGND VPWR VPWR _5943_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4942__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6349__B2 _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5874_ _5874_/A0 _5991_/A1 _5874_/S VGND VGND VPWR VPWR _5874_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3558__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7613_ _7627_/CLK _7613_/D fanout691/X VGND VGND VPWR VPWR _7613_/Q sky130_fd_sc_hd__dfrtp_1
X_4825_ _4825_/A _5071_/B _5071_/C _5089_/B VGND VGND VPWR VPWR _4825_/Y sky130_fd_sc_hd__nor4_1
XFILLER_166_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7544_ _7556_/CLK _7544_/D fanout732/X VGND VGND VPWR VPWR _7544_/Q sky130_fd_sc_hd__dfstp_2
X_4756_ _4823_/D _5134_/A _5068_/B VGND VGND VPWR VPWR _4756_/X sky130_fd_sc_hd__and3_1
XANTENNA__3583__A1 _7525_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3707_ _7547_/Q _5965_/A _5956_/B _3508_/X _7555_/Q VGND VGND VPWR VPWR _3707_/X
+ sky130_fd_sc_hd__a32o_1
X_4687_ _5138_/B _4687_/B _4687_/C VGND VGND VPWR VPWR _4687_/Y sky130_fd_sc_hd__nand3_4
X_7475_ _7475_/CLK _7475_/D fanout730/X VGND VGND VPWR VPWR _7475_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6426_ _6441_/D _6466_/B _6467_/A VGND VGND VPWR VPWR _6426_/X sky130_fd_sc_hd__and3_4
X_3638_ _7572_/Q _5983_/A _3637_/C _7452_/Q _5848_/A VGND VGND VPWR VPWR _3638_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6521__B2 _7281_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3200 _4266_/X VGND VGND VPWR VPWR hold3200/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3569_ _3682_/A _5947_/B _4509_/C VGND VGND VPWR VPWR _5893_/A sky130_fd_sc_hd__and3_4
X_6357_ _7059_/Q _6085_/X _6119_/X _7135_/Q _6356_/X VGND VGND VPWR VPWR _6357_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout594_A _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3211 _7036_/Q VGND VGND VPWR VPWR hold3211/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3886__A2 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3222 hold3222/A VGND VGND VPWR VPWR _4347_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3233 _7229_/Q VGND VGND VPWR VPWR hold3233/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_115_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5308_ _5308_/A _5308_/B _5308_/C VGND VGND VPWR VPWR _5311_/A sky130_fd_sc_hd__nor3_1
Xhold3244 _5804_/X VGND VGND VPWR VPWR hold3244/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6288_ _7112_/Q _6317_/C _6074_/X _6967_/Q _6287_/X VGND VGND VPWR VPWR _6288_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5088__A1 _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2510 _7201_/Q VGND VGND VPWR VPWR hold683/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3255 _5604_/X VGND VGND VPWR VPWR hold3255/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2521 _7324_/Q VGND VGND VPWR VPWR hold941/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3266 _7399_/Q VGND VGND VPWR VPWR hold3266/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3277 _7103_/Q VGND VGND VPWR VPWR _4425_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2532 hold887/X VGND VGND VPWR VPWR _4464_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3288 _6307_/X VGND VGND VPWR VPWR _7610_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5239_ _5222_/A _5453_/A _5453_/B _4934_/B _5237_/Y VGND VGND VPWR VPWR _5239_/X
+ sky130_fd_sc_hd__a311o_1
Xhold2543 hold609/X VGND VGND VPWR VPWR _5979_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3299 _7643_/Q VGND VGND VPWR VPWR _6819_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2554 hold835/X VGND VGND VPWR VPWR _5882_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2565 hold975/X VGND VGND VPWR VPWR _5791_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1820 hold257/X VGND VGND VPWR VPWR _4392_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3638__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4835__A1 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1831 _7344_/Q VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4835__B2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2576 _4484_/X VGND VGND VPWR VPWR hold738/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2587 _5810_/X VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1842 _4398_/X VGND VGND VPWR VPWR hold237/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2598 hold845/X VGND VGND VPWR VPWR _4458_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1853 _5742_/X VGND VGND VPWR VPWR hold358/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1864 _5907_/X VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6109__B _7590_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1875 hold253/X VGND VGND VPWR VPWR _4543_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1886 _7170_/Q VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1897 _7504_/Q VGND VGND VPWR VPWR hold437/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3810__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5563__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3574__B2 _7565_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6512__A1 _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6512__B2 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5903__S hold42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3877__A2 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3931__B _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__buf_8
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output311_A _7628_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6579__B2 _7532_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3659__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3801__A2 _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6200__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _5100_/A _4645_/D VGND VGND VPWR VPWR _4657_/D sky130_fd_sc_hd__nand2_2
XFILLER_175_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5590_ _5590_/A _5596_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5590_/X sky130_fd_sc_hd__and4_4
XFILLER_90_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4541_ _4541_/A0 hold198/X _4544_/S VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold416 hold416/A VGND VGND VPWR VPWR _7512_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4472_ _5853_/A0 _4472_/A1 _4472_/S VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__mux2_1
X_7260_ _7578_/CLK _7260_/D fanout747/X VGND VGND VPWR VPWR _7260_/Q sky130_fd_sc_hd__dfrtp_4
Xhold427 hold427/A VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6503__B2 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold438 hold438/A VGND VGND VPWR VPWR _7504_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3423_ _7458_/Q VGND VGND VPWR VPWR _3423_/Y sky130_fd_sc_hd__inv_2
Xhold449 hold449/A VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6211_ _6110_/A _6202_/X _6207_/X _6210_/X VGND VGND VPWR VPWR _6212_/C sky130_fd_sc_hd__a211o_1
XFILLER_143_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7191_ _7191_/CLK _7191_/D _6872_/A VGND VGND VPWR VPWR _7191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5813__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3868__A2 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6142_ _7456_/Q _6080_/X _6090_/X _7376_/Q _6141_/X VGND VGND VPWR VPWR _6142_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6267__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6099_/D _6081_/C _6112_/B VGND VGND VPWR VPWR _6073_/X sky130_fd_sc_hd__and3_2
XFILLER_85_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1105 hold3059/X VGND VGND VPWR VPWR hold1105/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 hold1116/A VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
Xhold1127 hold3130/X VGND VGND VPWR VPWR hold3131/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5024_ _5024_/A1 _4669_/X _4974_/B _5180_/A _5038_/A VGND VGND VPWR VPWR _5185_/B
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_57_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1138 hold3164/X VGND VGND VPWR VPWR _7415_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1149 hold2942/X VGND VGND VPWR VPWR hold2943/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5490__A1 _4997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6416__B_N _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6975_ _7636_/CLK _6975_/D VGND VGND VPWR VPWR _6975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5242__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3569__A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4164__S _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5926_ _5980_/A0 _5926_/A1 _5928_/S VGND VGND VPWR VPWR _5926_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5857_ _5857_/A _5893_/B VGND VGND VPWR VPWR _5865_/S sky130_fd_sc_hd__nand2_8
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4808_ _5410_/A _5061_/B _5453_/B VGND VGND VPWR VPWR _4809_/B sky130_fd_sc_hd__and3_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout607_A _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5788_ _5788_/A0 _5788_/A1 hold48/X VGND VGND VPWR VPWR _5788_/X sky130_fd_sc_hd__mux2_1
X_7527_ _7574_/CLK _7527_/D fanout739/X VGND VGND VPWR VPWR _7527_/Q sky130_fd_sc_hd__dfstp_4
X_4739_ _4730_/Y _4732_/Y _4738_/X VGND VGND VPWR VPWR _5139_/D sky130_fd_sc_hd__o21a_1
X_7458_ _7574_/CLK _7458_/D fanout745/X VGND VGND VPWR VPWR _7458_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6111__C _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6409_ _6441_/D _6433_/D _6434_/B _6462_/C VGND VGND VPWR VPWR _6409_/X sky130_fd_sc_hd__and4_4
Xhold950 _5773_/X VGND VGND VPWR VPWR _7380_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold961 hold961/A VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7389_ _7582_/CLK _7389_/D fanout716/X VGND VGND VPWR VPWR _7389_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold972 _4495_/X VGND VGND VPWR VPWR _7150_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5723__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap680 _5089_/C VGND VGND VPWR VPWR _4833_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold983 hold983/A VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold994 _4537_/X VGND VGND VPWR VPWR _7185_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3030 _6977_/Q VGND VGND VPWR VPWR _4287_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3041 _7450_/Q VGND VGND VPWR VPWR hold3041/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3052 hold3052/A VGND VGND VPWR VPWR _4441_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3063 _7629_/Q VGND VGND VPWR VPWR _6781_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3074 _4335_/X VGND VGND VPWR VPWR hold3074/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2340 _4393_/X VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3085 _7351_/Q VGND VGND VPWR VPWR hold3085/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3096 hold3096/A VGND VGND VPWR VPWR _5641_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2351 hold677/X VGND VGND VPWR VPWR _4369_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2362 hold769/X VGND VGND VPWR VPWR _5954_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2373 hold653/X VGND VGND VPWR VPWR _5586_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2384 _7571_/Q VGND VGND VPWR VPWR hold547/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1650 hold133/X VGND VGND VPWR VPWR _7232_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4284__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2395 _5763_/X VGND VGND VPWR VPWR hold584/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1661 _5797_/X VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1672 _7525_/Q VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1683 _3467_/Y VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1694 hold210/X VGND VGND VPWR VPWR _5887_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4582__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5233__B2 _4790_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5536__A2 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3547__A1 _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3547__B2 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_csclk _7399_/CLK VGND VGND VPWR VPWR _7576_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6249__B1 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3661__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4249__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk _7399_/CLK VGND VGND VPWR VPWR _7489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4773__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4923__D _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6760_ _7060_/Q _6447_/C _6651_/C _6419_/A _7161_/Q VGND VGND VPWR VPWR _6760_/X
+ sky130_fd_sc_hd__a32o_1
X_3972_ _7177_/Q _4539_/C _5619_/B _3647_/X _7167_/Q VGND VGND VPWR VPWR _3972_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5711_ _5972_/A1 _5711_/A1 _5712_/S VGND VGND VPWR VPWR _5711_/X sky130_fd_sc_hd__mux2_1
X_6691_ _7002_/Q _6419_/D _6421_/X _7007_/Q VGND VGND VPWR VPWR _6691_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5808__S _5811_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5642_ _5642_/A0 _5645_/A0 _5642_/S VGND VGND VPWR VPWR _5642_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5573_ _5231_/B _5573_/B _5573_/C _5573_/D VGND VGND VPWR VPWR _5574_/B sky130_fd_sc_hd__and4b_1
XANTENNA_hold2641_A _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_780 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7312_ _7576_/CLK _7312_/D fanout717/X VGND VGND VPWR VPWR _7312_/Q sky130_fd_sc_hd__dfstp_2
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4524_ _4524_/A0 _5788_/A1 _4526_/S VGND VGND VPWR VPWR _4524_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3555__C _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold213 _5682_/X VGND VGND VPWR VPWR _7299_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_18_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7197_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6488__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold235 hold235/A VGND VGND VPWR VPWR _7176_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7243_ _7329_/CLK _7243_/D fanout704/X VGND VGND VPWR VPWR _7243_/Q sky130_fd_sc_hd__dfstp_4
Xhold246 _6903_/Q VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4455_ _4455_/A _4479_/A _4455_/C _4533_/B VGND VGND VPWR VPWR _4460_/S sky130_fd_sc_hd__and4_4
Xhold257 hold257/A VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold268 hold268/A VGND VGND VPWR VPWR _7069_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold279 hold279/A VGND VGND VPWR VPWR _7307_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3406_ _7585_/Q VGND VGND VPWR VPWR _4099_/D sky130_fd_sc_hd__inv_2
Xfanout704 fanout706/X VGND VGND VPWR VPWR fanout704/X sky130_fd_sc_hd__buf_8
X_4386_ _5585_/A0 _4386_/A1 _4387_/S VGND VGND VPWR VPWR _4386_/X sky130_fd_sc_hd__mux2_1
X_7174_ _7176_/CLK _7174_/D fanout722/X VGND VGND VPWR VPWR _7174_/Q sky130_fd_sc_hd__dfstp_4
Xfanout715 fanout720/X VGND VGND VPWR VPWR fanout715/X sky130_fd_sc_hd__buf_8
Xfanout726 _6839_/A VGND VGND VPWR VPWR fanout726/X sky130_fd_sc_hd__buf_4
XFILLER_98_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout737 fanout740/X VGND VGND VPWR VPWR fanout737/X sky130_fd_sc_hd__buf_8
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _7464_/Q _6075_/A _6086_/X _6099_/X _7352_/Q VGND VGND VPWR VPWR _6125_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3710__B2 _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout748 fanout749/X VGND VGND VPWR VPWR fanout748/X sky130_fd_sc_hd__buf_8
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _4772_/A VGND VGND VPWR VPWR _4909_/D sky130_fd_sc_hd__clkbuf_16
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _7598_/Q _7597_/Q VGND VGND VPWR VPWR _6056_/X sky130_fd_sc_hd__and2b_1
XTAP_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5007_ _5059_/A _5180_/B VGND VGND VPWR VPWR _5007_/Y sky130_fd_sc_hd__nand2_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout557_A _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ _7238_/CLK _6958_/D fanout690/X VGND VGND VPWR VPWR _6958_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout724_A fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6106__C _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5909_ _5954_/A1 _5909_/A1 hold42/A VGND VGND VPWR VPWR _5909_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3777__B2 _7227_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6889_ _4169_/B2 _6889_/D _6839_/X VGND VGND VPWR VPWR _6889_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold1574_A _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6403__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6715__A1 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5151__B1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold780 _5629_/X VGND VGND VPWR VPWR _7255_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3481__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3122_A _6874_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6246__A3 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2170 _4237_/X VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5454__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input20_A mask_rev_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2181 _6925_/Q VGND VGND VPWR VPWR hold561/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2192 _5905_/X VGND VGND VPWR VPWR hold586/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6284__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1480 _7453_/Q VGND VGND VPWR VPWR hold64/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1491 _6889_/Q VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3768__A1 _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6706__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3656__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4193__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput307 _4134_/X VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
Xoutput318 hold1070/X VGND VGND VPWR VPWR hold1071/A sky130_fd_sc_hd__buf_6
Xoutput329 hold1105/X VGND VGND VPWR VPWR hold1106/A sky130_fd_sc_hd__buf_6
XFILLER_114_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _5654_/A1 _5951_/A1 _4248_/S VGND VGND VPWR VPWR _4240_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4171_ _4178_/A _4171_/B VGND VGND VPWR VPWR _7104_/D sky130_fd_sc_hd__and2_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5445__A1 _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6642__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6812_ _4427_/B _6812_/A2 _6812_/B1 wire536/A _6811_/X VGND VGND VPWR VPWR _6812_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6743_ _7170_/Q _6408_/D _6421_/X _7009_/Q _6742_/X VGND VGND VPWR VPWR _6749_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3955_ _7527_/Q _3529_/X _5776_/A _7383_/Q VGND VGND VPWR VPWR _3955_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4442__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6674_ _6957_/Q _6431_/Y _6067_/A VGND VGND VPWR VPWR _6674_/X sky130_fd_sc_hd__o21a_1
X_3886_ _7480_/Q _3535_/X _3673_/X _7198_/Q _3885_/X VGND VGND VPWR VPWR _3886_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5625_ _5625_/A0 _5625_/A1 _5629_/S VGND VGND VPWR VPWR _5625_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4184__A1 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5556_ _5533_/Y _5539_/X _5555_/X VGND VGND VPWR VPWR _5556_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4507_ _4507_/A0 _5625_/A1 _4508_/S VGND VGND VPWR VPWR _4507_/X sky130_fd_sc_hd__mux2_1
X_5487_ _4801_/B _4801_/C _4768_/Y _5408_/Y _5153_/C VGND VGND VPWR VPWR _5488_/C
+ sky130_fd_sc_hd__o41a_1
X_7226_ _7232_/CLK _7226_/D _4128_/B VGND VGND VPWR VPWR _7226_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5133__B1 _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4438_ _4438_/A0 _5990_/A1 _4439_/S VGND VGND VPWR VPWR _4438_/X sky130_fd_sc_hd__mux2_1
Xfanout501 _6116_/C VGND VGND VPWR VPWR _6097_/B sky130_fd_sc_hd__buf_8
XANTENNA__5684__A1 _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout512 _4844_/Y VGND VGND VPWR VPWR _5509_/A3 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout523 _4811_/D VGND VGND VPWR VPWR _5113_/A sky130_fd_sc_hd__clkbuf_16
X_7157_ _7266_/CLK _7157_/D fanout694/X VGND VGND VPWR VPWR _7157_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout545 _4447_/A1 VGND VGND VPWR VPWR _5990_/A1 sky130_fd_sc_hd__buf_6
X_4369_ _4369_/A0 _5736_/A1 _4369_/S VGND VGND VPWR VPWR _4369_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout556 _5826_/A1 VGND VGND VPWR VPWR _5997_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout567 _5950_/A1 VGND VGND VPWR VPWR _5815_/A1 sky130_fd_sc_hd__buf_8
X_6108_ _6104_/X _6105_/X _6107_/X _6121_/C VGND VGND VPWR VPWR _6108_/X sky130_fd_sc_hd__o31a_1
XFILLER_100_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout578 hold1567/X VGND VGND VPWR VPWR _5994_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__4858__A_N _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7088_ _7514_/CLK _7088_/D fanout743/X VGND VGND VPWR VPWR _7667_/A sky130_fd_sc_hd__dfrtp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 hold487/X VGND VGND VPWR VPWR _5993_/A1 sky130_fd_sc_hd__buf_8
XFILLER_100_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6633__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6039_ _6121_/C _6038_/X _6037_/X VGND VGND VPWR VPWR _7592_/D sky130_fd_sc_hd__o21ai_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__B _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1956_A _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input68_A mgmt_gpio_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_4__f_wb_clk_i clkbuf_3_2_0_wb_clk_i/X VGND VGND VPWR VPWR _7625_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6219__A3 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3989__A1 input93/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_808 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5866__B _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4770__B _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3667__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_19 _6495_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _7570_/Q _5983_/A _3637_/C _5643_/A input64/X VGND VGND VPWR VPWR _3740_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3610__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3671_ _5992_/A _4455_/C _4265_/B VGND VGND VPWR VPWR _5634_/A sky130_fd_sc_hd__and3_4
X_5410_ _5410_/A _5410_/B _5410_/C VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__and3_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6390_ _7020_/Q _6120_/X _6386_/X _6387_/X _6389_/X VGND VGND VPWR VPWR _6397_/A
+ sky130_fd_sc_hd__a2111o_1
X_5341_ _5180_/B _5058_/C _5202_/B VGND VGND VPWR VPWR _5343_/B sky130_fd_sc_hd__a21bo_2
XANTENNA__4929__C _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6458__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5272_ _4709_/Y _4798_/Y _5516_/A3 _4789_/Y _5271_/X VGND VGND VPWR VPWR _5272_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5666__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7011_ _7211_/CLK _7011_/D fanout698/X VGND VGND VPWR VPWR _7011_/Q sky130_fd_sc_hd__dfrtp_4
Xhold2906 _5622_/X VGND VGND VPWR VPWR hold2906/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4223_ _4254_/A0 _5969_/A1 _4231_/S VGND VGND VPWR VPWR _4223_/X sky130_fd_sc_hd__mux2_1
Xhold2917 hold2917/A VGND VGND VPWR VPWR _4331_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2928 _4306_/X VGND VGND VPWR VPWR hold2928/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2939 _4343_/X VGND VGND VPWR VPWR hold2939/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_4154_ _4153_/X input38/X _6898_/Q VGND VGND VPWR VPWR _4154_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4945__B _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3692__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4085_ _6895_/Q _4085_/A2 _6839_/B VGND VGND VPWR VPWR _4178_/A sky130_fd_sc_hd__o21ai_2
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3466__B1_N _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4987_ _5339_/D _5183_/A _5029_/A _5339_/C VGND VGND VPWR VPWR _5041_/C sky130_fd_sc_hd__nand4_1
XANTENNA__6394__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__A _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6726_ _6725_/X _6726_/A1 _6751_/S VGND VGND VPWR VPWR _6726_/X sky130_fd_sc_hd__mux2_1
XFILLER_149_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3938_ _7243_/Q _5992_/A _3485_/X _3860_/D _3937_/X VGND VGND VPWR VPWR _3938_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_134_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6657_ _7132_/Q _6409_/X _6420_/B _6988_/Q _6655_/X VGND VGND VPWR VPWR _6657_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_149_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3869_ _7148_/Q _3652_/X _3654_/X _7118_/Q _3859_/X VGND VGND VPWR VPWR _3869_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4157__A1 _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5608_ _5608_/A0 _5736_/A1 _5611_/S VGND VGND VPWR VPWR _5608_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6588_ _7460_/Q _4101_/X _6574_/C _6463_/X _7428_/Q VGND VGND VPWR VPWR _6588_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ _5488_/Y _5539_/B _5568_/B VGND VGND VPWR VPWR _5539_/X sky130_fd_sc_hd__and3b_1
XFILLER_191_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7209_ _7210_/CLK _7209_/D fanout702/X VGND VGND VPWR VPWR _7209_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout364 _4376_/B VGND VGND VPWR VPWR _5938_/C sky130_fd_sc_hd__buf_8
XFILLER_143_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5409__A1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6606__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout386 _4265_/B VGND VGND VPWR VPWR _5659_/B sky130_fd_sc_hd__buf_12
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout397 hold1685/X VGND VGND VPWR VPWR _3848_/A2 sky130_fd_sc_hd__buf_8
XFILLER_100_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4574__C _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input122_A wb_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4632__A2 _4984_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5686__B _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5906__S hold42/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR _4177_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_128_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3653__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6612__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4084__B1 _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5820__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4910_ _4840_/D _5399_/A _4924_/B _4910_/D VGND VGND VPWR VPWR _4928_/B sky130_fd_sc_hd__and4b_2
XTAP_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5890_ _5890_/A0 _5980_/A0 hold91/X VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5596__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4841_ _4841_/A _4841_/B _4841_/C VGND VGND VPWR VPWR _4851_/A sky130_fd_sc_hd__nor3_1
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6376__A2 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5584__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7560_ _7563_/CLK _7560_/D fanout739/X VGND VGND VPWR VPWR _7560_/Q sky130_fd_sc_hd__dfstp_2
X_4772_ _4772_/A _4772_/B _4797_/B VGND VGND VPWR VPWR _4775_/C sky130_fd_sc_hd__and3_4
X_6511_ _7361_/Q _6462_/X _6502_/X _6506_/X _6510_/X VGND VGND VPWR VPWR _6511_/X
+ sky130_fd_sc_hd__a2111o_1
X_3723_ _6992_/Q _5731_/B _5623_/B _3531_/X _7339_/Q VGND VGND VPWR VPWR _3723_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6128__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7491_ _7491_/CLK _7491_/D fanout730/X VGND VGND VPWR VPWR _7491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_158_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5816__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4139__A1 input89/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6442_ _7495_/Q _6600_/B _6651_/C _6422_/X _7287_/Q VGND VGND VPWR VPWR _6442_/X
+ sky130_fd_sc_hd__a32o_1
X_3654_ _4455_/A _4479_/A _4455_/C VGND VGND VPWR VPWR _3654_/X sky130_fd_sc_hd__and3_2
XANTENNA__5887__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6373_ _7145_/Q _6082_/C _6097_/B _6144_/B VGND VGND VPWR VPWR _6373_/X sky130_fd_sc_hd__o211a_1
XFILLER_161_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_0_0_wb_clk_i clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR clkbuf_3_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_8
X_3585_ _7285_/Q _5731_/A _5659_/B _5857_/A _7461_/Q VGND VGND VPWR VPWR _3585_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3563__C _3563_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5324_ _5324_/A _5324_/B VGND VGND VPWR VPWR _5340_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2703 _7212_/Q VGND VGND VPWR VPWR hold843/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4956__A _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5255_ _4879_/D _4747_/B _5073_/B _4601_/Y VGND VGND VPWR VPWR _5255_/X sky130_fd_sc_hd__o31a_4
XANTENNA__6300__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2714 hold787/X VGND VGND VPWR VPWR _5817_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5103__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3860__A _7183_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2725 hold857/X VGND VGND VPWR VPWR _4465_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4206_ _4206_/A0 _5815_/A1 _4211_/S VGND VGND VPWR VPWR _4206_/X sky130_fd_sc_hd__mux2_1
Xhold2736 _7357_/Q VGND VGND VPWR VPWR hold927/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4311__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2747 hold761/X VGND VGND VPWR VPWR _5605_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2758 _7311_/Q VGND VGND VPWR VPWR hold541/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5186_ _5034_/B _5180_/B _5030_/C _5026_/A VGND VGND VPWR VPWR _5186_/X sky130_fd_sc_hd__a31o_1
Xhold2769 _7044_/Q VGND VGND VPWR VPWR hold953/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4167__S _7255_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4137_ _7073_/Q _4136_/Y _3996_/A VGND VGND VPWR VPWR _6881_/D sky130_fd_sc_hd__o21a_4
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6603__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4068_ _4098_/A1 _4062_/B _4062_/Y _4076_/B _4067_/Y VGND VGND VPWR VPWR _6890_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5811__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6897__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4691__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5024__C1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6367__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4378__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3738__C _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ _7134_/Q _6409_/X _6422_/X _6964_/Q _6708_/X VGND VGND VPWR VPWR _6709_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5726__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5878__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3889__B1 _5713_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4569__C _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3473__C _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4866__A _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__B1 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4369__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output291_A _6925_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3592__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5869__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3664__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6040__B _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6530__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4479__C _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4541__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_max_cap602_A _4075_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__B2 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5040_ _5158_/A _5339_/D _5183_/A _5339_/C VGND VGND VPWR VPWR _5041_/B sky130_fd_sc_hd__nand4_1
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 hold3240/X VGND VGND VPWR VPWR hold3241/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4926__D _5260_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ _6991_/CLK _6991_/D fanout693/X VGND VGND VPWR VPWR _6991_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__6597__A2 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5942_ _5942_/A0 _5978_/A0 _5946_/S VGND VGND VPWR VPWR _5942_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3804__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6349__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5873_ _5873_/A0 _5990_/A1 _5874_/S VGND VGND VPWR VPWR _5873_/X sky130_fd_sc_hd__mux2_1
X_7612_ _7627_/CLK _7612_/D fanout691/X VGND VGND VPWR VPWR _7612_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_hold2769_A _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3558__C _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4824_ _4824_/A _5531_/D _4824_/C _5531_/C VGND VGND VPWR VPWR _4830_/C sky130_fd_sc_hd__nand4_1
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7543_ _7573_/CLK _7543_/D fanout733/X VGND VGND VPWR VPWR _7543_/Q sky130_fd_sc_hd__dfstp_1
X_4755_ _4755_/A _5138_/B _5061_/B _5005_/A VGND VGND VPWR VPWR _4755_/Y sky130_fd_sc_hd__nand4_4
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3706_ _7507_/Q _3526_/X _3535_/X _7483_/Q _3705_/X VGND VGND VPWR VPWR _3706_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__3583__A2 _4431_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7474_ _7565_/CLK _7474_/D fanout746/X VGND VGND VPWR VPWR _7474_/Q sky130_fd_sc_hd__dfrtp_4
X_4686_ _5138_/B _4687_/B _4687_/C VGND VGND VPWR VPWR _5404_/A sky130_fd_sc_hd__and3_2
XFILLER_174_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6425_ _6455_/B _6434_/B _6462_/C VGND VGND VPWR VPWR _6425_/X sky130_fd_sc_hd__and3_4
X_3637_ _5992_/A _3860_/D _3637_/C VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__and3_4
XANTENNA__4532__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6356_ _7069_/Q _6110_/A _6332_/C _6075_/X _7165_/Q VGND VGND VPWR VPWR _6356_/X
+ sky130_fd_sc_hd__a32o_1
X_3568_ _3568_/A _3568_/B _3568_/C _3568_/D VGND VGND VPWR VPWR _3570_/C sky130_fd_sc_hd__nor4_2
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3201 _7157_/Q VGND VGND VPWR VPWR hold3201/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3212 hold3212/A VGND VGND VPWR VPWR _4365_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3223 _4347_/X VGND VGND VPWR VPWR hold3223/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5307_ _5297_/A _5404_/C _5410_/B _5086_/B _5061_/B VGND VGND VPWR VPWR _5308_/C
+ sky130_fd_sc_hd__a32o_1
Xhold3234 hold3234/A VGND VGND VPWR VPWR _5597_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6287_ _6962_/Q _6112_/B _6121_/B _6379_/B1 _7122_/Q VGND VGND VPWR VPWR _6287_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA_fanout587_A hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3245 _6919_/Q VGND VGND VPWR VPWR hold3245/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3499_ _7502_/Q hold41/A _3498_/X _7382_/Q _3495_/X VGND VGND VPWR VPWR _3524_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2500 hold863/X VGND VGND VPWR VPWR _5914_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2511 hold683/X VGND VGND VPWR VPWR _4556_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3256 _7343_/Q VGND VGND VPWR VPWR hold3256/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__A1 _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2522 hold941/X VGND VGND VPWR VPWR _5710_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3267 hold3267/A VGND VGND VPWR VPWR _5795_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6285__B2 _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2533 _4464_/X VGND VGND VPWR VPWR hold888/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5238_ _5222_/A _5453_/A _5453_/B _4932_/X VGND VGND VPWR VPWR _5238_/X sky130_fd_sc_hd__a31o_1
Xhold3278 _7102_/Q VGND VGND VPWR VPWR _7108_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3289 _7609_/Q VGND VGND VPWR VPWR _6284_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2544 _5979_/X VGND VGND VPWR VPWR hold610/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2555 _7531_/Q VGND VGND VPWR VPWR hold647/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1810 hold395/X VGND VGND VPWR VPWR _5931_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2566 _7668_/A VGND VGND VPWR VPWR hold617/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1821 _4392_/X VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4599__A_N _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4836__D _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1832 hold425/X VGND VGND VPWR VPWR _5733_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2577 _7397_/Q VGND VGND VPWR VPWR hold905/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout754_A _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1843 _7245_/Q VGND VGND VPWR VPWR hold429/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2588 _7420_/Q VGND VGND VPWR VPWR hold979/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5169_ _4672_/X _4956_/B _4980_/X _4692_/Y _4814_/Y VGND VGND VPWR VPWR _5169_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6037__A1 _6036_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1854 _7309_/Q VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2599 _4458_/X VGND VGND VPWR VPWR hold846/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6109__C _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1865 _7268_/Q VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1876 _4543_/X VGND VGND VPWR VPWR hold254/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1887 hold280/X VGND VGND VPWR VPWR _4519_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1898 hold437/X VGND VGND VPWR VPWR _5913_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6588__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5796__A0 _5949_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7075__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6760__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6512__A2 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5720__A0 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A mgmt_gpio_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3877__A3 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6276__B2 _7406_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3931__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4287__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6579__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output304_A _4167_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__B _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3801__A3 _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_727 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6200__A1 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6200__B2 _7515_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3675__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4270__S _4270_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4540_ _4540_/A0 _5582_/A0 _4544_/S VGND VGND VPWR VPWR _4540_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold406 hold406/A VGND VGND VPWR VPWR _7037_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4471_ _4555_/A0 _4471_/A1 _4472_/S VGND VGND VPWR VPWR _4471_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6503__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold428 hold428/A VGND VGND VPWR VPWR _7313_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold439 hold439/A VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6210_ _7419_/Q _6072_/X _6099_/X _7355_/Q _6209_/X VGND VGND VPWR VPWR _6210_/X
+ sky130_fd_sc_hd__a221o_1
X_3422_ _7466_/Q VGND VGND VPWR VPWR _3422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5711__A0 _5972_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4514__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7190_ _7191_/CLK _7190_/D fanout701/X VGND VGND VPWR VPWR _7190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6141_ _7512_/Q _6075_/A _6317_/C _6110_/X _7432_/Q VGND VGND VPWR VPWR _6141_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4937__C _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6110_/A _6144_/A _6144_/B VGND VGND VPWR VPWR _6072_/X sky130_fd_sc_hd__and3_4
XFILLER_39_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1106 hold1106/A VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold1117 hold3143/X VGND VGND VPWR VPWR hold3144/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 _5840_/X VGND VGND VPWR VPWR _7439_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5023_ _5023_/A _5023_/B VGND VGND VPWR VPWR _5025_/A sky130_fd_sc_hd__nor2_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 hold3119/X VGND VGND VPWR VPWR hold3120/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5778__A0 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4445__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ _7636_/CLK _6974_/D VGND VGND VPWR VPWR _6974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5242__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3569__B _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5925_ _5979_/A0 _5925_/A1 _5928_/S VGND VGND VPWR VPWR _5925_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5856_ hold20/X _5856_/A1 _5856_/S VGND VGND VPWR VPWR _5856_/X sky130_fd_sc_hd__mux2_1
X_4807_ _5410_/A _4807_/B _5453_/B VGND VGND VPWR VPWR _4809_/A sky130_fd_sc_hd__and3_1
X_5787_ _5787_/A0 _5922_/A0 hold48/X VGND VGND VPWR VPWR _5787_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6742__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7526_ _7572_/CLK hold78/X fanout733/X VGND VGND VPWR VPWR _7526_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4738_ _4706_/Y _4712_/Y _4734_/Y _4737_/Y _4723_/Y VGND VGND VPWR VPWR _4738_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout502_A _6089_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7457_ _7542_/CLK _7457_/D fanout719/X VGND VGND VPWR VPWR _7457_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4669_ _4570_/Y _4667_/B _4860_/A VGND VGND VPWR VPWR _4669_/X sky130_fd_sc_hd__o21a_4
XFILLER_135_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6408_ _6408_/A _6408_/B _6408_/C _6408_/D VGND VGND VPWR VPWR _6431_/A sky130_fd_sc_hd__nor4_4
XANTENNA__4505__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold940 _4487_/X VGND VGND VPWR VPWR _7143_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7388_ _7421_/CLK _7388_/D fanout716/X VGND VGND VPWR VPWR _7388_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 hold951/A VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap670 _4608_/Y VGND VGND VPWR VPWR _4899_/A2 sky130_fd_sc_hd__buf_4
Xhold962 hold962/A VGND VGND VPWR VPWR _7356_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap681 _4788_/C VGND VGND VPWR VPWR _5089_/C sky130_fd_sc_hd__clkbuf_4
Xhold973 hold973/A VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6339_ _6335_/X _6336_/X _6338_/X _6121_/C VGND VGND VPWR VPWR _6339_/X sky130_fd_sc_hd__o31a_1
Xhold984 _4536_/X VGND VGND VPWR VPWR _7184_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3020 hold3020/A VGND VGND VPWR VPWR _5858_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3031 hold3031/A VGND VGND VPWR VPWR hold3031/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3042 hold3042/A VGND VGND VPWR VPWR _5852_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4847__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3053 _7631_/Q VGND VGND VPWR VPWR _6784_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3064 hold3064/A VGND VGND VPWR VPWR hold3064/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3075 _7664_/A VGND VGND VPWR VPWR hold3075/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2330 hold603/X VGND VGND VPWR VPWR _5694_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2341 _7387_/Q VGND VGND VPWR VPWR hold557/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3086 hold3086/A VGND VGND VPWR VPWR _5741_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3097 _5641_/X VGND VGND VPWR VPWR hold3097/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2352 _4369_/X VGND VGND VPWR VPWR hold678/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2363 _5954_/X VGND VGND VPWR VPWR hold770/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2374 _5586_/X VGND VGND VPWR VPWR hold654/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1640 _7288_/Q VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2385 hold547/X VGND VGND VPWR VPWR _5988_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1651 _7270_/Q VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2396 _7012_/Q VGND VGND VPWR VPWR hold877/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1662 _7536_/Q VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1673 hold136/X VGND VGND VPWR VPWR _5936_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1684 hold75/X VGND VGND VPWR VPWR _3507_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1695 _5887_/X VGND VGND VPWR VPWR hold211/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_72_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4582__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input98_A usr2_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6733__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3547__A2 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3661__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4773__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3971_ _7209_/Q _5581_/A _3962_/X _3965_/X _3970_/X VGND VGND VPWR VPWR _3988_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_189_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5710_ _5881_/A1 _5710_/A1 _5712_/S VGND VGND VPWR VPWR _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6690_ _7193_/Q _6443_/X _6468_/X _7143_/Q _6689_/X VGND VGND VPWR VPWR _6697_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5641_ _5641_/A0 _5732_/A1 _5642_/S VGND VGND VPWR VPWR _5641_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6185__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5932__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5572_ _5572_/A _5572_/B _5572_/C VGND VGND VPWR VPWR _5572_/X sky130_fd_sc_hd__and3_1
XFILLER_129_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7311_ _7576_/CLK _7311_/D fanout717/X VGND VGND VPWR VPWR _7311_/Q sky130_fd_sc_hd__dfstp_4
X_4523_ _4523_/A0 _4547_/A0 _4526_/S VGND VGND VPWR VPWR _4523_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5824__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold214 _7377_/Q VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7242_ _7327_/CLK _7242_/D fanout703/X VGND VGND VPWR VPWR _7242_/Q sky130_fd_sc_hd__dfstp_4
Xhold225 hold225/A VGND VGND VPWR VPWR _7524_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4454_ _4454_/A0 _5853_/A0 _4454_/S VGND VGND VPWR VPWR _4454_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4499__A0 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold247 _3455_/X VGND VGND VPWR VPWR _3456_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold258 hold258/A VGND VGND VPWR VPWR _7059_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3405_ _7306_/Q VGND VGND VPWR VPWR _3405_/Y sky130_fd_sc_hd__inv_2
X_7173_ _7176_/CLK _7173_/D fanout722/X VGND VGND VPWR VPWR _7173_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout705 fanout706/X VGND VGND VPWR VPWR fanout705/X sky130_fd_sc_hd__buf_4
X_4385_ _4548_/A0 _4385_/A1 _4387_/S VGND VGND VPWR VPWR _4385_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout716 fanout720/X VGND VGND VPWR VPWR fanout716/X sky130_fd_sc_hd__buf_6
X_6124_ _6124_/A1 _6777_/S _6122_/Y _6123_/X VGND VGND VPWR VPWR _7602_/D sky130_fd_sc_hd__a22o_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout727 fanout728/X VGND VGND VPWR VPWR _6839_/A sky130_fd_sc_hd__buf_6
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3710__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout738 fanout740/X VGND VGND VPWR VPWR fanout738/X sky130_fd_sc_hd__buf_4
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 fanout750/X VGND VGND VPWR VPWR fanout749/X sky130_fd_sc_hd__buf_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6055_/A1 _6051_/Y _6054_/X VGND VGND VPWR VPWR _7597_/D sky130_fd_sc_hd__a21bo_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6660__A1 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5006_ _5495_/C1 _5528_/A3 _5046_/A _4690_/Y VGND VGND VPWR VPWR _5006_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_38_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout452_A hold40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ _7238_/CLK _6957_/D fanout690/X VGND VGND VPWR VPWR _6957_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3777__A2 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ _5998_/A1 _5908_/A1 hold42/A VGND VGND VPWR VPWR _5908_/X sky130_fd_sc_hd__mux2_1
X_6888_ _4169_/B2 _6888_/D _6838_/X VGND VGND VPWR VPWR _6888_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout717_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6176__B1 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5839_ _5866_/B _5983_/A _5992_/D VGND VGND VPWR VPWR _5847_/S sky130_fd_sc_hd__and3_4
XFILLER_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6403__B _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6715__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5923__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7509_ _7525_/CLK _7509_/D fanout748/X VGND VGND VPWR VPWR _7509_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4858__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_3__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X VGND VGND VPWR VPWR _7587_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold770 hold770/A VGND VGND VPWR VPWR _7541_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold792 _4496_/X VGND VGND VPWR VPWR _7151_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input152_A wb_dat_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3701__A2 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2160 _7526_/Q VGND VGND VPWR VPWR hold2160/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2171 _7653_/A VGND VGND VPWR VPWR hold481/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2182 hold561/X VGND VGND VPWR VPWR _4210_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2193 _7358_/Q VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1470 hold186/X VGND VGND VPWR VPWR _5971_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input13_A mask_rev_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1481 hold64/X VGND VGND VPWR VPWR _5855_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1492 hold18/X VGND VGND VPWR VPWR _4201_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5909__S hold42/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3768__A2 _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6706__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5509__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3656__C _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6182__A3 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5644__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput308 _4135_/X VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
Xoutput319 hold1129/X VGND VGND VPWR VPWR hold1130/A sky130_fd_sc_hd__buf_6
XANTENNA__3940__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3672__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5590__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4170_ _4178_/A _4427_/B VGND VGND VPWR VPWR _7106_/D sky130_fd_sc_hd__and2_1
XFILLER_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5445__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2215_A _7334_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ _4427_/D _6811_/A2 _6811_/B1 _4427_/C VGND VGND VPWR VPWR _6811_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5819__S _5820_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6742_ _7069_/Q _4101_/X _6441_/X _6443_/X _7195_/Q VGND VGND VPWR VPWR _6742_/X
+ sky130_fd_sc_hd__a32o_1
X_3954_ _7511_/Q _5920_/A _4533_/A _7182_/Q _3953_/X VGND VGND VPWR VPWR _3954_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6158__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6673_ _7182_/Q _6466_/C _6574_/C _6654_/X _6672_/X VGND VGND VPWR VPWR _6673_/X
+ sky130_fd_sc_hd__a311o_2
X_3885_ _7392_/Q _5740_/A _4431_/A _3526_/X _7504_/Q VGND VGND VPWR VPWR _3885_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5905__A0 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5624_ _5624_/A0 _5736_/A1 _5629_/S VGND VGND VPWR VPWR _5624_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5555_ _5504_/B _5551_/X _5572_/B _5550_/Y VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__a31o_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4506_ _4506_/A0 _4548_/A0 _4508_/S VGND VGND VPWR VPWR _4506_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ _5569_/A _5569_/B VGND VGND VPWR VPWR _5486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7225_ _7232_/CLK _7225_/D _4128_/B VGND VGND VPWR VPWR _7225_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5133__A1 _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4437_ _4437_/A0 _5980_/A0 _4439_/S VGND VGND VPWR VPWR _4437_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6330__B1 _6328_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_766 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout502 _6089_/C VGND VGND VPWR VPWR _6116_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_99_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_703 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout513 _5067_/C VGND VGND VPWR VPWR _5453_/C sky130_fd_sc_hd__buf_8
XFILLER_101_800 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7156_ _7185_/CLK _7156_/D fanout738/X VGND VGND VPWR VPWR _7156_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout524 _4705_/Y VGND VGND VPWR VPWR _5561_/A1 sky130_fd_sc_hd__buf_6
X_4368_ _4368_/A0 _5647_/A0 _4369_/S VGND VGND VPWR VPWR _4368_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3695__A1 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout546 hold1428/A VGND VGND VPWR VPWR _5953_/A1 sky130_fd_sc_hd__buf_6
Xfanout557 _5826_/A1 VGND VGND VPWR VPWR _5979_/A0 sky130_fd_sc_hd__buf_4
XANTENNA_input5_A mask_rev_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6107_ _7295_/Q _6136_/B _6121_/B _6379_/B1 _7391_/Q VGND VGND VPWR VPWR _6107_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_112_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout568 _5950_/A1 VGND VGND VPWR VPWR _4548_/A0 sky130_fd_sc_hd__clkbuf_8
X_7087_ _7514_/CLK _7087_/D fanout743/X VGND VGND VPWR VPWR _7666_/A sky130_fd_sc_hd__dfrtp_1
Xfanout579 _4553_/A0 VGND VGND VPWR VPWR _4547_/A0 sky130_fd_sc_hd__buf_6
X_4299_ _4302_/S _3734_/B _4298_/Y VGND VGND VPWR VPWR _6984_/D sky130_fd_sc_hd__o21ai_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6038_ _6019_/A _6929_/Q _6116_/C _6121_/B VGND VGND VPWR VPWR _6038_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6633__B2 _7294_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5729__S _5730_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7368__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6149__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1851_A _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1949_A _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_64_csclk _7399_/CLK VGND VGND VPWR VPWR _7472_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6164__A3 _7289_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_39_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6321__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3686__A1 _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3989__A2 _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7201_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6388__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5866__C _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3667__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6043__B _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _5740_/A _5992_/A _4455_/C VGND VGND VPWR VPWR _3670_/X sky130_fd_sc_hd__and3_2
XFILLER_9_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6155__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _5340_/A _5340_/B _5423_/B _5340_/D VGND VGND VPWR VPWR _5343_/C sky130_fd_sc_hd__nand4_1
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5271_ _5255_/X _4789_/Y _5473_/B _5269_/X VGND VGND VPWR VPWR _5271_/X sky130_fd_sc_hd__o211a_1
X_7010_ _7160_/CLK _7010_/D fanout700/X VGND VGND VPWR VPWR _7010_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4222_ _4222_/A0 _4221_/X _4232_/S VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__mux2_1
Xhold2907 _7189_/Q VGND VGND VPWR VPWR hold2907/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2918 _4331_/X VGND VGND VPWR VPWR hold2918/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A1 _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2929 _7159_/Q VGND VGND VPWR VPWR hold2929/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4153_ _6942_/Q _7221_/Q _6839_/B VGND VGND VPWR VPWR _4153_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4084_ _6895_/Q _4085_/A2 _6839_/B VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__o21a_2
XFILLER_110_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6379__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4986_ _5339_/A _5339_/C VGND VGND VPWR VPWR _4986_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4680__C _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3577__B _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6725_ _6715_/X _6717_/X _6724_/X _6431_/Y _6959_/Q VGND VGND VPWR VPWR _6725_/X
+ sky130_fd_sc_hd__o32a_1
X_3937_ _7311_/Q _5983_/A _3563_/C _3936_/X VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3601__A1 _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6656_ _7177_/Q _6058_/X _6457_/X _7061_/Q _6651_/X VGND VGND VPWR VPWR _6656_/X
+ sky130_fd_sc_hd__a221o_1
X_3868_ _7312_/Q _3521_/X _3553_/X input72/X _3867_/X VGND VGND VPWR VPWR _3868_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout415_A _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5607_ _5607_/A0 _5625_/A1 _5611_/S VGND VGND VPWR VPWR _5607_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4157__A2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6587_ _7300_/Q _6420_/A _6576_/X _6578_/X _6586_/X VGND VGND VPWR VPWR _6587_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6551__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3799_ _7441_/Q _3931_/B _5695_/A _4545_/A _7194_/Q VGND VGND VPWR VPWR _3799_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_191_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5538_ _5538_/A _5538_/B _5538_/C VGND VGND VPWR VPWR _5568_/B sky130_fd_sc_hd__and3_1
XANTENNA__3904__A2 _4394_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_40_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5469_ _5070_/X _5468_/X _5260_/C VGND VGND VPWR VPWR _5469_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7208_ _7633_/CLK _7208_/D _6780_/B VGND VGND VPWR VPWR _7208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7139_ _7197_/CLK _7139_/D fanout728/X VGND VGND VPWR VPWR _7139_/Q sky130_fd_sc_hd__dfstp_4
Xfanout365 _3496_/Y VGND VGND VPWR VPWR _4376_/B sky130_fd_sc_hd__buf_6
XANTENNA__6606__A1 _7309_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout387 _3557_/X VGND VGND VPWR VPWR _4265_/B sky130_fd_sc_hd__buf_12
XFILLER_86_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout398 _5614_/B VGND VGND VPWR VPWR _4479_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_47_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4574__D _4805_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input115_A wb_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__A1 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__B2 _7154_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6144__A _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5593__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6790__A0 _3643_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5983__A _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6137__A3 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input80_A spi_sck VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__buf_2
XANTENNA__6542__B1 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4765__C _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4608__B1 _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4084__A1 _6895_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4840_ _4888_/B _4888_/C _4910_/D _4840_/D VGND VGND VPWR VPWR _4840_/X sky130_fd_sc_hd__and4b_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4771_ _4700_/Y _4717_/Y _4770_/Y _4766_/Y VGND VGND VPWR VPWR _4776_/B sky130_fd_sc_hd__o211ai_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold2282_A _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6510_ _7537_/Q _6427_/A _6466_/C _6468_/C _6509_/X VGND VGND VPWR VPWR _6510_/X
+ sky130_fd_sc_hd__a41o_1
X_3722_ _6961_/Q _3657_/X _3717_/X _3719_/X _3721_/X VGND VGND VPWR VPWR _3732_/C
+ sky130_fd_sc_hd__a2111o_2
XANTENNA__3595__B1 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7490_ _7562_/CLK _7490_/D fanout740/X VGND VGND VPWR VPWR _7490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ _6433_/D _7598_/Q _7597_/Q _6441_/D VGND VGND VPWR VPWR _6441_/X sky130_fd_sc_hd__and4bb_4
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3653_ _5612_/A _4388_/B _4346_/C VGND VGND VPWR VPWR _4340_/A sky130_fd_sc_hd__and3_4
XANTENNA__6533__B1 _6451_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2547_A _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ _7180_/Q _6317_/B _6091_/X _6110_/X _7175_/Q VGND VGND VPWR VPWR _6372_/X
+ sky130_fd_sc_hd__a32o_1
X_3584_ _7405_/Q _5794_/A _3565_/X _7469_/Q _3583_/X VGND VGND VPWR VPWR _3587_/C
+ sky130_fd_sc_hd__a221o_2
X_5323_ _5183_/C _5049_/C _5339_/C _5203_/A _5339_/D VGND VGND VPWR VPWR _5324_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5832__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5254_ _4707_/Y _4709_/Y _4774_/Y _5516_/A3 VGND VGND VPWR VPWR _5254_/X sky130_fd_sc_hd__o22a_1
XFILLER_88_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2704 hold843/X VGND VGND VPWR VPWR _5585_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4956__B _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2715 _5817_/X VGND VGND VPWR VPWR hold788/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4205_ _4205_/A0 _5645_/A0 _4211_/S VGND VGND VPWR VPWR _4205_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3860__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2726 _4465_/X VGND VGND VPWR VPWR hold858/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4448__S _4448_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2737 hold927/X VGND VGND VPWR VPWR _5747_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4311__A2 _3996_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5185_ _5185_/A _5185_/B _5185_/C VGND VGND VPWR VPWR _5185_/Y sky130_fd_sc_hd__nand3_1
Xhold2748 _5605_/X VGND VGND VPWR VPWR hold762/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_3_6_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_6_0_csclk/X sky130_fd_sc_hd__clkbuf_8
Xhold2759 hold541/X VGND VGND VPWR VPWR _5696_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4136_ _7075_/Q _7072_/Q VGND VGND VPWR VPWR _4136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4862__A3 _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4067_ _6890_/Q _7071_/Q _4067_/C VGND VGND VPWR VPWR _4067_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4075__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_750 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5272__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4691__B _5012_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout532_A _4600_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4969_ _4873_/X _5528_/A3 _4672_/X _4679_/Y _4427_/B VGND VGND VPWR VPWR _4969_/Y
+ sky130_fd_sc_hd__o41ai_4
XANTENNA__6772__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3586__B1 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6708_ _7038_/Q _6462_/C _6651_/C _6707_/X VGND VGND VPWR VPWR _6708_/X sky130_fd_sc_hd__a31o_1
X_6639_ _7350_/Q _6452_/X _6468_/X _7414_/Q _6638_/X VGND VGND VPWR VPWR _6647_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6524__B1 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4212__A hold90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__7199__SET_B fanout728/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5742__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3510__B1 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4882__A _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3813__B2 _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3498__A _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__B1 _5013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6358__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7424__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5318__A1 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6515__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output284_A _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3664__C _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6818__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__A2 _6086_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4268__S _4270_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6990_ _6991_/CLK _6990_/D fanout693/X VGND VGND VPWR VPWR _6990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_80_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_8_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5941_ _5941_/A0 _5986_/A1 _5946_/S VGND VGND VPWR VPWR _5941_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3804__A1 _7521_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4942__D _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5872_ _5872_/A0 _5980_/A0 _5874_/S VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5006__B1 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7611_ _7627_/CLK _7611_/D fanout693/X VGND VGND VPWR VPWR _7611_/Q sky130_fd_sc_hd__dfrtp_1
X_4823_ _5295_/A _4823_/B _4833_/A _4823_/D VGND VGND VPWR VPWR _4824_/C sky130_fd_sc_hd__nand4_1
XANTENNA__6754__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5827__S hold33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4754_ _4803_/A _5297_/B VGND VGND VPWR VPWR _4760_/D sky130_fd_sc_hd__nand2_1
X_7542_ _7542_/CLK _7542_/D fanout713/X VGND VGND VPWR VPWR _7542_/Q sky130_fd_sc_hd__dfrtp_4
X_3705_ _7045_/Q _4370_/A _3665_/X _7126_/Q VGND VGND VPWR VPWR _3705_/X sky130_fd_sc_hd__a22o_1
XFILLER_186_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7473_ _7537_/CLK _7473_/D fanout709/X VGND VGND VPWR VPWR _7473_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__5309__B2 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4685_ _4593_/A _4591_/Y _4593_/Y VGND VGND VPWR VPWR _4822_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__3583__A3 _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6424_ _6427_/A _6455_/B _6447_/B VGND VGND VPWR VPWR _6424_/X sky130_fd_sc_hd__and3_4
X_3636_ input8/X _3486_/X _3529_/X _7532_/Q _3635_/X VGND VGND VPWR VPWR _3642_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6355_ _6355_/A1 _4116_/X _6067_/X _6354_/X VGND VGND VPWR VPWR _7612_/D sky130_fd_sc_hd__o31a_1
X_3567_ _7334_/Q _5713_/A _3563_/X _3566_/X _3560_/X VGND VGND VPWR VPWR _3568_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6809__A1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3202 hold3202/A VGND VGND VPWR VPWR _4504_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5306_ _5306_/A _5306_/B VGND VGND VPWR VPWR _5308_/B sky130_fd_sc_hd__nand2_1
Xhold3213 _7177_/Q VGND VGND VPWR VPWR hold3213/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3224 _7224_/Q VGND VGND VPWR VPWR hold3224/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6286_ _7011_/Q _6384_/A4 _6120_/B _6110_/A VGND VGND VPWR VPWR _6286_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3235 _6941_/Q VGND VGND VPWR VPWR hold3235/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3498_ _5740_/A _3682_/A _4455_/A VGND VGND VPWR VPWR _3498_/X sky130_fd_sc_hd__and3_4
Xhold3246 hold3246/A VGND VGND VPWR VPWR _4204_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3590__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2501 _7355_/Q VGND VGND VPWR VPWR hold621/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2512 _4556_/X VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3257 hold3257/A VGND VGND VPWR VPWR _5732_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5237_ _5208_/Y _5237_/B _5237_/C VGND VGND VPWR VPWR _5237_/Y sky130_fd_sc_hd__nand3b_1
Xhold2523 _5710_/X VGND VGND VPWR VPWR hold942/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3268 _7219_/Q VGND VGND VPWR VPWR _3645_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2534 _7372_/Q VGND VGND VPWR VPWR hold931/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3279 _6792_/S VGND VGND VPWR VPWR _6789_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2545 _7412_/Q VGND VGND VPWR VPWR hold945/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1800 hold45/X VGND VGND VPWR VPWR _3475_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2556 hold647/X VGND VGND VPWR VPWR _5943_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1811 _5931_/X VGND VGND VPWR VPWR hold396/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1822 _7304_/Q VGND VGND VPWR VPWR hold351/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2567 hold617/X VGND VGND VPWR VPWR _4436_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5168_ _4849_/X _5061_/X _5167_/Y _5294_/A VGND VGND VPWR VPWR _5168_/X sky130_fd_sc_hd__o31a_1
Xhold1833 _5733_/X VGND VGND VPWR VPWR hold426/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2578 hold905/X VGND VGND VPWR VPWR _5792_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1844 hold429/X VGND VGND VPWR VPWR _5616_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2589 hold979/X VGND VGND VPWR VPWR _5818_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1855 hold238/X VGND VGND VPWR VPWR _5693_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4119_ _6009_/B _4107_/Y _4105_/Y _7256_/Q _6929_/Q VGND VGND VPWR VPWR _6931_/D
+ sky130_fd_sc_hd__a32o_1
Xhold1866 hold286/X VGND VGND VPWR VPWR _5647_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1877 _7019_/Q VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout747_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5099_ _4798_/Y _4960_/A _5098_/Y VGND VGND VPWR VPWR _5099_/Y sky130_fd_sc_hd__o21ai_1
Xhold1888 _4519_/X VGND VGND VPWR VPWR hold281/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5245__B1 _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1899 _5913_/X VGND VGND VPWR VPWR hold438/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6588__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6745__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3559__B1 _3558_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1764_A _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6422__A _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6760__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3574__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5038__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3484__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3731__B1 _3727_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4596__B _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input43_A mgmt_gpio_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3931__D _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6579__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5251__A3 _5342_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3659__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6736__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5647__S _5649_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6200__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4211__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3675__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4470_ _5914_/A1 _4470_/A1 _4472_/S VGND VGND VPWR VPWR _4470_/X sky130_fd_sc_hd__mux2_1
Xhold407 hold407/A VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5199__A_N _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold418 hold418/A VGND VGND VPWR VPWR _7353_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6503__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3421_ _7474_/Q VGND VGND VPWR VPWR _3421_/Y sky130_fd_sc_hd__inv_2
Xhold429 hold429/A VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6140_ _7416_/Q _6072_/X _6097_/X _7440_/Q _6139_/X VGND VGND VPWR VPWR _6140_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_98_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6267__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _7589_/Q _7588_/Q _6121_/B VGND VGND VPWR VPWR _6071_/X sky130_fd_sc_hd__and3b_2
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 hold2842/X VGND VGND VPWR VPWR hold2843/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5022_ _5029_/A _5180_/A _5216_/A VGND VGND VPWR VPWR _5023_/A sky130_fd_sc_hd__and3_1
Xhold1118 hold3145/X VGND VGND VPWR VPWR _7041_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 hold3047/X VGND VGND VPWR VPWR hold1129/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6973_ _7630_/CLK _6973_/D VGND VGND VPWR VPWR _6973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3789__B1 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5924_ _5978_/A0 _5924_/A1 _5928_/S VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2879_A _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3569__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4450__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5855_ _5990_/A1 _5855_/A1 _5856_/S VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4806_ _5100_/A _5260_/B VGND VGND VPWR VPWR _4806_/Y sky130_fd_sc_hd__nand2_2
XFILLER_166_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4202__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5786_ _5786_/A0 _5993_/A1 hold48/X VGND VGND VPWR VPWR _5786_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6742__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7525_ _7525_/CLK _7525_/D fanout746/X VGND VGND VPWR VPWR _7525_/Q sky130_fd_sc_hd__dfrtp_4
X_4737_ _5100_/A _5079_/B VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__5950__A1 _5950_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7456_ _7576_/CLK _7456_/D fanout718/X VGND VGND VPWR VPWR _7456_/Q sky130_fd_sc_hd__dfstp_2
X_4668_ _4984_/B _4805_/B _4668_/C _4797_/B VGND VGND VPWR VPWR _4974_/C sky130_fd_sc_hd__nand4_4
XFILLER_174_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2__f_wb_clk_i clkbuf_3_1_0_wb_clk_i/X VGND VGND VPWR VPWR _6999_/CLK sky130_fd_sc_hd__clkbuf_16
X_3619_ _7614_/Q _7253_/Q _7255_/Q VGND VGND VPWR VPWR _3619_/X sky130_fd_sc_hd__mux2_8
X_6407_ _6427_/A _6466_/C _6468_/C VGND VGND VPWR VPWR _6408_/D sky130_fd_sc_hd__and3_4
XANTENNA__5702__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold930 hold930/A VGND VGND VPWR VPWR _7577_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold941 hold941/A VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4599_ _4888_/C _4888_/B VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__nand2b_4
X_7387_ _7580_/CLK _7387_/D fanout734/X VGND VGND VPWR VPWR _7387_/Q sky130_fd_sc_hd__dfrtp_4
Xhold952 hold952/A VGND VGND VPWR VPWR _7200_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout697_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap671 _5387_/B VGND VGND VPWR VPWR _5399_/B sky130_fd_sc_hd__buf_8
Xhold963 hold963/A VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6338_ _7013_/Q _6136_/B _6120_/B _6337_/X VGND VGND VPWR VPWR _6338_/X sky130_fd_sc_hd__a31o_1
Xhold3010 hold3010/A VGND VGND VPWR VPWR hold3010/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold974 hold974/A VGND VGND VPWR VPWR _6963_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold985 hold985/A VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3021 _5858_/X VGND VGND VPWR VPWR hold3021/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold996 hold996/A VGND VGND VPWR VPWR _7140_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3032 _7383_/Q VGND VGND VPWR VPWR hold3032/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3043 _5852_/X VGND VGND VPWR VPWR hold3043/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6269_ _7534_/Q _6080_/A _6091_/X _6121_/X _7310_/Q VGND VGND VPWR VPWR _6269_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3054 hold3054/A VGND VGND VPWR VPWR hold3054/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2320 _5909_/X VGND VGND VPWR VPWR hold748/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4269__A1 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3065 _7375_/Q VGND VGND VPWR VPWR hold3065/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2331 _5694_/X VGND VGND VPWR VPWR hold604/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3076 hold3076/A VGND VGND VPWR VPWR _4432_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2342 hold557/X VGND VGND VPWR VPWR _5781_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3087 _5741_/X VGND VGND VPWR VPWR hold3087/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3098 _7271_/Q VGND VGND VPWR VPWR hold3098/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2353 _7332_/Q VGND VGND VPWR VPWR hold795/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2364 _7540_/Q VGND VGND VPWR VPWR hold797/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2375 _7250_/Q VGND VGND VPWR VPWR hold611/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1630 _3449_/X VGND VGND VPWR VPWR _3459_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1641 hold379/X VGND VGND VPWR VPWR _5670_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2386 _7052_/Q VGND VGND VPWR VPWR hold805/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1652 hold312/X VGND VGND VPWR VPWR _5649_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2397 hold877/X VGND VGND VPWR VPWR _4336_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1663 hold385/X VGND VGND VPWR VPWR _5949_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6417__A _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1674 _5936_/X VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1685 _3507_/X VGND VGND VPWR VPWR hold1685/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1696 _7568_/Q VGND VGND VPWR VPWR hold381/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5769__A1 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6136__B _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4441__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6718__B1 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6194__A1 _7323_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5941__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4400__A _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6249__A2 _6072_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5930__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5209__B1 _4946_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3970_ _7495_/Q hold41/A _3969_/X _3931_/X _3968_/X VGND VGND VPWR VPWR _3970_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4432__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6709__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5640_ _5640_/A _5640_/B _5640_/C _5640_/D VGND VGND VPWR VPWR _5642_/S sky130_fd_sc_hd__and4_1
XANTENNA__6185__A1 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6185__B2 _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5571_ _5038_/B _5339_/B _5030_/C _5570_/X _5435_/D VGND VGND VPWR VPWR _5572_/C
+ sky130_fd_sc_hd__a311oi_4
X_7310_ _7541_/CLK _7310_/D fanout710/X VGND VGND VPWR VPWR _7310_/Q sky130_fd_sc_hd__dfrtp_4
X_4522_ _4522_/A0 _5876_/A1 _4526_/S VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold204 hold204/A VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6488__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7241_ _7327_/CLK _7241_/D fanout703/X VGND VGND VPWR VPWR _7241_/Q sky130_fd_sc_hd__dfstp_2
Xhold226 hold226/A VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4453_ _4453_/A0 _4555_/A0 _4454_/S VGND VGND VPWR VPWR _4453_/X sky130_fd_sc_hd__mux2_1
Xhold237 hold237/A VGND VGND VPWR VPWR _7064_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold248 _3456_/X VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3404_ _4674_/A VGND VGND VPWR VPWR _5089_/B sky130_fd_sc_hd__inv_12
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4310__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7172_ _7176_/CLK _7172_/D fanout722/X VGND VGND VPWR VPWR _7172_/Q sky130_fd_sc_hd__dfrtp_4
X_4384_ _4547_/A0 _4384_/A1 _4387_/S VGND VGND VPWR VPWR _4384_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout706 fanout720/X VGND VGND VPWR VPWR fanout706/X sky130_fd_sc_hd__buf_4
X_6123_ _7279_/Q _6036_/Y _6623_/B1 _6067_/B VGND VGND VPWR VPWR _6123_/X sky130_fd_sc_hd__o211a_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout717 fanout720/X VGND VGND VPWR VPWR fanout717/X sky130_fd_sc_hd__buf_6
Xfanout728 fanout750/X VGND VGND VPWR VPWR fanout728/X sky130_fd_sc_hd__buf_8
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 fanout740/X VGND VGND VPWR VPWR fanout739/X sky130_fd_sc_hd__buf_8
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6054_ _6050_/Y _6067_/B _7597_/Q _6019_/Y VGND VGND VPWR VPWR _6054_/X sky130_fd_sc_hd__a211o_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5005_/A _5005_/B _5005_/C VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__nand3_4
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4671__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6902__CLK _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A3 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6956_ _7578_/CLK hold57/X fanout747/X VGND VGND VPWR VPWR _6956_/Q sky130_fd_sc_hd__dfrtp_1
X_5907_ _5952_/A1 _5907_/A1 hold42/X VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__mux2_1
X_6887_ _4169_/B2 _6887_/D _6837_/X VGND VGND VPWR VPWR _6887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6176__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5838_ _5838_/A0 hold20/X _5838_/S VGND VGND VPWR VPWR _5838_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__B2 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5769_ _5769_/A0 _5976_/A0 _5775_/S VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7508_ _7574_/CLK _7508_/D fanout745/X VGND VGND VPWR VPWR _7508_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6479__A2 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7439_ _7519_/CLK _7439_/D fanout741/X VGND VGND VPWR VPWR _7439_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__5687__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold760 hold760/A VGND VGND VPWR VPWR _7030_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5151__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold771 hold771/A VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold782 hold782/A VGND VGND VPWR VPWR _7349_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5439__B1 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input145_A wb_dat_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2150 hold2150/A VGND VGND VPWR VPWR _5793_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2161 hold2161/A VGND VGND VPWR VPWR _5937_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2172 hold481/X VGND VGND VPWR VPWR _4249_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2183 _7409_/Q VGND VGND VPWR VPWR hold595/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2194 hold244/X VGND VGND VPWR VPWR _5748_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1460 _6954_/Q VGND VGND VPWR VPWR hold140/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_18_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1471 _5971_/X VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold3108_A _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1482 _5855_/X VGND VGND VPWR VPWR hold65/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1493 _4201_/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4414__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5914__A1 _5914_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput309 _7672_/X VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3672__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__A2 _4690_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6642__A2 _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6810_ _6809_/X _6810_/A1 _6822_/S VGND VGND VPWR VPWR _7640_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6741_ _7160_/Q _6419_/A _6447_/X _7185_/Q _6740_/X VGND VGND VPWR VPWR _6749_/B
+ sky130_fd_sc_hd__a221o_1
X_3953_ _7132_/Q _4473_/A _5619_/B _3506_/X _7351_/Q VGND VGND VPWR VPWR _3953_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4950__D _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6158__A1 _7377_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6158__B2 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6672_ _6962_/Q _6422_/X _6656_/X _6666_/X _6671_/X VGND VGND VPWR VPWR _6672_/X
+ sky130_fd_sc_hd__a2111o_1
X_3884_ _7528_/Q _3529_/X _3661_/X _7032_/Q _3883_/X VGND VGND VPWR VPWR _3884_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5623_ _5640_/C _5623_/B _5640_/D VGND VGND VPWR VPWR _5629_/S sky130_fd_sc_hd__and3_4
XANTENNA__5835__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3916__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5554_ _5554_/A _5554_/B _5554_/C VGND VGND VPWR VPWR _5572_/B sky130_fd_sc_hd__and3_1
XFILLER_117_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3863__B _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4505_ _4505_/A0 hold198/X _4508_/S VGND VGND VPWR VPWR _4505_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5485_ _5408_/Y _4713_/X _5143_/C _5303_/A VGND VGND VPWR VPWR _5569_/B sky130_fd_sc_hd__o211a_1
XANTENNA__5669__A0 hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4436_ _4436_/A0 _5979_/A0 _4439_/S VGND VGND VPWR VPWR _4436_/X sky130_fd_sc_hd__mux2_1
X_7224_ _7232_/CLK _7224_/D _4128_/B VGND VGND VPWR VPWR _7224_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout503 _6022_/X VGND VGND VPWR VPWR _6136_/B sky130_fd_sc_hd__buf_8
XFILLER_160_778 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4367_ _4367_/A0 _4548_/A0 _4369_/S VGND VGND VPWR VPWR _4367_/X sky130_fd_sc_hd__mux2_1
Xfanout514 wire516/X VGND VGND VPWR VPWR _5282_/C sky130_fd_sc_hd__clkbuf_8
X_7155_ _7185_/CLK _7155_/D fanout725/X VGND VGND VPWR VPWR _7155_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout525 _4705_/Y VGND VGND VPWR VPWR _5563_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout547 hold1428/A VGND VGND VPWR VPWR _5881_/A1 sky130_fd_sc_hd__buf_4
XFILLER_113_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6106_ _7591_/Q _7590_/Q _6136_/B VGND VGND VPWR VPWR _6106_/X sky130_fd_sc_hd__and3_2
XFILLER_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7086_ _7514_/CLK _7086_/D fanout743/X VGND VGND VPWR VPWR _7665_/A sky130_fd_sc_hd__dfrtp_1
Xfanout558 _5673_/A0 VGND VGND VPWR VPWR _5826_/A1 sky130_fd_sc_hd__buf_6
Xfanout569 _5968_/A1 VGND VGND VPWR VPWR _5950_/A1 sky130_fd_sc_hd__clkbuf_8
X_4298_ _4302_/S _4298_/B VGND VGND VPWR VPWR _4298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6633__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6037_ _6036_/Y _6019_/A _6019_/Y VGND VGND VPWR VPWR _6037_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout562_A _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ _7578_/CLK _6939_/D fanout747/X VGND VGND VPWR VPWR _6939_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6149__A1 _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6554__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5745__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__B1 _4485_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_csclk _4169_/X VGND VGND VPWR VPWR clkbuf_0_csclk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__4134__A_N _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5046__A _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3492__C _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6321__A1 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold590 hold590/A VGND VGND VPWR VPWR _7331_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4885__A _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3686__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4635__A1 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3989__A3 _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1290 _5591_/X VGND VGND VPWR VPWR _7224_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4399__A0 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3667__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3610__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5899__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2158_A _7158_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5270_ _4698_/Y _5561_/A1 _4946_/Y _4789_/Y _5480_/B2 VGND VGND VPWR VPWR _5473_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6312__A1 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4323__A0 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4221_ _4253_/A0 _5986_/A1 _4231_/S VGND VGND VPWR VPWR _4221_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2908 hold2908/A VGND VGND VPWR VPWR _4542_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2919 _7466_/Q VGND VGND VPWR VPWR hold2919/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4874__B2 _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4152_ _6947_/Q input77/X _4173_/B VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__mux2_8
XANTENNA__6076__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6615__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4083_ _7600_/Q _7250_/Q _7255_/Q VGND VGND VPWR VPWR _4117_/B sky130_fd_sc_hd__mux2_8
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ _5328_/A _5328_/B _5339_/C VGND VGND VPWR VPWR _5030_/C sky130_fd_sc_hd__and3_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6724_ _6431_/A _6411_/Y _6431_/C _6723_/X VGND VGND VPWR VPWR _6724_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3936_ _7543_/Q _4479_/A _5956_/B _3654_/X _7117_/Q VGND VGND VPWR VPWR _3936_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_176_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_2_0_csclk clkbuf_0_csclk/X VGND VGND VPWR VPWR clkbuf_3_2_0_csclk/X sky130_fd_sc_hd__clkbuf_8
X_6655_ _7066_/Q _4101_/X _6441_/X _6425_/X _7016_/Q VGND VGND VPWR VPWR _6655_/X
+ sky130_fd_sc_hd__a32o_1
X_3867_ _7336_/Q _3531_/X _3667_/X _7022_/Q _3863_/X VGND VGND VPWR VPWR _3867_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_191_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5606_ _5606_/A0 _5815_/A1 _5611_/S VGND VGND VPWR VPWR _5606_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4157__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6551__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6586_ _7540_/Q _6408_/D _6582_/X _6585_/X VGND VGND VPWR VPWR _6586_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6551__B2 _7347_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3798_ _7569_/Q _5983_/A _4479_/A _3654_/X _7119_/Q VGND VGND VPWR VPWR _3798_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_192_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5537_ _4706_/Y _4735_/Y _4760_/D _5536_/Y VGND VGND VPWR VPWR _5538_/C sky130_fd_sc_hd__o211a_1
XFILLER_117_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5106__A2 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5468_ _5100_/A _5079_/B _4807_/B _4823_/D _5134_/A VGND VGND VPWR VPWR _5468_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_160_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7207_ _7630_/CLK _7207_/D _6780_/B VGND VGND VPWR VPWR _7207_/Q sky130_fd_sc_hd__dfrtp_1
X_4419_ _4419_/A0 _4418_/X _4423_/S VGND VGND VPWR VPWR _4419_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5399_ _5399_/A _5399_/B _5399_/C _5399_/D VGND VGND VPWR VPWR _5481_/B sky130_fd_sc_hd__nand4_1
X_7138_ _7197_/CLK _7138_/D fanout742/X VGND VGND VPWR VPWR _7138_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout366 hold31/X VGND VGND VPWR VPWR _3931_/B sky130_fd_sc_hd__buf_8
XANTENNA__6606__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout388 _3548_/X VGND VGND VPWR VPWR _5619_/B sky130_fd_sc_hd__clkbuf_16
X_7069_ _7191_/CLK _7069_/D _6872_/A VGND VGND VPWR VPWR _7069_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout399 _5965_/A VGND VGND VPWR VPWR _3637_/C sky130_fd_sc_hd__buf_6
XANTENNA__4617__A1 _4570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__C _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A wb_adr_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6144__B _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6542__A1 _7474_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6542__B2 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4553__A0 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input73_A pad_flash_io0_di VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4608__A1 _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4084__A2 _4085_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5596__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4770_ _5260_/C _5113_/A _5404_/C _5410_/B VGND VGND VPWR VPWR _4770_/Y sky130_fd_sc_hd__nand4_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5893__B _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3721_ input16/X _3490_/X _5581_/A _7213_/Q _3720_/X VGND VGND VPWR VPWR _3721_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3595__B2 _7533_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6440_ _7575_/Q _6427_/X _6432_/X _6439_/X _6430_/X VGND VGND VPWR VPWR _6440_/Y
+ sky130_fd_sc_hd__a2111oi_4
XANTENNA__6533__A1 _7354_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3652_ _3860_/D _4479_/A _4491_/C VGND VGND VPWR VPWR _3652_/X sky130_fd_sc_hd__and3_2
XANTENNA__6533__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_162_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6371_ _7044_/Q _6089_/X _6082_/C _7064_/Q _6100_/X VGND VGND VPWR VPWR _6371_/X
+ sky130_fd_sc_hd__a32o_1
X_3583_ _7525_/Q _4431_/A _5938_/C _3553_/X input41/X VGND VGND VPWR VPWR _3583_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_173_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_csclk_A _7416_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3898__A2 _4551_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5322_ _5496_/B _5320_/X _5321_/X _5294_/Y VGND VGND VPWR VPWR _5322_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_154_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6297__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5253_ _5134_/A _5282_/B _5524_/A3 _5107_/X VGND VGND VPWR VPWR _5278_/D sky130_fd_sc_hd__a31oi_1
Xhold2705 _5585_/X VGND VGND VPWR VPWR hold844/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4204_ _4204_/A0 _5732_/A1 _4211_/S VGND VGND VPWR VPWR _4204_/X sky130_fd_sc_hd__mux2_1
Xhold2716 _7433_/Q VGND VGND VPWR VPWR hold981/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3860__C _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5184_ _5495_/C1 _5528_/A3 _5046_/A _5183_/Y VGND VGND VPWR VPWR _5184_/X sky130_fd_sc_hd__o31a_1
Xhold2727 _7035_/Q VGND VGND VPWR VPWR hold775/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2738 _5747_/X VGND VGND VPWR VPWR hold928/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2749 _7581_/Q VGND VGND VPWR VPWR hold965/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4135_ _6896_/Q _4135_/B VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__and2b_4
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_63_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7542_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4066_ _6891_/Q _4098_/A1 _4058_/A _4067_/C _4065_/Y VGND VGND VPWR VPWR _4066_/Y
+ sky130_fd_sc_hd__o41ai_1
XFILLER_37_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4691__C _5328_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3822__A2 _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4968_ _4873_/X _5528_/A3 _4672_/X _4679_/Y _4427_/B VGND VGND VPWR VPWR _4968_/X
+ sky130_fd_sc_hd__o41a_1
X_6707_ _7063_/Q _6466_/C _6441_/X _6058_/X _7179_/Q VGND VGND VPWR VPWR _6707_/X
+ sky130_fd_sc_hd__a32o_1
X_3919_ _7304_/Q _5686_/A _3914_/X _3915_/X _3918_/X VGND VGND VPWR VPWR _3919_/X
+ sky130_fd_sc_hd__a2111o_4
X_4899_ _4667_/A _4899_/A2 _4657_/C wire649/X _5213_/C VGND VGND VPWR VPWR _4899_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__5327__A2 _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6638_ _7478_/Q _6574_/B _6441_/X _6443_/X _7454_/Q VGND VGND VPWR VPWR _6638_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6524__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6524__B2 _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4535__A0 _4553_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_818 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6569_ _6569_/A _6569_/B _6569_/C _6569_/D VGND VGND VPWR VPWR _6570_/C sky130_fd_sc_hd__nor4_2
XANTENNA__3889__A2 _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6288__B1 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_csclk clkbuf_3_5_0_csclk/X VGND VGND VPWR VPWR _7186_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4866__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_csclk_A clkbuf_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3510__B2 input33/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__7070__RESET_B _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5263__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3813__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__B _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5015__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5318__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6515__B2 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5933__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6279__B1 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3453__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5254__B2 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5940_ _5940_/A0 _5985_/A1 _5946_/S VGND VGND VPWR VPWR _5940_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3804__A2 hold77/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5871_ _5871_/A0 _5979_/A0 _5871_/S VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6203__B1 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7610_ _7610_/CLK _7610_/D fanout693/X VGND VGND VPWR VPWR _7610_/Q sky130_fd_sc_hd__dfrtp_1
X_4822_ _5138_/A _5138_/C _5029_/A _4822_/D VGND VGND VPWR VPWR _5531_/D sky130_fd_sc_hd__nand4_4
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7541_ _7541_/CLK _7541_/D fanout713/X VGND VGND VPWR VPWR _7541_/Q sky130_fd_sc_hd__dfrtp_4
X_4753_ _4778_/A _4767_/B _4753_/C VGND VGND VPWR VPWR _5297_/B sky130_fd_sc_hd__and3_2
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4313__A _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3704_ _6878_/Q _5866_/B _3514_/X _3703_/X VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__a31o_1
X_7472_ _7472_/CLK _7472_/D fanout719/X VGND VGND VPWR VPWR _7472_/Q sky130_fd_sc_hd__dfstp_2
X_4684_ _4825_/A _4593_/A _4592_/X VGND VGND VPWR VPWR _5138_/B sky130_fd_sc_hd__a21oi_4
X_6423_ _6463_/A _6455_/B _6462_/C VGND VGND VPWR VPWR _6423_/X sky130_fd_sc_hd__and3_4
Xclkbuf_4_1__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X VGND VGND VPWR VPWR _7594_/CLK sky130_fd_sc_hd__clkbuf_16
X_3635_ _7492_/Q _5947_/B _5965_/B _3565_/X _7468_/Q VGND VGND VPWR VPWR _3635_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6354_ _6009_/B _6354_/A2 _6777_/S _6353_/X VGND VGND VPWR VPWR _6354_/X sky130_fd_sc_hd__a211o_1
X_3566_ _7366_/Q _4364_/A _5965_/B _3565_/X _7470_/Q VGND VGND VPWR VPWR _3566_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3203 _6957_/Q VGND VGND VPWR VPWR hold3203/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3740__A1 _7570_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5305_ _4716_/Y _4723_/Y _4978_/Y _4713_/X _5304_/X VGND VGND VPWR VPWR _5306_/B
+ sky130_fd_sc_hd__o221a_1
Xhold3214 hold3214/A VGND VGND VPWR VPWR _4528_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3740__B2 input64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3497_ hold40/X _4328_/A _5947_/B VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__and3_4
X_6285_ _7001_/Q _6097_/B _6120_/B _6332_/C _7031_/Q VGND VGND VPWR VPWR _6285_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3225 hold3225/A VGND VGND VPWR VPWR _5591_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3236 hold3236/A VGND VGND VPWR VPWR _4235_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3247 _7327_/Q VGND VGND VPWR VPWR hold3247/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3590__C _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2502 hold621/X VGND VGND VPWR VPWR _5745_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3258 _5732_/X VGND VGND VPWR VPWR hold3258/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2513 _7428_/Q VGND VGND VPWR VPWR hold955/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6285__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5236_ _4799_/C _4885_/X _4927_/B VGND VGND VPWR VPWR _5237_/C sky130_fd_sc_hd__a21oi_1
Xhold2524 _7269_/Q VGND VGND VPWR VPWR hold659/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3269 _3645_/X VGND VGND VPWR VPWR _7219_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2535 hold931/X VGND VGND VPWR VPWR _5764_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2546 hold945/X VGND VGND VPWR VPWR _5809_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1801 _3475_/X VGND VGND VPWR VPWR _3500_/B sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2557 _5943_/X VGND VGND VPWR VPWR hold648/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4983__A _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1812 _7206_/Q VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1823 hold351/X VGND VGND VPWR VPWR _5688_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5167_ _5167_/A _5529_/A _5496_/B _5496_/A VGND VGND VPWR VPWR _5167_/Y sky130_fd_sc_hd__nand4_1
Xhold2568 _7047_/Q VGND VGND VPWR VPWR hold935/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1834 _7448_/Q VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2579 _7131_/Q VGND VGND VPWR VPWR hold731/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1845 _7069_/Q VGND VGND VPWR VPWR hold267/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4118_ _4107_/A _6009_/B _6019_/A _4116_/X VGND VGND VPWR VPWR _6930_/D sky130_fd_sc_hd__a211o_1
Xhold1856 _5693_/X VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1867 _5647_/X VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5098_ _4748_/A _5091_/A _4797_/X _5097_/Y VGND VGND VPWR VPWR _5098_/Y sky130_fd_sc_hd__a31oi_1
Xhold1878 hold320/X VGND VGND VPWR VPWR _4344_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5245__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1889 _7326_/Q VGND VGND VPWR VPWR hold178/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6442__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5245__B2 _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4049_ _6908_/Q _4058_/A _6910_/Q _6909_/Q VGND VGND VPWR VPWR _4050_/S sky130_fd_sc_hd__and4b_1
XFILLER_25_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3559__A1 _7542_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5181__B1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4877__B _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3731__A1 _4177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_161_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6276__A3 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3138_A _7031_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input36_A mgmt_gpio_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3495__B1 _3494_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3798__A1 _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3798__B2 _7119_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4117__B _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6736__A1 _7044_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6200__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3675__C _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6051__C _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire350 _6733_/Y VGND VGND VPWR VPWR wire350/X sky130_fd_sc_hd__clkbuf_4
Xhold408 _4505_/X VGND VGND VPWR VPWR _7158_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold419 hold419/A VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3420_ _7482_/Q VGND VGND VPWR VPWR _3420_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4787__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3722__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _6332_/B _6119_/B _6116_/C _6119_/A VGND VGND VPWR VPWR _6070_/X sky130_fd_sc_hd__and4bb_4
XANTENNA__6267__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5475__A1 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 hold2844/X VGND VGND VPWR VPWR _6947_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5021_ _5021_/A _5021_/B _5021_/C _5021_/D VGND VGND VPWR VPWR _5023_/B sky130_fd_sc_hd__nand4_1
Xhold1119 hold3138/X VGND VGND VPWR VPWR hold3139/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2405_A _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6972_ _7000_/CLK _6972_/D VGND VGND VPWR VPWR _6972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3789__A1 _7346_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5923_ _5986_/A1 _5923_/A1 _5928_/S VGND VGND VPWR VPWR _5923_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5838__S _5838_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5854_ _5998_/A1 _5854_/A1 _5856_/S VGND VGND VPWR VPWR _5854_/X sky130_fd_sc_hd__mux2_1
X_4805_ _4984_/B _4805_/B _5260_/B VGND VGND VPWR VPWR _5453_/B sky130_fd_sc_hd__and3_4
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5785_ hold47/X _5785_/B _5992_/D VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__and3_1
XFILLER_166_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7524_ _7574_/CLK _7524_/D fanout733/X VGND VGND VPWR VPWR _7524_/Q sky130_fd_sc_hd__dfrtp_4
X_4736_ _4786_/D _4767_/A _4831_/C VGND VGND VPWR VPWR _5074_/B sky130_fd_sc_hd__and3b_4
XFILLER_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7455_ _7528_/CLK _7455_/D fanout729/X VGND VGND VPWR VPWR _7455_/Q sky130_fd_sc_hd__dfstp_2
X_4667_ _4667_/A _4667_/B _4667_/C VGND VGND VPWR VPWR _4667_/Y sky130_fd_sc_hd__nor3_2
XFILLER_119_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6406_ _7594_/Q _7597_/Q _7598_/Q _6455_/B VGND VGND VPWR VPWR _6408_/C sky130_fd_sc_hd__and4bb_4
X_3618_ _7332_/Q _3933_/A _5731_/B _3521_/X _7316_/Q VGND VGND VPWR VPWR _3618_/X
+ sky130_fd_sc_hd__a32o_1
Xhold920 _4360_/X VGND VGND VPWR VPWR _7032_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4697__B _4797_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold931 hold931/A VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7386_ _7548_/CLK _7386_/D fanout732/X VGND VGND VPWR VPWR _7386_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4598_ _4888_/C _4888_/B VGND VGND VPWR VPWR _5399_/A sky130_fd_sc_hd__and2b_4
Xhold942 hold942/A VGND VGND VPWR VPWR _7324_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3713__A1 _7291_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold953 hold953/A VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3713__B2 _3503_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6337_ _6964_/Q _6112_/B _6121_/B _6379_/B1 _7124_/Q VGND VGND VPWR VPWR _6337_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold964 _4501_/X VGND VGND VPWR VPWR _7155_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout592_A hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold975 hold975/A VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3000 hold3000/A VGND VGND VPWR VPWR hold3000/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3549_ _5992_/A _3637_/C _4455_/C VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__and3_4
Xhold3011 _6996_/Q VGND VGND VPWR VPWR _4315_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold986 _5896_/X VGND VGND VPWR VPWR _7489_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3022 _7632_/Q VGND VGND VPWR VPWR _6786_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3033 hold3033/A VGND VGND VPWR VPWR _5777_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold997 hold997/A VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6268_ _7478_/Q _6032_/Y _6267_/X _6144_/C VGND VGND VPWR VPWR _6268_/X sky130_fd_sc_hd__a211o_1
Xhold3044 _7391_/Q VGND VGND VPWR VPWR hold3044/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2310 hold573/X VGND VGND VPWR VPWR _4243_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3055 _7431_/Q VGND VGND VPWR VPWR hold3055/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5466__A1 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2321 _7228_/Q VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3066 hold3066/A VGND VGND VPWR VPWR _5768_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2332 _7321_/Q VGND VGND VPWR VPWR hold717/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3077 _7244_/Q VGND VGND VPWR VPWR hold3077/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6663__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5219_ _4741_/Y _4886_/Y _4896_/Y _4903_/Y _5218_/Y VGND VGND VPWR VPWR _5219_/Y
+ sky130_fd_sc_hd__o2111ai_1
Xhold3088 _7656_/A VGND VGND VPWR VPWR hold3088/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2343 _5781_/X VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3099 hold3099/A VGND VGND VPWR VPWR _5651_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2354 hold795/X VGND VGND VPWR VPWR _5719_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6199_ _7483_/Q _6112_/X _6197_/X _6198_/X _6196_/X VGND VGND VPWR VPWR _6212_/B
+ sky130_fd_sc_hd__a2111o_2
Xhold2365 hold797/X VGND VGND VPWR VPWR _5953_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1620 _5675_/X VGND VGND VPWR VPWR hold171/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2376 hold611/X VGND VGND VPWR VPWR _5624_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1631 _3459_/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1642 _5670_/X VGND VGND VPWR VPWR hold380/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2387 hold805/X VGND VGND VPWR VPWR _4384_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1653 _5649_/X VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2398 _4336_/X VGND VGND VPWR VPWR hold878/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1664 _5949_/X VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6417__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1675 _7574_/Q VGND VGND VPWR VPWR hold99/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1686 _3848_/A2 VGND VGND VPWR VPWR _5749_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1697 hold381/X VGND VGND VPWR VPWR _5985_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6136__C _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5748__S _5748_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6718__A1 _7184_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6194__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3952__A1 _7391_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3792__A _3792_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_31_csclk_A clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__A1 _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4400__B _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4879__B_N _4887_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6654__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4128__A _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4968__B1 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6709__A1 _7134_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3640__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4196__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2188_A _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5570_ _4996_/A _5038_/B _5425_/X _5189_/X VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__a31o_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3943__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4521_ _4551_/B _4521_/B _4533_/B VGND VGND VPWR VPWR _4526_/S sky130_fd_sc_hd__and3_2
XFILLER_172_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold205 hold205/A VGND VGND VPWR VPWR _7499_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7240_ _7327_/CLK _7240_/D fanout703/X VGND VGND VPWR VPWR _7240_/Q sky130_fd_sc_hd__dfstp_4
Xhold216 hold216/A VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6488__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4452_ _4452_/A0 _5914_/A1 _4454_/S VGND VGND VPWR VPWR _4452_/X sky130_fd_sc_hd__mux2_1
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold238 hold238/A VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5696__A1 hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold249 _3485_/C VGND VGND VPWR VPWR _3511_/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_3403_ _7075_/Q VGND VGND VPWR VPWR _3403_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4948__D _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7171_ _7181_/CLK _7171_/D fanout724/X VGND VGND VPWR VPWR _7171_/Q sky130_fd_sc_hd__dfrtp_2
X_4383_ _5582_/A0 _4383_/A1 _4387_/S VGND VGND VPWR VPWR _4383_/X sky130_fd_sc_hd__mux2_1
Xfanout707 fanout709/X VGND VGND VPWR VPWR fanout707/X sky130_fd_sc_hd__buf_8
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6122_/A _6122_/B VGND VGND VPWR VPWR _6122_/Y sky130_fd_sc_hd__nand2_8
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout718 fanout719/X VGND VGND VPWR VPWR fanout718/X sky130_fd_sc_hd__buf_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout729 fanout730/X VGND VGND VPWR VPWR fanout729/X sky130_fd_sc_hd__buf_8
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6052_/X _6019_/A _6050_/Y _6019_/Y _6441_/D VGND VGND VPWR VPWR _7596_/D
+ sky130_fd_sc_hd__a32o_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5004_/A1 _5089_/B _4675_/A _4675_/B _4675_/C VGND VGND VPWR VPWR _5005_/C
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA_hold2891_A _7498_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _7578_/CLK hold86/X fanout747/X VGND VGND VPWR VPWR _6955_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5620__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5906_ _5978_/A0 _5906_/A1 hold42/A VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__mux2_1
X_6886_ _4169_/B2 _6886_/D _6836_/X VGND VGND VPWR VPWR _6886_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3631__B1 _3553_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5837_ _5837_/A0 _5999_/A1 _5838_/S VGND VGND VPWR VPWR _5837_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__A2 _3444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout605_A _3444_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5768_ _5768_/A0 _5993_/A1 _5775_/S VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__mux2_1
X_7507_ _7531_/CLK _7507_/D fanout743/X VGND VGND VPWR VPWR _7507_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3934__A1 _4175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4719_ _4786_/D _4909_/D _4772_/B _4767_/A VGND VGND VPWR VPWR _5387_/D sky130_fd_sc_hd__and4bb_4
XFILLER_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5699_ _5699_/A0 _5951_/A1 _5703_/S VGND VGND VPWR VPWR _5699_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7438_ _7579_/CLK hold36/X fanout731/X VGND VGND VPWR VPWR _7438_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold750 hold750/A VGND VGND VPWR VPWR _7070_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7369_ _7542_/CLK _7369_/D fanout719/X VGND VGND VPWR VPWR _7369_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold761 hold761/A VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold772 hold772/A VGND VGND VPWR VPWR _7285_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold794 _5598_/X VGND VGND VPWR VPWR _7230_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6636__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2140 _7534_/Q VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2151 _7550_/Q VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2162 _7462_/Q VGND VGND VPWR VPWR hold62/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4111__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2173 _4249_/X VGND VGND VPWR VPWR hold482/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_input138_A wb_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2184 hold595/X VGND VGND VPWR VPWR _5806_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1450 _4191_/X VGND VGND VPWR VPWR _4202_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2195 _5748_/X VGND VGND VPWR VPWR hold245/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1461 hold140/X VGND VGND VPWR VPWR _4256_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1472 hold187/X VGND VGND VPWR VPWR _7556_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1483 hold65/X VGND VGND VPWR VPWR _7453_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1494 hold19/X VGND VGND VPWR VPWR hold1494/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3870__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3003_A _7257_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5611__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4965__A3 _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5678__A1 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_798 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4350__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6627__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3461__S _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6642__A3 _6428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6057__B _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6740_ _7059_/Q _6447_/C _6769_/A3 _6435_/X _7049_/Q VGND VGND VPWR VPWR _6740_/X
+ sky130_fd_sc_hd__a32o_1
X_3952_ _7391_/Q _5740_/A _5785_/B _3951_/X VGND VGND VPWR VPWR _3952_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3613__B1 _5920_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6671_ _7157_/Q _6419_/A _6670_/X _6430_/X VGND VGND VPWR VPWR _6671_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6158__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3883_ _7123_/Q _5740_/A _4551_/A _4515_/B _3882_/X VGND VGND VPWR VPWR _3883_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_176_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5622_ _3933_/Y _5732_/A1 _5622_/B1 _5640_/D VGND VGND VPWR VPWR _5622_/X sky130_fd_sc_hd__o211a_1
XFILLER_136_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5553_ _5216_/A _5339_/C _5328_/X _5552_/X _5015_/X VGND VGND VPWR VPWR _5554_/C
+ sky130_fd_sc_hd__a311oi_1
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _4504_/A0 _5582_/A0 _4508_/S VGND VGND VPWR VPWR _4504_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3863__C _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5484_ _5484_/A1 _5580_/A2 _5482_/Y _5560_/B _5464_/Y VGND VGND VPWR VPWR _7205_/D
+ sky130_fd_sc_hd__a221o_1
X_7223_ _7232_/CLK _7223_/D _4128_/B VGND VGND VPWR VPWR _7223_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_105_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4435_ _4435_/A0 _5978_/A0 _4439_/S VGND VGND VPWR VPWR _4435_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5851__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout504 _6022_/X VGND VGND VPWR VPWR _6384_/A4 sky130_fd_sc_hd__buf_4
X_7154_ _7185_/CLK _7154_/D fanout725/X VGND VGND VPWR VPWR _7154_/Q sky130_fd_sc_hd__dfstp_4
X_4366_ _4366_/A0 hold198/X _4369_/S VGND VGND VPWR VPWR _4366_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6618__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout526 _4703_/Y VGND VGND VPWR VPWR _5480_/A1 sky130_fd_sc_hd__buf_6
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6105_ _7303_/Q _6121_/A _6121_/B _6071_/X _7287_/Q VGND VGND VPWR VPWR _6105_/X
+ sky130_fd_sc_hd__a32o_1
Xfanout548 _4446_/A1 VGND VGND VPWR VPWR hold1428/A sky130_fd_sc_hd__buf_6
X_7085_ _7514_/CLK _7085_/D fanout743/X VGND VGND VPWR VPWR _7664_/A sky130_fd_sc_hd__dfrtp_1
Xfanout559 _5726_/A1 VGND VGND VPWR VPWR _5625_/A1 sky130_fd_sc_hd__buf_8
X_4297_ _4302_/S _3795_/B _4296_/Y VGND VGND VPWR VPWR _6983_/D sky130_fd_sc_hd__o21ai_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6116_/C _6121_/B _6121_/C VGND VGND VPWR VPWR _6036_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__6633__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ _7575_/CLK _6938_/D fanout735/X VGND VGND VPWR VPWR _6938_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6414__C _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6869_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6869_/X sky130_fd_sc_hd__and2_1
XANTENNA__6149__A2 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__7095__RESET_B fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__A1 _7408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__B2 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5761__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6321__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4332__A1 _5625_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 hold580/A VGND VGND VPWR VPWR _7241_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold591 hold591/A VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6609__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5832__A1 _5985_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1280 hold3239/X VGND VGND VPWR VPWR _6988_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3989__A4 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1291 hold3247/X VGND VGND VPWR VPWR hold3248/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5936__S _5937_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3610__A3 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6560__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_173_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6312__A2 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4220_ _4220_/A0 _4219_/X _4232_/S VGND VGND VPWR VPWR _4220_/X sky130_fd_sc_hd__mux2_1
Xhold2909 _4542_/X VGND VGND VPWR VPWR hold2909/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3677__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4151_ _6933_/Q _4168_/D _6899_/Q VGND VGND VPWR VPWR _4151_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4287__S _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6076__A1 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4082_ _6894_/Q _4082_/A2 _7073_/Q _4123_/B VGND VGND VPWR VPWR _6879_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5823__A1 _5994_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6379__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4984_ _4984_/A _4984_/B _4984_/C VGND VGND VPWR VPWR _5216_/C sky130_fd_sc_hd__and3_1
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6723_ _7144_/Q _6468_/X _6719_/X _6720_/X _6722_/X VGND VGND VPWR VPWR _6723_/X
+ sky130_fd_sc_hd__a2111o_1
X_3935_ input52/X _4431_/A _4479_/A _5974_/A _7559_/Q VGND VGND VPWR VPWR _3935_/X
+ sky130_fd_sc_hd__a32o_1
X_6654_ _7051_/Q _6434_/X _6466_/X _7209_/Q _6653_/X VGND VGND VPWR VPWR _6654_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3866_ input53/X _4431_/A _5992_/C _3549_/X input44/X VGND VGND VPWR VPWR _3866_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_176_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6000__A1 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5605_ _5605_/A0 _5645_/A0 _5611_/S VGND VGND VPWR VPWR _5605_/X sky130_fd_sc_hd__mux2_1
X_6585_ _7316_/Q _6419_/D _6424_/X _7572_/Q _6584_/X VGND VGND VPWR VPWR _6585_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5354__A3 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3797_ _3797_/A1 _3996_/A _3795_/Y _3796_/X VGND VGND VPWR VPWR _3797_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6551__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5536_ _4997_/A _5404_/D _5297_/B _5410_/A VGND VGND VPWR VPWR _5536_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5467_ _5467_/A _5467_/B _5467_/C VGND VGND VPWR VPWR _5521_/B sky130_fd_sc_hd__and3_2
XANTENNA__5106__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4314__A1 _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7206_ _7633_/CLK _7206_/D _6780_/B VGND VGND VPWR VPWR _7206_/Q sky130_fd_sc_hd__dfrtp_1
X_4418_ _4446_/A0 _4446_/A1 _4422_/S VGND VGND VPWR VPWR _4418_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5398_ _5480_/B2 _4748_/Y _5528_/A3 _4832_/Y _4826_/Y VGND VGND VPWR VPWR _5482_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_160_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7137_ _7197_/CLK _7137_/D fanout741/X VGND VGND VPWR VPWR _7137_/Q sky130_fd_sc_hd__dfrtp_4
X_4349_ _4349_/A0 _5815_/A1 _4351_/S VGND VGND VPWR VPWR _4349_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout672_A _5134_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout356 _6068_/Y VGND VGND VPWR VPWR _6777_/S sky130_fd_sc_hd__buf_8
XANTENNA__6409__C _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout367 hold31/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__buf_8
X_7068_ _7268_/CLK _7068_/D _6869_/A VGND VGND VPWR VPWR _7068_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_74_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout389 _3548_/X VGND VGND VPWR VPWR _3738_/B sky130_fd_sc_hd__buf_4
XANTENNA__5814__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6019_ _6019_/A _6929_/Q VGND VGND VPWR VPWR _6019_/Y sky130_fd_sc_hd__nor2_8
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold250_A _3563_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4871__A_N _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6425__B _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4871__D _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4101__A_N _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4250__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1954_A _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6542__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input66_A mgmt_gpio_in[37] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4305__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_151_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4608__A2 _4747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5805__A1 hold198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6230__B2 _7452_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _3470_/X _3485_/X _4509_/C _3669_/X _6971_/Q VGND VGND VPWR VPWR _3720_/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA__3595__A2 _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3651_ _5830_/C _5938_/C _4388_/B VGND VGND VPWR VPWR _3651_/X sky130_fd_sc_hd__and3_2
Xclkbuf_4_0__f_wb_clk_i clkbuf_3_0_0_wb_clk_i/X VGND VGND VPWR VPWR _7601_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6533__A2 _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6370_ _6367_/X _6368_/X _6369_/X _6082_/C VGND VGND VPWR VPWR _6370_/X sky130_fd_sc_hd__o31a_1
XANTENNA_hold2268_A _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3582_ _7381_/Q _3498_/X _3564_/X _7365_/Q _3581_/X VGND VGND VPWR VPWR _3587_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3898__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5321_ _4595_/Y _4601_/Y _4622_/Y _4846_/Y _4956_/B VGND VGND VPWR VPWR _5321_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_170_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6297__B2 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5252_ _5252_/A _5252_/B _5252_/C VGND VGND VPWR VPWR _5252_/Y sky130_fd_sc_hd__nor3_1
XFILLER_88_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2706 _7225_/Q VGND VGND VPWR VPWR hold757/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4203_ _5640_/B _5619_/A _5596_/A _5640_/D VGND VGND VPWR VPWR _4203_/X sky130_fd_sc_hd__and4_1
XFILLER_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2717 hold981/X VGND VGND VPWR VPWR _5833_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3860__D _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5183_ _5183_/A _5183_/B _5183_/C _5339_/D VGND VGND VPWR VPWR _5183_/Y sky130_fd_sc_hd__nand4_1
Xhold2728 hold775/X VGND VGND VPWR VPWR _4363_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2739 _7223_/Q VGND VGND VPWR VPWR hold765/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4134_ _6897_/Q _4134_/B VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__and2b_4
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4065_ _4062_/B _4098_/A1 _6891_/Q _4062_/Y VGND VGND VPWR VPWR _4065_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__3807__B1 _3531_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3822__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4967_ _4966_/X _4965_/X _4964_/Y _4854_/X VGND VGND VPWR VPWR _4967_/Y sky130_fd_sc_hd__o31ai_4
XANTENNA__6772__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3586__A2 _3506_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6706_ _7013_/Q _6423_/X _6462_/X _7033_/Q _6705_/X VGND VGND VPWR VPWR _6706_/X
+ sky130_fd_sc_hd__a221o_1
X_3918_ input96/X _3933_/A _4265_/B _3916_/X _3917_/X VGND VGND VPWR VPWR _3918_/X
+ sky130_fd_sc_hd__a311o_1
X_4898_ _5005_/A _4948_/B _4898_/C _5222_/B VGND VGND VPWR VPWR _4898_/Y sky130_fd_sc_hd__nand4_4
XANTENNA_fanout518_A _4983_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6637_ _7302_/Q _6420_/A _6632_/X _6634_/X _6636_/X VGND VGND VPWR VPWR _6647_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_20_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3849_ input45/X _3549_/X _3846_/X _3847_/X _3848_/X VGND VGND VPWR VPWR _3849_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__6524__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6568_ _7547_/Q _6419_/A _6435_/X _7515_/Q _6567_/X VGND VGND VPWR VPWR _6569_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4212__C _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3889__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5519_ _4717_/Y _4722_/Y _5083_/X _4718_/Y VGND VGND VPWR VPWR _5521_/D sky130_fd_sc_hd__o211a_1
X_6499_ _7489_/Q _6463_/A _6441_/X _6425_/X _7337_/Q VGND VGND VPWR VPWR _6499_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6288__A1 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold1702_A _7513_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3510__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5799__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__7457__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input120_A wb_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3813__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3498__C _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6515__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4526__A1 _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6279__A1 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _5870_/A0 _5978_/A0 _5871_/S VGND VGND VPWR VPWR _5870_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5006__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6203__A1 _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4821_ _5058_/D _4856_/A _5072_/B VGND VGND VPWR VPWR _4821_/Y sky130_fd_sc_hd__nand3_4
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6754__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7540_ _7541_/CLK _7540_/D fanout713/X VGND VGND VPWR VPWR _7540_/Q sky130_fd_sc_hd__dfrtp_4
X_4752_ _4706_/Y _4741_/Y _4751_/Y _4687_/Y _4746_/Y VGND VGND VPWR VPWR _4760_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3703_ _7387_/Q _5776_/A _3658_/X _7116_/Q VGND VGND VPWR VPWR _3703_/X sky130_fd_sc_hd__a22o_1
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7471_ _7471_/CLK _7471_/D fanout729/X VGND VGND VPWR VPWR _7471_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_146_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4683_ _4562_/Y _4585_/Y _4687_/C VGND VGND VPWR VPWR _5138_/A sky130_fd_sc_hd__o21a_4
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6506__A2 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5714__A0 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6422_ _6467_/A _6468_/C _6651_/B VGND VGND VPWR VPWR _6422_/X sky130_fd_sc_hd__and3_4
XANTENNA__4517__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3634_ _7500_/Q hold41/A _3526_/X _7508_/Q _3633_/X VGND VGND VPWR VPWR _3642_/A
+ sky130_fd_sc_hd__a221o_1
X_6353_ _6959_/Q _6036_/Y _6341_/X _6352_/X _6067_/A VGND VGND VPWR VPWR _6353_/X
+ sky130_fd_sc_hd__o221a_1
X_3565_ hold40/A hold32/A _5938_/B VGND VGND VPWR VPWR _3565_/X sky130_fd_sc_hd__and3_4
XFILLER_143_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5304_ _4667_/A _4692_/Y _4712_/Y _4716_/Y _4755_/Y VGND VGND VPWR VPWR _5304_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_115_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3740__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6284_ _6283_/X _6284_/A1 _6777_/S VGND VGND VPWR VPWR _6284_/X sky130_fd_sc_hd__mux2_1
Xhold3204 hold3204/A VGND VGND VPWR VPWR _4260_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3215 _4528_/X VGND VGND VPWR VPWR hold3215/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3496_ _3511_/A _3496_/B VGND VGND VPWR VPWR _3496_/Y sky130_fd_sc_hd__nor2_2
Xhold3226 _6927_/Q VGND VGND VPWR VPWR hold3226/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3237 _6988_/Q VGND VGND VPWR VPWR hold3237/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _5235_/A _5444_/D _5235_/C VGND VGND VPWR VPWR _5237_/B sky130_fd_sc_hd__and3_1
Xhold3248 hold3248/A VGND VGND VPWR VPWR _5714_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2503 _5745_/X VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3259 _6911_/Q VGND VGND VPWR VPWR hold3259/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2514 hold955/X VGND VGND VPWR VPWR _5827_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2525 hold659/X VGND VGND VPWR VPWR _5648_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2536 _5764_/X VGND VGND VPWR VPWR hold932/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1802 _3500_/X VGND VGND VPWR VPWR hold1802/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2547 _7402_/Q VGND VGND VPWR VPWR hold911/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1813 hold29/X VGND VGND VPWR VPWR _3458_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__B2 _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5166_ wire375/X _5166_/A2 _5203_/C _5060_/A VGND VGND VPWR VPWR _5496_/B sky130_fd_sc_hd__a31oi_4
XFILLER_69_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2558 _7017_/Q VGND VGND VPWR VPWR hold921/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1824 _5688_/X VGND VGND VPWR VPWR hold352/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2569 hold935/X VGND VGND VPWR VPWR _4378_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1835 hold433/X VGND VGND VPWR VPWR _5850_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4117_ _6009_/B _4117_/B VGND VGND VPWR VPWR _4117_/Y sky130_fd_sc_hd__nand2_2
Xhold1846 hold267/X VGND VGND VPWR VPWR _4404_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1857 _7440_/Q VGND VGND VPWR VPWR hold447/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1868 _7145_/Q VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5097_ _5097_/A _5097_/B _5444_/B VGND VGND VPWR VPWR _5097_/Y sky130_fd_sc_hd__nand3_1
Xhold1879 _4344_/X VGND VGND VPWR VPWR hold321/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6442__B2 _7287_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4048_ _4062_/A _3998_/Y _3403_/Y _4113_/B1 _4048_/B1 VGND VGND VPWR VPWR _4048_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5650__C1 _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout635_A _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5999_ _5999_/A0 _5999_/A1 _6000_/S VGND VGND VPWR VPWR _5999_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6745__A2 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3559__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7669_ _7669_/A VGND VGND VPWR VPWR _7669_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5705__A0 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5038__C _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3731__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input168_A wb_sel_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6130__B1 _6276_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput290 _6924_/Q VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3495__A1 _7414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4893__B _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4385__S _4387_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input29_A mask_rev_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3798__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6197__B1 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6736__A2 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6332__C _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6051__D _6434_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire351 _6631_/Y VGND VGND VPWR VPWR wire351/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3970__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5325__A2_N _4977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7539_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold409 hold409/A VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5172__B2 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5024_/A1 _4669_/X _4974_/B _5404_/D _5180_/A VGND VGND VPWR VPWR _5021_/D
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__5475__A2 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1109 hold3132/X VGND VGND VPWR VPWR hold3133/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6971_ _7176_/CLK _6971_/D fanout722/X VGND VGND VPWR VPWR _6971_/Q sky130_fd_sc_hd__dfrtp_4
X_5922_ _5922_/A0 _5922_/A1 _5928_/S VGND VGND VPWR VPWR _5922_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3789__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5853_ _5853_/A0 _5853_/A1 _5856_/S VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6188__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7035_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5935__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4804_ _4700_/Y _4798_/Y _4803_/Y _4800_/Y VGND VGND VPWR VPWR _4809_/C sky130_fd_sc_hd__o211ai_1
X_5784_ hold20/X _5784_/A1 _5784_/S VGND VGND VPWR VPWR _5784_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4735_ _5404_/B _5404_/C VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__nand2_1
X_7523_ _7561_/CLK _7523_/D fanout738/X VGND VGND VPWR VPWR _7523_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5854__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2934_A _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7454_ _7573_/CLK hold23/X fanout733/X VGND VGND VPWR VPWR _7454_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _4860_/A _4831_/A VGND VGND VPWR VPWR _4667_/C sky130_fd_sc_hd__nand2b_2
XANTENNA__4978__B _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6405_ _6466_/A _6466_/B _6466_/C _6462_/C VGND VGND VPWR VPWR _6408_/B sky130_fd_sc_hd__and4_4
X_3617_ _5596_/A _5596_/B _5659_/B VGND VGND VPWR VPWR _3617_/X sky130_fd_sc_hd__and3_4
Xhold910 hold910/A VGND VGND VPWR VPWR _7341_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7385_ _7421_/CLK _7385_/D fanout716/X VGND VGND VPWR VPWR _7385_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6360__B1 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold921 hold921/A VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4597_ _4910_/D _4856_/A VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__4697__C _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap640 _4082_/A2 VGND VGND VPWR VPWR _4085_/A2 sky130_fd_sc_hd__buf_4
Xhold932 hold932/A VGND VGND VPWR VPWR _7372_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold943 hold943/A VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold954 hold954/A VGND VGND VPWR VPWR _7044_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3713__A2 hold90/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6336_ _6969_/Q _6136_/B _6121_/B _6332_/C _7033_/Q VGND VGND VPWR VPWR _6336_/X
+ sky130_fd_sc_hd__a32o_1
X_3548_ _4551_/A _3576_/B _3576_/C VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__and3_2
Xhold965 hold965/A VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3001 _6981_/Q VGND VGND VPWR VPWR _4293_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold976 _5791_/X VGND VGND VPWR VPWR _7396_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3012 hold3012/A VGND VGND VPWR VPWR hold3012/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold987 hold987/A VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold998 hold998/A VGND VGND VPWR VPWR _6937_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3023 hold3023/A VGND VGND VPWR VPWR hold3023/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4994__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6267_ _7454_/Q _6144_/A _6116_/A _6267_/B1 _7526_/Q VGND VGND VPWR VPWR _6267_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3034 _5777_/X VGND VGND VPWR VPWR hold3034/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout585_A _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3479_ _7398_/Q _5803_/A _4431_/A _5848_/A _7454_/Q VGND VGND VPWR VPWR _3479_/X
+ sky130_fd_sc_hd__a32o_4
Xhold2300 hold667/X VGND VGND VPWR VPWR _4254_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3045 hold3045/A VGND VGND VPWR VPWR _5786_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2311 _4243_/X VGND VGND VPWR VPWR hold574/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3056 hold3056/A VGND VGND VPWR VPWR _5831_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5466__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2322 hold553/X VGND VGND VPWR VPWR _5595_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3067 _7295_/Q VGND VGND VPWR VPWR hold3067/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5218_ _5079_/X _5216_/X _5065_/A VGND VGND VPWR VPWR _5218_/Y sky130_fd_sc_hd__o21ai_1
Xhold2333 hold717/X VGND VGND VPWR VPWR _5707_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3078 hold3078/A VGND VGND VPWR VPWR _5615_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3089 hold3089/A VGND VGND VPWR VPWR _4409_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2344 _7403_/Q VGND VGND VPWR VPWR hold567/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6198_ _6082_/C _6089_/X _7379_/Q _6119_/X _7403_/Q VGND VGND VPWR VPWR _6198_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2355 _5719_/X VGND VGND VPWR VPWR hold796/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1610 _5627_/X VGND VGND VPWR VPWR hold167/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2366 _5953_/X VGND VGND VPWR VPWR hold798/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1621 _7328_/Q VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1632 hold47/X VGND VGND VPWR VPWR _5767_/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2377 _7146_/Q VGND VGND VPWR VPWR hold679/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5149_ _4687_/Y _4777_/X _4821_/Y _4698_/Y _4723_/Y VGND VGND VPWR VPWR _5150_/C
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout752_A input164/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2388 _4384_/X VGND VGND VPWR VPWR hold806/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1643 _7260_/Q VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1654 hold313/X VGND VGND VPWR VPWR _7270_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2399 _7057_/Q VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1665 _7320_/Q VGND VGND VPWR VPWR hold369/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1676 hold99/X VGND VGND VPWR VPWR _5991_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1687 _5679_/X VGND VGND VPWR VPWR hold376/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1698 _5985_/X VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6179__B1 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6718__A2 _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5764__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3952__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5154__A1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold3150_A _7503_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4901__A1 _4726_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3704__A2 _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4400__C _5596_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3468__A1 _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7401__RESET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output302_A _3619_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6709__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6185__A3 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6590__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4520_ _4520_/A0 _5817_/A1 _4520_/S VGND VGND VPWR VPWR _4520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3943__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_722 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ _4451_/A0 _4553_/A0 _4454_/S VGND VGND VPWR VPWR _4451_/X sky130_fd_sc_hd__mux2_1
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold217 hold217/A VGND VGND VPWR VPWR _7513_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6342__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold2250_A _7233_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold239 hold239/A VGND VGND VPWR VPWR _7309_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3402_ _4058_/A VGND VGND VPWR VPWR _4062_/A sky130_fd_sc_hd__inv_4
X_7170_ _7213_/CLK _7170_/D fanout701/X VGND VGND VPWR VPWR _7170_/Q sky130_fd_sc_hd__dfrtp_2
X_4382_ _4551_/A _4551_/B _4455_/C _4533_/B VGND VGND VPWR VPWR _4387_/S sky130_fd_sc_hd__nand4_4
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ _6121_/A _6121_/B _6121_/C VGND VGND VPWR VPWR _6121_/X sky130_fd_sc_hd__and3_4
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout708 fanout709/X VGND VGND VPWR VPWR fanout708/X sky130_fd_sc_hd__buf_8
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout719 fanout720/X VGND VGND VPWR VPWR fanout719/X sky130_fd_sc_hd__clkbuf_16
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _7594_/Q _6429_/C _6433_/D _6441_/D VGND VGND VPWR VPWR _6052_/X sky130_fd_sc_hd__a31o_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _4675_/A _4675_/B _4675_/C _4591_/B VGND VGND VPWR VPWR _5005_/B sky130_fd_sc_hd__a31o_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5849__S _5856_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2884_A _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4959__B2 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6954_ _7575_/CLK _6954_/D fanout735/X VGND VGND VPWR VPWR _6954_/Q sky130_fd_sc_hd__dfrtp_1
X_5905_ _5950_/A1 _5905_/A1 hold42/X VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3631__A1 _4173_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6885_ _4169_/B2 _6885_/D _6835_/X VGND VGND VPWR VPWR _6885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3631__B2 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5908__A0 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5836_ _5836_/A0 _5998_/A1 _5838_/S VGND VGND VPWR VPWR _5836_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6176__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4989__A _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5767_ _5767_/A _5983_/A _5992_/D VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__and3_4
XANTENNA__6581__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_148_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7506_ _7565_/CLK _7506_/D fanout743/X VGND VGND VPWR VPWR _7506_/Q sky130_fd_sc_hd__dfrtp_4
X_4718_ _4803_/A _4765_/B VGND VGND VPWR VPWR _4718_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3934__A2 _3552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5698_ _5698_/A0 _5968_/A1 _5703_/S VGND VGND VPWR VPWR _5698_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5136__A1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4649_ _4591_/Y _4616_/Y _4675_/A _4675_/B VGND VGND VPWR VPWR _4726_/C sky130_fd_sc_hd__nand4bb_4
XANTENNA__6333__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7437_ _7576_/CLK _7437_/D fanout717/X VGND VGND VPWR VPWR _7437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold740 hold740/A VGND VGND VPWR VPWR _7126_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7368_ _7472_/CLK _7368_/D fanout719/X VGND VGND VPWR VPWR _7368_/Q sky130_fd_sc_hd__dfstp_1
Xhold751 hold751/A VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold762 hold762/A VGND VGND VPWR VPWR _7236_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold773 hold773/A VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold784 hold784/A VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6319_ _7183_/Q _6097_/X _6317_/X _6318_/X _6316_/X VGND VGND VPWR VPWR _6327_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold795 hold795/A VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7299_ _7329_/CLK _7299_/D fanout704/X VGND VGND VPWR VPWR _7299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6636__B2 _7510_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2130 _5910_/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2141 hold66/X VGND VGND VPWR VPWR _5946_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2152 hold60/X VGND VGND VPWR VPWR _5964_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2163 hold62/X VGND VGND VPWR VPWR _5865_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2174 hold482/X VGND VGND VPWR VPWR _6948_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1440 hold10/X VGND VGND VPWR VPWR _4447_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2185 _5806_/X VGND VGND VPWR VPWR hold596/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1451 _4198_/X VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2196 _7345_/Q VGND VGND VPWR VPWR hold637/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1462 _4256_/X VGND VGND VPWR VPWR hold141/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1473 _7485_/Q VGND VGND VPWR VPWR hold1473/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1484 _7662_/A VGND VGND VPWR VPWR hold70/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__A1 _7138_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1495 _4422_/A1 VGND VGND VPWR VPWR _5991_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__B2 _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5759__S hold27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4890__C _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3622__A1 _7234_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input96_A usr1_vdd_pwrgood VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5375__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6572__B1 _6570_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6324__B1 _6094_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _7152_/Q _5740_/A _4352_/B _3661_/X _7031_/Q VGND VGND VPWR VPWR _3951_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3613__A1 _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3613__B2 _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6670_ _7142_/Q _6468_/X _6667_/X _6669_/X VGND VGND VPWR VPWR _6670_/X sky130_fd_sc_hd__a211o_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3882_ _7352_/Q _4473_/A _5956_/B _4370_/A _7042_/Q VGND VGND VPWR VPWR _3882_/X
+ sky130_fd_sc_hd__a32o_1
X_5621_ _5612_/A _5590_/A _5619_/A _5621_/B1 VGND VGND VPWR VPWR _5621_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5366__A1 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6563__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3916__A2 _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5552_ _5180_/B _5342_/B _5013_/C _5339_/A VGND VGND VPWR VPWR _5552_/X sky130_fd_sc_hd__o211a_1
X_4503_ _4539_/C _5632_/B _5619_/C VGND VGND VPWR VPWR _4508_/S sky130_fd_sc_hd__and3_4
XANTENNA__3863__D _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6315__B1 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5483_ _5073_/A _5495_/C1 _4826_/Y _5374_/X _7107_/Q VGND VGND VPWR VPWR _5560_/B
+ sky130_fd_sc_hd__o311a_1
X_4434_ _4434_/A0 _5986_/A1 _4439_/S VGND VGND VPWR VPWR _4434_/X sky130_fd_sc_hd__mux2_1
X_7222_ _7255_/CLK _7222_/D _4128_/B VGND VGND VPWR VPWR _7222_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_144_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7153_ _7185_/CLK _7153_/D fanout737/X VGND VGND VPWR VPWR _7153_/Q sky130_fd_sc_hd__dfrtp_4
X_4365_ _4365_/A0 _5582_/A0 _4369_/S VGND VGND VPWR VPWR _4365_/X sky130_fd_sc_hd__mux2_1
Xfanout505 _6112_/B VGND VGND VPWR VPWR _6144_/A sky130_fd_sc_hd__buf_8
X_6104_ _7327_/Q _6079_/X _6091_/X _7399_/Q _6103_/X VGND VGND VPWR VPWR _6104_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout538 _6000_/A1 VGND VGND VPWR VPWR _5955_/A1 sky130_fd_sc_hd__buf_8
XFILLER_58_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7084_ _7646_/CLK _7084_/D fanout751/X VGND VGND VPWR VPWR _7084_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout549 _4446_/A1 VGND VGND VPWR VPWR _5998_/A1 sky130_fd_sc_hd__buf_6
X_4296_ _4302_/S _4296_/B VGND VGND VPWR VPWR _4296_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6035_ _6099_/D _6081_/C VGND VGND VPWR VPWR _6035_/Y sky130_fd_sc_hd__nor2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout548_A _4446_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ _7551_/CLK _6937_/D fanout734/X VGND VGND VPWR VPWR _7655_/A sky130_fd_sc_hd__dfrtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_74_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6868_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6868_/X sky130_fd_sc_hd__and2_1
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5819_ _5819_/A0 _5999_/A1 _5820_/S VGND VGND VPWR VPWR _5819_/X sky130_fd_sc_hd__mux2_1
X_6799_ _4427_/D _6799_/A2 _6799_/B1 _4427_/C VGND VGND VPWR VPWR _6799_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold570 _5685_/X VGND VGND VPWR VPWR _7302_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold581 hold581/A VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold592 hold592/A VGND VGND VPWR VPWR _7435_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input150_A wb_dat_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5293__B1 _4428_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1270 _4367_/X VGND VGND VPWR VPWR _7038_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3843__A1 _7481_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input11_A mask_rev_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3843__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1281 hold3221/X VGND VGND VPWR VPWR hold3222/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1292 hold3249/X VGND VGND VPWR VPWR _7327_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5348__A1 _5094_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4795__C _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4150_ _6934_/Q _4150_/A1 _6898_/Q VGND VGND VPWR VPWR _4150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6783__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4081_ _4076_/B _4050_/S _4080_/X _4121_/A VGND VGND VPWR VPWR _6880_/D sky130_fd_sc_hd__a22o_1
XFILLER_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3501__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _5038_/A _5183_/A _4983_/C VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__and3_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6722_ _7124_/Q _6420_/C _6467_/X _7154_/Q _6721_/X VGND VGND VPWR VPWR _6722_/X
+ sky130_fd_sc_hd__a221o_1
X_3934_ _4175_/A _3552_/X _3652_/X _7147_/Q VGND VGND VPWR VPWR _3934_/X sky130_fd_sc_hd__a22o_1
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3865_ _7223_/Q _5612_/A _5640_/A _5619_/A VGND VGND VPWR VPWR _3865_/X sky130_fd_sc_hd__and4_2
X_6653_ _7046_/Q _6435_/X _6443_/X _7192_/Q _6652_/X VGND VGND VPWR VPWR _6653_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6536__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5604_ _5604_/A0 _5948_/A1 _5611_/S VGND VGND VPWR VPWR _5604_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2847_A _7303_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3796_ _7216_/Q _3856_/A _7073_/Q _6893_/Q VGND VGND VPWR VPWR _3796_/X sky130_fd_sc_hd__o211a_1
X_6584_ _7593_/Q _7580_/Q _6408_/C _6583_/X VGND VGND VPWR VPWR _6584_/X sky130_fd_sc_hd__a31o_1
XFILLER_145_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5535_ _5535_/A _5535_/B _5535_/C VGND VGND VPWR VPWR _5539_/B sky130_fd_sc_hd__and3_1
XFILLER_191_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5862__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5466_ _5480_/B2 _4722_/Y _4720_/Y _5563_/A1 VGND VGND VPWR VPWR _5467_/C sky130_fd_sc_hd__a211o_1
XFILLER_105_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4417_ _4417_/A0 _4416_/X _4423_/S VGND VGND VPWR VPWR _4417_/X sky130_fd_sc_hd__mux2_1
X_7205_ _7633_/CLK _7205_/D _6780_/B VGND VGND VPWR VPWR _7205_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4314__A2 _3856_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5397_ _4668_/C _4827_/X _5110_/X _5396_/X VGND VGND VPWR VPWR _5397_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout498_A _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3522__B1 _3521_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4348_ _4348_/A0 _5645_/A0 _4351_/S VGND VGND VPWR VPWR _4348_/X sky130_fd_sc_hd__mux2_1
X_7136_ _7176_/CLK _7136_/D fanout724/X VGND VGND VPWR VPWR _7136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout357 _6068_/Y VGND VGND VPWR VPWR _6573_/S sky130_fd_sc_hd__buf_4
XANTENNA_input3_A debug_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7067_ _7191_/CLK _7067_/D _6872_/A VGND VGND VPWR VPWR _7067_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout368 _5866_/B VGND VGND VPWR VPWR _4551_/B sky130_fd_sc_hd__buf_8
Xfanout379 _6869_/B VGND VGND VPWR VPWR _6873_/B sky130_fd_sc_hd__buf_4
X_4279_ _4289_/S _3996_/B _4278_/Y VGND VGND VPWR VPWR _6972_/D sky130_fd_sc_hd__o21ai_1
X_6018_ _6018_/A _6018_/B _6018_/C VGND VGND VPWR VPWR _7587_/D sky130_fd_sc_hd__and3_1
XFILLER_39_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3411__A _7554_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6775__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3589__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6527__B1 _6455_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6542__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5750__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5772__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3761__B1 _3542_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4896__B _4997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input59_A mgmt_gpio_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5502__A1 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3230_A _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3513__B1 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3570__A_N _3491_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3816__B2 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6766__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6230__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_158_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ _4551_/B _4455_/A _4551_/C VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__and3_2
XFILLER_173_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6070__C _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6533__A3 _6428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3581_ _7493_/Q _5947_/B _5965_/B _3549_/X input50/X VGND VGND VPWR VPWR _3581_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5741__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5320_ _4956_/A _4834_/Y _5529_/A _5422_/D _5319_/X VGND VGND VPWR VPWR _5320_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3752__B1 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5251_ _4966_/A _5203_/A _5342_/B _4847_/X VGND VGND VPWR VPWR _5252_/A sky130_fd_sc_hd__a31o_1
XFILLER_142_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4202_ _4202_/A0 _5955_/A1 _4202_/S VGND VGND VPWR VPWR _4202_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2707 hold757/X VGND VGND VPWR VPWR _5592_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5182_ _5034_/C _5018_/B _5180_/X _5181_/X _5179_/Y VGND VGND VPWR VPWR _5185_/A
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2718 _5833_/X VGND VGND VPWR VPWR hold982/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2729 _6958_/Q VGND VGND VPWR VPWR hold743/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4133_ input85/X _4076_/B _6897_/Q VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__mux2_2
XFILLER_29_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4064_ _6891_/Q _4063_/Y _4062_/B _4064_/B1 _4062_/Y VGND VGND VPWR VPWR _4064_/X
+ sky130_fd_sc_hd__o32a_1
X_4966_ _4966_/A _5248_/A _5248_/C VGND VGND VPWR VPWR _4966_/X sky130_fd_sc_hd__and3_1
X_6705_ _7028_/Q _6462_/C _6459_/C _6408_/B _7043_/Q VGND VGND VPWR VPWR _6705_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3917_ input12/X _3490_/X _3542_/X _6920_/Q _3865_/X VGND VGND VPWR VPWR _3917_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__6509__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4897_ _4622_/Y _4956_/A _4726_/Y _4895_/Y VGND VGND VPWR VPWR _4897_/X sky130_fd_sc_hd__o31a_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5158__A _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6636_ _7526_/Q _6446_/X _6466_/X _7510_/Q _6635_/X VGND VGND VPWR VPWR _6636_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout413_A _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ _7226_/Q _3848_/A2 _5659_/B _5713_/A _7329_/Q VGND VGND VPWR VPWR _3848_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_20_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5732__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A _4997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3779_ _7009_/Q _3659_/X _4485_/A _7145_/Q VGND VGND VPWR VPWR _3779_/X sky130_fd_sc_hd__a22o_1
X_6567_ _7499_/Q _6447_/C _6769_/A3 _6455_/X _7459_/Q VGND VGND VPWR VPWR _6567_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3743__B1 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5518_ _5518_/A _5518_/B _5518_/C VGND VGND VPWR VPWR _5562_/C sky130_fd_sc_hd__and3_1
X_6498_ _6497_/X _6522_/A1 _6777_/S VGND VGND VPWR VPWR _6498_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6288__A2 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5449_ _4667_/A _4667_/C _5065_/Y _4913_/B _5228_/D VGND VGND VPWR VPWR _5450_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4299__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7119_ _7561_/CLK _7119_/D fanout741/X VGND VGND VPWR VPWR _7119_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1897_A _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input113_A wb_adr_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _4169_/A2 sky130_fd_sc_hd__clkbuf_16
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4223__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5971__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5723__A1 hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6279__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5006__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6203__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7218__CLK_N _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4820_ _5058_/D _4856_/A _5072_/B VGND VGND VPWR VPWR _5138_/D sky130_fd_sc_hd__and3_4
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4214__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6754__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4751_ _5134_/A _5158_/A _5059_/B _5077_/B _4898_/C VGND VGND VPWR VPWR _4751_/Y
+ sky130_fd_sc_hd__a221oi_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5962__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3702_ _7371_/Q _5758_/A _3698_/X _3699_/X _3701_/X VGND VGND VPWR VPWR _3732_/A
+ sky130_fd_sc_hd__a2111o_2
X_4682_ _4593_/A _4674_/A _5005_/A VGND VGND VPWR VPWR _4687_/C sky130_fd_sc_hd__a21boi_4
X_7470_ _7525_/CLK _7470_/D fanout745/X VGND VGND VPWR VPWR _7470_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6421_ _6455_/B _6467_/A _6462_/C VGND VGND VPWR VPWR _6421_/X sky130_fd_sc_hd__and3_4
X_3633_ _7484_/Q _5938_/C _5956_/B _3520_/X _7444_/Q VGND VGND VPWR VPWR _3633_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_161_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4610__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3564_ _4364_/A _5590_/A _5596_/B VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__and3_4
X_6352_ _7028_/Q _6099_/X _6343_/X _6347_/X _6351_/X VGND VGND VPWR VPWR _6352_/X
+ sky130_fd_sc_hd__a2111o_1
X_5303_ _5303_/A _5538_/A _5405_/D _5303_/D VGND VGND VPWR VPWR _5306_/A sky130_fd_sc_hd__and4_1
X_6283_ _6649_/S _7608_/Q _6281_/X _6282_/X VGND VGND VPWR VPWR _6283_/X sky130_fd_sc_hd__a22o_2
Xhold3205 _7006_/Q VGND VGND VPWR VPWR hold3205/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3495_ _7414_/Q _5803_/A _3590_/C _3494_/X _7478_/Q VGND VGND VPWR VPWR _3495_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3216 _7051_/Q VGND VGND VPWR VPWR hold3216/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3227 hold3227/A VGND VGND VPWR VPWR _4213_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3238 hold3238/A VGND VGND VPWR VPWR _4304_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5234_ _4933_/A _4864_/X _5342_/B _5102_/B _4790_/C VGND VGND VPWR VPWR _5235_/C
+ sky130_fd_sc_hd__a32oi_1
Xhold3249 _5714_/X VGND VGND VPWR VPWR hold3249/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2504 _7027_/Q VGND VGND VPWR VPWR hold917/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2515 _7637_/Q VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2526 _7341_/Q VGND VGND VPWR VPWR hold909/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2537 _7199_/Q VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6690__A2 _6443_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5493__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5165_ _4595_/Y _4748_/Y _4832_/Y _4834_/Y _5480_/B2 VGND VGND VPWR VPWR _5529_/A
+ sky130_fd_sc_hd__o32a_2
Xhold1803 _5614_/X VGND VGND VPWR VPWR _5618_/S sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2548 hold911/X VGND VGND VPWR VPWR _5798_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1814 _3457_/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2559 hold921/X VGND VGND VPWR VPWR _4342_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1825 _7480_/Q VGND VGND VPWR VPWR hold435/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4983__C _4983_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1836 _5850_/X VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4116_ _6009_/B _4117_/B VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__and2_4
XFILLER_69_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1847 _4404_/X VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5096_ _5096_/A _5248_/C VGND VGND VPWR VPWR _5097_/B sky130_fd_sc_hd__nand2_1
Xhold1858 hold447/X VGND VGND VPWR VPWR _5841_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6905__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1869 hold218/X VGND VGND VPWR VPWR _4489_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ _4047_/A0 _4121_/A _4047_/S VGND VGND VPWR VPWR _6899_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6442__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5650__B1 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout530_A _4997_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4205__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _5998_/A0 _5998_/A1 _6000_/S VGND VGND VPWR VPWR _5998_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5953__A1 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3559__A3 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4949_ _4949_/A _4949_/B _4949_/C VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__nor3_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3964__B1 _3537_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7668_ _7668_/A VGND VGND VPWR VPWR _7668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6619_ _7397_/Q _6420_/C _6467_/X _7421_/Q _6600_/X VGND VGND VPWR VPWR _6619_/X
+ sky130_fd_sc_hd__a221o_1
X_7599_ _7627_/CLK _7599_/D fanout690/X VGND VGND VPWR VPWR _7599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3716__B1 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5181__A2 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput280 _6920_/Q VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput291 _6925_/Q VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
XFILLER_160_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4141__B1 _4140_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6681__A2 _6427_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3495__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4444__A1 _5996_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_689 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5944__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3955__B1 _5776_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output282_A _7240_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire352 _6440_/Y VGND VGND VPWR VPWR wire352/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3707__B1 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5172__A2 _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6672__A2 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6791__S _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6970_ _7176_/CLK _6970_/D fanout722/X VGND VGND VPWR VPWR _6970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5921_ _5975_/A0 _5921_/A1 _5928_/S VGND VGND VPWR VPWR _5921_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3789__A3 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5852_ _5978_/A0 _5852_/A1 _5856_/S VGND VGND VPWR VPWR _5852_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6188__A1 _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6188__B2 _7306_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4803_ _4803_/A _4823_/B VGND VGND VPWR VPWR _4803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5783_ _5999_/A1 _5783_/A1 _5784_/S VGND VGND VPWR VPWR _5783_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2662_A _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7522_ _7522_/CLK _7522_/D fanout748/X VGND VGND VPWR VPWR _7522_/Q sky130_fd_sc_hd__dfrtp_4
X_4734_ _4831_/C _4801_/B VGND VGND VPWR VPWR _4734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7453_ _7573_/CLK _7453_/D fanout733/X VGND VGND VPWR VPWR _7453_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4665_ _4767_/A _4786_/D VGND VGND VPWR VPWR _4797_/B sky130_fd_sc_hd__and2b_4
XFILLER_175_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6404_ _7597_/Q _7598_/Q VGND VGND VPWR VPWR _6404_/Y sky130_fd_sc_hd__nor2_1
X_3616_ _7348_/Q _5731_/A _5731_/B VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__and3_1
Xhold900 hold900/A VGND VGND VPWR VPWR _7389_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7384_ _7582_/CLK _7384_/D fanout717/X VGND VGND VPWR VPWR _7384_/Q sky130_fd_sc_hd__dfstp_2
Xhold911 hold911/A VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4596_ _4879_/D _4747_/B VGND VGND VPWR VPWR _4596_/X sky130_fd_sc_hd__and2b_4
XANTENNA__6360__B2 _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold922 hold922/A VGND VGND VPWR VPWR _7017_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap641 _5072_/D VGND VGND VPWR VPWR _5524_/A3 sky130_fd_sc_hd__clkbuf_2
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6335_ _7003_/Q _6116_/C _6120_/B _6317_/C _7114_/Q VGND VGND VPWR VPWR _6335_/X
+ sky130_fd_sc_hd__a32o_1
Xhold944 _5828_/X VGND VGND VPWR VPWR _7429_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3547_ _6926_/Q _3542_/X _5668_/A _7294_/Q _3546_/X VGND VGND VPWR VPWR _3568_/B
+ sky130_fd_sc_hd__a221o_4
Xhold955 hold955/A VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold966 hold966/A VGND VGND VPWR VPWR _7581_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3002 hold3002/A VGND VGND VPWR VPWR hold3002/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_89_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3013 _6974_/Q VGND VGND VPWR VPWR _4281_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3024 _6995_/Q VGND VGND VPWR VPWR _4313_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold988 _4477_/X VGND VGND VPWR VPWR _7135_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6266_ _7398_/Q _6267_/B1 _6075_/A _6265_/X _6263_/X VGND VGND VPWR VPWR _6266_/X
+ sky130_fd_sc_hd__a2111o_1
X_3478_ _4551_/A _5938_/A _5866_/B VGND VGND VPWR VPWR _5848_/A sky130_fd_sc_hd__and3_4
Xhold999 hold999/A VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3035 _7635_/Q VGND VGND VPWR VPWR _6791_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3046 _6972_/Q VGND VGND VPWR VPWR _4278_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2301 _4254_/X VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2312 _7386_/Q VGND VGND VPWR VPWR hold675/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3057 _5831_/X VGND VGND VPWR VPWR hold3057/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2323 _7331_/Q VGND VGND VPWR VPWR hold589/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3068 hold3068/A VGND VGND VPWR VPWR _5678_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_103_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6663__A2 _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5217_ _4907_/B _5342_/B _4940_/D _5079_/X VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__a31o_1
Xhold3079 _7511_/Q VGND VGND VPWR VPWR hold3079/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2334 _5707_/X VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout480_A _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1600 _5932_/X VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6197_ _7411_/Q _6144_/C _6097_/B _6270_/C1 VGND VGND VPWR VPWR _6197_/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout578_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2345 hold567/X VGND VGND VPWR VPWR _5799_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2356 _7246_/Q VGND VGND VPWR VPWR hold741/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1611 _7452_/Q VGND VGND VPWR VPWR hold226/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1622 hold361/X VGND VGND VPWR VPWR _5715_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2367 _7434_/Q VGND VGND VPWR VPWR hold685/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2378 hold679/X VGND VGND VPWR VPWR _4490_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1633 _5767_/X VGND VGND VPWR VPWR _5775_/S sky130_fd_sc_hd__clkdlybuf4s50_2
X_5148_ _5148_/A _5308_/A _5148_/C VGND VGND VPWR VPWR _5150_/B sky130_fd_sc_hd__nor3_1
Xhold2389 _7337_/Q VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1644 hold263/X VGND VGND VPWR VPWR _5637_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1655 _7336_/Q VGND VGND VPWR VPWR hold401/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1666 hold369/X VGND VGND VPWR VPWR _5706_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1677 _5991_/X VGND VGND VPWR VPWR hold100/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5079_ _5100_/A _5079_/B _5248_/C VGND VGND VPWR VPWR _5079_/X sky130_fd_sc_hd__and3_1
Xhold1688 hold376/X VGND VGND VPWR VPWR _7296_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1699 _7666_/A VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1595_A _7529_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4515__A _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A1 _7450_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__B2 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6718__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5049__C _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__1111_ clkbuf_0__1111_/X VGND VGND VPWR VPWR _6789_/A2 sky130_fd_sc_hd__clkbuf_16
XANTENNA__3952__A3 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4888__C _4888_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5065__B _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3704__A3 _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5780__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3143_A _7041_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_69_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input41_A mgmt_gpio_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6654__A2 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5081__A _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5862__A0 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2890 hold2890/A VGND VGND VPWR VPWR _5626_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4968__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3640__A2 _5803_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6590__A1 _7348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_734 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4450_ _4450_/A0 _5876_/A1 _4454_/S VGND VGND VPWR VPWR _4450_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold207 hold207/A VGND VGND VPWR VPWR _7529_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold218 hold218/A VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold229 hold229/A VGND VGND VPWR VPWR _7532_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3401_ _6890_/Q VGND VGND VPWR VPWR _3401_/Y sky130_fd_sc_hd__inv_2
X_4381_ _4381_/A0 _5817_/A1 _4381_/S VGND VGND VPWR VPWR _4381_/X sky130_fd_sc_hd__mux2_1
X_6120_ _6121_/A _6120_/B _6121_/C VGND VGND VPWR VPWR _6120_/X sky130_fd_sc_hd__and3_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 fanout720/X VGND VGND VPWR VPWR fanout709/X sky130_fd_sc_hd__buf_6
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6441_/D _6433_/D _6067_/B _6434_/B VGND VGND VPWR VPWR _6051_/Y sky130_fd_sc_hd__nand4_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4656__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5853__A0 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5024_/A1 _4669_/X _4974_/B _5038_/C _5158_/A VGND VGND VPWR VPWR _5025_/D
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__4408__A1 _5975_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4959__A2 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6953_ _7575_/CLK _6953_/D fanout735/X VGND VGND VPWR VPWR _6953_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5904_ hold198/X _5904_/A1 hold42/X VGND VGND VPWR VPWR _5904_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold2877_A _7226_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ _4169_/B2 _6884_/D _6834_/X VGND VGND VPWR VPWR _6884_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3631__A2 _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _5835_/A0 _5997_/A1 _5838_/S VGND VGND VPWR VPWR _5835_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5865__S _5865_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5766_ hold20/X _5766_/A1 hold27/X VGND VGND VPWR VPWR _5766_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6581__B2 _7492_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7505_ _7561_/CLK _7505_/D fanout738/X VGND VGND VPWR VPWR _7505_/Q sky130_fd_sc_hd__dfrtp_4
X_4717_ _5387_/C _4717_/B VGND VGND VPWR VPWR _4717_/Y sky130_fd_sc_hd__nand2_4
X_5697_ _5697_/A0 _5994_/A1 _5703_/S VGND VGND VPWR VPWR _5697_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7436_ _7548_/CLK _7436_/D fanout732/X VGND VGND VPWR VPWR _7436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ _4648_/A _4825_/A VGND VGND VPWR VPWR _4726_/B sky130_fd_sc_hd__nand2_4
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4344__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold730 hold730/A VGND VGND VPWR VPWR _7015_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold741 hold741/A VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7367_ _7580_/CLK _7367_/D fanout735/X VGND VGND VPWR VPWR _7367_/Q sky130_fd_sc_hd__dfstp_4
X_4579_ _4831_/A _4767_/A _4909_/D _4772_/B VGND VGND VPWR VPWR _4643_/C sky130_fd_sc_hd__and4_4
XFILLER_162_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold752 _4514_/X VGND VGND VPWR VPWR _7166_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold763 hold763/A VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap471 _4870_/A VGND VGND VPWR VPWR _4947_/C sky130_fd_sc_hd__buf_4
Xhold774 _4193_/X VGND VGND VPWR VPWR _6912_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6318_ _7067_/Q _6317_/B _6332_/C _6092_/X _7178_/Q VGND VGND VPWR VPWR _6318_/X
+ sky130_fd_sc_hd__a32o_1
Xhold785 hold785/A VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_70_csclk_A clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold796 hold796/A VGND VGND VPWR VPWR _7332_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7298_ _7334_/CLK _7298_/D fanout711/X VGND VGND VPWR VPWR _7298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6636__A2 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5439__A3 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6249_ _7421_/Q _6072_/X _6099_/X _7357_/Q _6248_/X VGND VGND VPWR VPWR _6257_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2120 _4228_/X VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3414__A _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2131 _7067_/Q VGND VGND VPWR VPWR hold326/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2142 _5946_/X VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2153 _5964_/X VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2164 _5865_/X VGND VGND VPWR VPWR hold63/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2175 _7657_/A VGND VGND VPWR VPWR hold533/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1430 hold117/X VGND VGND VPWR VPWR _7234_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1441 _4447_/X VGND VGND VPWR VPWR hold1441/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2186 _6917_/Q VGND VGND VPWR VPWR hold565/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2197 hold637/X VGND VGND VPWR VPWR _5734_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1452 hold143/X VGND VGND VPWR VPWR _6916_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1463 _6924_/Q VGND VGND VPWR VPWR hold1463/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1474 hold1474/A VGND VGND VPWR VPWR _5891_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 hold70/X VGND VGND VPWR VPWR _4421_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_61_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7329_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1496 _5928_/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3622__A2 _3617_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5775__S _5775_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input89_A spimemio_flash_io2_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3689__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_14_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7180_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6088__B1 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6627__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4638__A1 _4667_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_29_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7563_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3950_ _7359_/Q _4364_/A _5965_/B _3946_/X _3949_/X VGND VGND VPWR VPWR _3961_/C
+ sky130_fd_sc_hd__a311o_1
XANTENNA__6073__C _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3613__A2 _3508_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3881_ _6875_/Q _4551_/B _4352_/B _3880_/X VGND VGND VPWR VPWR _3881_/X sky130_fd_sc_hd__a31o_1
X_5620_ _5620_/A0 _5732_/A1 _5620_/S VGND VGND VPWR VPWR _5620_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6563__B2 _7339_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_829 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5551_ _4975_/X _5424_/X _5340_/A _5169_/X _5438_/D VGND VGND VPWR VPWR _5551_/X
+ sky130_fd_sc_hd__o2111a_1
X_4502_ _5853_/A0 _4502_/A1 _4502_/S VGND VGND VPWR VPWR _4502_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5482_ _5482_/A _5482_/B _5560_/A VGND VGND VPWR VPWR _5482_/Y sky130_fd_sc_hd__nand3_1
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4326__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7221_ _7075_/CLK _7221_/D _6873_/X VGND VGND VPWR VPWR _7221_/Q sky130_fd_sc_hd__dfrtn_1
XFILLER_144_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4433_ _4433_/A0 _5922_/A0 _4439_/S VGND VGND VPWR VPWR _4433_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7152_ _7201_/CLK _7152_/D fanout726/X VGND VGND VPWR VPWR _7152_/Q sky130_fd_sc_hd__dfrtp_4
X_4364_ _4364_/A _4364_/B _5619_/C VGND VGND VPWR VPWR _4369_/S sky130_fd_sc_hd__and3_2
Xfanout506 _6021_/X VGND VGND VPWR VPWR _6112_/B sky130_fd_sc_hd__buf_12
X_6103_ _7335_/Q _6121_/A _6120_/B _6332_/C _7359_/Q VGND VGND VPWR VPWR _6103_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6618__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout517 _5138_/D VGND VGND VPWR VPWR _5029_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7083_ _7514_/CLK _7083_/D fanout743/X VGND VGND VPWR VPWR _7663_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4295_ _4302_/S _3856_/B _4294_/Y VGND VGND VPWR VPWR _6982_/D sky130_fd_sc_hd__o21ai_1
Xfanout539 hold1494/X VGND VGND VPWR VPWR _6000_/A1 sky130_fd_sc_hd__buf_8
XFILLER_98_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4629__A1 _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6034_ _6099_/D _6019_/Y _6033_/X VGND VGND VPWR VPWR _7591_/D sky130_fd_sc_hd__a21o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4644__A4 _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3852__A2 _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5054__A1 _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5054__B2 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ _7551_/CLK _6936_/D fanout734/X VGND VGND VPWR VPWR _7654_/A sky130_fd_sc_hd__dfrtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout443_A _3860_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3604__A2 hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6867_ _6869_/A _6872_/B VGND VGND VPWR VPWR _6867_/X sky130_fd_sc_hd__and2_1
XFILLER_168_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5818_ _5818_/A0 _5881_/A1 _5820_/S VGND VGND VPWR VPWR _5818_/X sky130_fd_sc_hd__mux2_1
X_6798_ _6797_/X _6798_/B _6798_/C VGND VGND VPWR VPWR _6822_/S sky130_fd_sc_hd__nand3b_4
X_5749_ _5803_/A _5749_/B _5947_/C VGND VGND VPWR VPWR _5757_/S sky130_fd_sc_hd__and3_4
XANTENNA__3907__A3 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7419_ _7471_/CLK _7419_/D fanout730/X VGND VGND VPWR VPWR _7419_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4868__A1 _4571_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold560 hold560/A VGND VGND VPWR VPWR _7294_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold571 hold571/A VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 hold582/A VGND VGND VPWR VPWR _7259_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6609__A2 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input143_A wb_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6490__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6455__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1260 hold2925/X VGND VGND VPWR VPWR _6964_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1271 hold2950/X VGND VGND VPWR VPWR hold2951/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3843__A2 _3535_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1282 hold3223/X VGND VGND VPWR VPWR _7021_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1293 hold3245/X VGND VGND VPWR VPWR hold3246/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6242__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4703__A _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4556__A0 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4795__D _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4080_ _6908_/Q _6882_/Q _4062_/A _4001_/Y VGND VGND VPWR VPWR _4080_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6076__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5284__A1 _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6481__B1 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3834__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold2206_A _7242_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5036__A1 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6233__B1 _6121_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3501__B _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4982_ _4996_/A _5339_/D _5183_/A _5203_/C VGND VGND VPWR VPWR _5044_/C sky130_fd_sc_hd__nand4_2
X_6721_ _7058_/Q _6466_/D _6651_/C _6452_/X _7023_/Q VGND VGND VPWR VPWR _6721_/X
+ sky130_fd_sc_hd__a32o_1
X_3933_ _3933_/A _5619_/A VGND VGND VPWR VPWR _3933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6652_ _7137_/Q _6419_/C _6446_/X _7187_/Q VGND VGND VPWR VPWR _6652_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3864_ _5612_/A _5640_/A _5619_/A VGND VGND VPWR VPWR _3864_/X sky130_fd_sc_hd__and3_1
XANTENNA__6536__A1 _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6536__B2 _7522_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4547__A0 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5603_ _5619_/A _5632_/B _5640_/D VGND VGND VPWR VPWR _5611_/S sky130_fd_sc_hd__and3_4
X_6583_ _7436_/Q _6747_/B _6747_/C _6408_/A _7556_/Q VGND VGND VPWR VPWR _6583_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3795_ _3856_/A _3795_/B VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5534_ _5158_/B _5410_/C _5410_/A _5160_/D _5317_/C VGND VGND VPWR VPWR _5535_/C
+ sky130_fd_sc_hd__a311oi_2
XFILLER_117_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _4601_/Y _4700_/Y _5509_/A3 _5077_/Y VGND VGND VPWR VPWR _5467_/B sky130_fd_sc_hd__a31o_1
X_7204_ _7633_/CLK _7204_/D _6780_/B VGND VGND VPWR VPWR _7204_/Q sky130_fd_sc_hd__dfrtp_1
X_4416_ _4445_/A0 _5853_/A0 _4422_/S VGND VGND VPWR VPWR _4416_/X sky130_fd_sc_hd__mux2_1
X_5396_ _4817_/X _5453_/C _5394_/Y _5395_/X VGND VGND VPWR VPWR _5396_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3522__A1 _7446_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7135_ _7184_/CLK _7135_/D fanout724/X VGND VGND VPWR VPWR _7135_/Q sky130_fd_sc_hd__dfrtp_4
X_4347_ _4347_/A0 _5948_/A1 _4351_/S VGND VGND VPWR VPWR _4347_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout393_A _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout358 _3553_/X VGND VGND VPWR VPWR _4231_/S sky130_fd_sc_hd__buf_12
X_7066_ _7160_/CLK _7066_/D _6872_/A VGND VGND VPWR VPWR _7066_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout369 hold31/X VGND VGND VPWR VPWR _5866_/B sky130_fd_sc_hd__buf_8
X_4278_ _4289_/S _4278_/B VGND VGND VPWR VPWR _4278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6472__B1 _7279_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6017_ _7585_/Q _7586_/Q _7587_/Q _6017_/D VGND VGND VPWR VPWR _6018_/C sky130_fd_sc_hd__nand4_1
XANTENNA_fanout560_A _5726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3825__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clkbuf_0_wbbd_sck/X VGND VGND VPWR VPWR _3443__2/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__6775__A1 _6961_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5578__A2 _4722_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6919_ _7255_/CLK _6919_/D fanout688/X VGND VGND VPWR VPWR _6919_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__4250__A2 hold365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__A _5619_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6527__A1 _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6527__B2 _7458_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4538__A0 _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold390 _5790_/X VGND VGND VPWR VPWR _7395_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3513__B2 _7310_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3816__A2 _5947_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1090 hold3014/X VGND VGND VPWR VPWR hold1090/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6518__A1 _7393_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5248__B _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3580_ _7501_/Q hold41/A _3542_/X _6925_/Q _3579_/X VGND VGND VPWR VPWR _3587_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_127_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3752__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3752__B2 _7482_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6297__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5250_ _4910_/D _5399_/A _4953_/X _5249_/Y VGND VGND VPWR VPWR _5252_/C sky130_fd_sc_hd__a31o_1
XANTENNA__6151__C1 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4201_ _4201_/A0 _4201_/A1 _4429_/B VGND VGND VPWR VPWR _4201_/X sky130_fd_sc_hd__mux2_2
XFILLER_69_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5181_ _5203_/C _5183_/C _5180_/A _5216_/A VGND VGND VPWR VPWR _5181_/X sky130_fd_sc_hd__o211a_1
Xhold2708 _7156_/Q VGND VGND VPWR VPWR hold809/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2719 _7196_/Q VGND VGND VPWR VPWR hold755/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2323_A _7331_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4132_ _4132_/A VGND VGND VPWR VPWR _4132_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4063_ _3401_/Y _6892_/Q _7071_/Q VGND VGND VPWR VPWR _4063_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3512__A _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A2 _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6206__B1 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6221__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4965_ _4966_/A _5203_/A _5029_/A _4847_/X VGND VGND VPWR VPWR _4965_/X sky130_fd_sc_hd__a31o_2
X_6704_ _7114_/Q _6462_/C _6426_/X _6703_/X VGND VGND VPWR VPWR _6704_/X sky130_fd_sc_hd__a31o_1
X_3916_ _7368_/Q _5758_/A _5776_/A _7384_/Q _3860_/X VGND VGND VPWR VPWR _3916_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_189_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6509__B2 _7569_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4896_ _4966_/A _4997_/A _5222_/B _5222_/C VGND VGND VPWR VPWR _4896_/Y sky130_fd_sc_hd__nand4_2
XFILLER_177_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6635_ _7342_/Q _6425_/X _6460_/X _7390_/Q VGND VGND VPWR VPWR _6635_/X sky130_fd_sc_hd__a22o_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ _7246_/Q _5947_/A _5614_/B _3598_/X VGND VGND VPWR VPWR _3847_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3991__B2 _7112_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6566_ _7555_/Q _6408_/A _6408_/D _7539_/Q _6565_/X VGND VGND VPWR VPWR _6569_/C
+ sky130_fd_sc_hd__a221o_1
X_3778_ _7059_/Q _4539_/C _4364_/B _3739_/X VGND VGND VPWR VPWR _3782_/C sky130_fd_sc_hd__a31o_1
XANTENNA__4997__B _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3743__A1 _7562_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5517_ _5561_/A1 _4796_/Y _5471_/X _5516_/X VGND VGND VPWR VPWR _5518_/B sky130_fd_sc_hd__o31a_1
XANTENNA__3743__B2 input38/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6497_ _6649_/S _7615_/Q _6495_/Y _6496_/X VGND VGND VPWR VPWR _6497_/X sky130_fd_sc_hd__a22o_1
XFILLER_133_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5448_ _5445_/X _5448_/B _5508_/A _5448_/D VGND VGND VPWR VPWR _5452_/B sky130_fd_sc_hd__and4b_1
XFILLER_154_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6693__B1 _6466_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5379_ _5480_/A1 _5509_/A3 _4737_/Y _5563_/A1 VGND VGND VPWR VPWR _5379_/X sky130_fd_sc_hd__a211o_1
XANTENNA_fanout775_A _4887_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7118_ _7561_/CLK _7118_/D fanout741/X VGND VGND VPWR VPWR _7118_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6445__B1 _6420_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7049_ _7471_/CLK _7049_/D fanout729/X VGND VGND VPWR VPWR _7049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3422__A _7466_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6748__A1 _7024_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A wb_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6452__B _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3982__A1 _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3982__B2 _7487_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5783__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input71_A mgmt_gpio_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4700__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6684__B1 _6460_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5812__A _5866_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5239__A1 _5222_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4998__B1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _5260_/A _5260_/B _5094_/A VGND VGND VPWR VPWR _4898_/C sky130_fd_sc_hd__and3_2
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3701_ _7475_/Q _3494_/X _3529_/X _7531_/Q _3700_/X VGND VGND VPWR VPWR _3701_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4681_ _5158_/A _4952_/B VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6420_ _6420_/A _6420_/B _6420_/C _6419_/Y VGND VGND VPWR VPWR _6431_/C sky130_fd_sc_hd__nor4b_4
X_3632_ _3632_/A _3632_/B _3632_/C _3632_/D VGND VGND VPWR VPWR _3643_/B sky130_fd_sc_hd__nor4_2
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3725__A1 _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6351_ _7164_/Q _6075_/X _6350_/X _6332_/X _6349_/X VGND VGND VPWR VPWR _6351_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_162_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4610__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3563_ _7302_/Q _5965_/B _3563_/C VGND VGND VPWR VPWR _3563_/X sky130_fd_sc_hd__and3_1
XFILLER_127_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2440_A _7259_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5302_ _4741_/Y _4755_/Y _4687_/Y _5135_/Y _5297_/Y VGND VGND VPWR VPWR _5303_/D
+ sky130_fd_sc_hd__o221a_1
X_6282_ _7286_/Q _6036_/Y _6623_/B1 VGND VGND VPWR VPWR _6282_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3494_ _5590_/A hold32/A _5722_/B VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__and3_4
Xhold3206 hold3206/A VGND VGND VPWR VPWR _4329_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3217 hold3217/A VGND VGND VPWR VPWR _4383_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5233_ _4954_/C _4933_/A _4943_/B _5102_/B _4790_/C VGND VGND VPWR VPWR _5233_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3228 _4213_/X VGND VGND VPWR VPWR hold3228/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3239 _4304_/X VGND VGND VPWR VPWR hold3239/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5722__A hold40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2505 hold917/X VGND VGND VPWR VPWR _4354_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2516 hold485/X VGND VGND VPWR VPWR _4181_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4150__A1 _4150_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2527 hold909/X VGND VGND VPWR VPWR _5729_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2538 hold833/X VGND VGND VPWR VPWR _4554_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5164_ _5164_/A _5164_/B VGND VGND VPWR VPWR _5167_/A sky130_fd_sc_hd__nor2_1
Xhold1804 _5618_/X VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2549 _5798_/X VGND VGND VPWR VPWR hold912/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1815 hold30/X VGND VGND VPWR VPWR _3557_/C sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1826 hold435/X VGND VGND VPWR VPWR _5886_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4115_ _4424_/B _4115_/B VGND VGND VPWR VPWR _7101_/D sky130_fd_sc_hd__nand2b_1
Xhold1837 _7286_/Q VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5095_ _4748_/A _4596_/X _5096_/A _5093_/Y VGND VGND VPWR VPWR _5097_/A sky130_fd_sc_hd__a31oi_2
Xhold1848 _7272_/Q VGND VGND VPWR VPWR hold413/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1859 _7134_/Q VGND VGND VPWR VPWR hold363/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4046_ _6910_/Q _6909_/Q _6908_/Q _4058_/A VGND VGND VPWR VPWR _4047_/S sky130_fd_sc_hd__and4_1
XANTENNA__6442__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5650__A1 _5650_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ _5997_/A0 _5997_/A1 _6000_/S VGND VGND VPWR VPWR _5997_/X sky130_fd_sc_hd__mux2_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4948_ _4966_/A _4948_/B _4948_/C _5248_/C VGND VGND VPWR VPWR _4949_/B sky130_fd_sc_hd__and4_1
X_7667_ _7667_/A VGND VGND VPWR VPWR _7667_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4879_ _4840_/D _4887_/B _4945_/A _4879_/D VGND VGND VPWR VPWR _4918_/D sky130_fd_sc_hd__and4bb_4
XFILLER_165_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6618_ _7549_/Q _6419_/A _6455_/X _7461_/Q _6602_/X VGND VGND VPWR VPWR _6618_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7598_ _7610_/CLK _7598_/D fanout694/X VGND VGND VPWR VPWR _7598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6549_ _7571_/Q _6424_/X _6427_/X _7579_/Q VGND VGND VPWR VPWR _6549_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3417__A _7506_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput270 _6913_/Q VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XANTENNA__6130__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput281 _7239_/Q VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
Xoutput292 _6926_/Q VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
XANTENNA__4141__A1 _7578_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3495__A3 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5641__A1 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5778__S _5784_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6463__A _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5079__A _5100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3955__A1 _7527_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5157__B1 _4977_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire353 _6118_/Y VGND VGND VPWR VPWR _6122_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_139_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire375 _5127_/A VGND VGND VPWR VPWR wire375/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output275_A _6918_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4380__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_152_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6657__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5880__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5920_ _5920_/A _5992_/D VGND VGND VPWR VPWR _5928_/S sky130_fd_sc_hd__nand2_8
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5851_ _5914_/A1 _5851_/A1 _5856_/S VGND VGND VPWR VPWR _5851_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6188__A2 _6097_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4802_ _4802_/A _5404_/C VGND VGND VPWR VPWR _4802_/Y sky130_fd_sc_hd__nand2_1
X_5782_ _5953_/A1 _5782_/A1 _5784_/S VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7521_ _7531_/CLK _7521_/D fanout743/X VGND VGND VPWR VPWR _7521_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3946__A1 _7295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4733_ _4733_/A _4733_/B _4772_/A VGND VGND VPWR VPWR _5404_/C sky130_fd_sc_hd__and3_4
XFILLER_159_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7452_ _7572_/CLK _7452_/D fanout733/X VGND VGND VPWR VPWR _7452_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_175_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4664_ _4568_/Y _4984_/C _4861_/B VGND VGND VPWR VPWR _4974_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5699__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6403_ _6463_/A _6427_/A _6468_/C VGND VGND VPWR VPWR _6408_/A sky130_fd_sc_hd__and3_4
XFILLER_119_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3615_ _7292_/Q _5668_/A _3549_/X input49/X _3614_/X VGND VGND VPWR VPWR _3623_/C
+ sky130_fd_sc_hd__a221o_1
X_7383_ _7580_/CLK _7383_/D fanout733/X VGND VGND VPWR VPWR _7383_/Q sky130_fd_sc_hd__dfstp_4
Xhold901 hold901/A VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6360__A2 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4595_ _5295_/A _5295_/D VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__nand2_8
Xhold912 hold912/A VGND VGND VPWR VPWR _7402_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold923 hold923/A VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6334_ _7144_/Q _6121_/C _6116_/C _6121_/B VGND VGND VPWR VPWR _6334_/X sky130_fd_sc_hd__o211a_1
Xhold934 _4494_/X VGND VGND VPWR VPWR _7149_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3546_ _7422_/Q hold32/A hold90/A _3545_/X _7350_/Q VGND VGND VPWR VPWR _3546_/X
+ sky130_fd_sc_hd__a32o_1
Xhold945 hold945/A VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap653 _5549_/A3 VGND VGND VPWR VPWR _5055_/C sky130_fd_sc_hd__buf_2
Xhold956 _5827_/X VGND VGND VPWR VPWR _7428_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold967 hold967/A VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold978 hold978/A VGND VGND VPWR VPWR _7120_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3003 _7257_/Q VGND VGND VPWR VPWR _4078_/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold989 hold989/A VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6265_ _7390_/Q _6274_/A3 _6079_/X _7334_/Q _6264_/X VGND VGND VPWR VPWR _6265_/X
+ sky130_fd_sc_hd__a221o_1
Xhold3014 hold3014/A VGND VGND VPWR VPWR hold3014/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3025 hold3025/A VGND VGND VPWR VPWR hold3025/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_3477_ _3557_/C _3477_/B VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__nor2_4
XFILLER_89_749 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4994__C _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3036 hold3036/A VGND VGND VPWR VPWR hold3036/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3047 hold3047/A VGND VGND VPWR VPWR hold3047/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2302 _7579_/Q VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5216_ _5216_/A _5342_/B _5216_/C VGND VGND VPWR VPWR _5216_/X sky130_fd_sc_hd__and3_2
Xhold3058 _7630_/Q VGND VGND VPWR VPWR _6783_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2313 hold675/X VGND VGND VPWR VPWR _5780_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2324 hold589/X VGND VGND VPWR VPWR _5718_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3069 _7056_/Q VGND VGND VPWR VPWR hold3069/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6196_ _7443_/Q _6097_/X _6121_/X _7307_/Q _6195_/X VGND VGND VPWR VPWR _6196_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6663__A3 _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2335 _7308_/Q VGND VGND VPWR VPWR hold803/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1601 _7517_/Q VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2346 _5799_/X VGND VGND VPWR VPWR hold568/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5871__A1 _5979_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2357 hold741/X VGND VGND VPWR VPWR _5617_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1612 hold226/X VGND VGND VPWR VPWR _5854_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1623 _5715_/X VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ _4778_/A _4758_/X _5410_/B _5086_/B _5152_/B2 VGND VGND VPWR VPWR _5148_/C
+ sky130_fd_sc_hd__a32o_1
Xhold2368 hold685/X VGND VGND VPWR VPWR _5834_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2379 _7277_/Q VGND VGND VPWR VPWR hold821/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1634 _5770_/X VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_151_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1645 _5637_/X VGND VGND VPWR VPWR hold264/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1656 hold401/X VGND VGND VPWR VPWR _5724_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1667 _5706_/X VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5078_ _4571_/Y _4843_/A _4727_/Y _5516_/A3 _5077_/Y VGND VGND VPWR VPWR _5467_/A
+ sky130_fd_sc_hd__o32a_1
Xhold1678 _6951_/Q VGND VGND VPWR VPWR hold188/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1689 _7470_/Q VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4029_ _6902_/Q _6901_/Q _6900_/Q _4025_/A VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__a31o_1
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4515__B _4515_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3937__A1 _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1755_A _7512_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6351__A2 _6075_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5154__A3 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4362__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6639__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6103__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3456__A_N _4181_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input34_A mask_rev_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2880 hold2880/A VGND VGND VPWR VPWR _5942_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2891 _7498_/Q VGND VGND VPWR VPWR hold2891/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3625__B1 hold77/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5090__A2 _4960_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3640__A3 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4050__A0 _6897_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6590__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__A3 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5971__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold219 hold219/A VGND VGND VPWR VPWR _7145_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_3400_ _3400_/A VGND VGND VPWR VPWR _3400_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4353__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2069_A _7408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4380_ _4380_/A0 _5585_/A0 _4381_/S VGND VGND VPWR VPWR _4380_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__B1 _4687_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6050_ _7594_/Q _6429_/C _6441_/D _6433_/D VGND VGND VPWR VPWR _6050_/Y sky130_fd_sc_hd__nand4_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6087__B _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5001_ _5024_/A1 _4669_/X _4974_/B _5404_/D _5038_/C VGND VGND VPWR VPWR _5025_/C
+ sky130_fd_sc_hd__o2111ai_4
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5605__A1 _5645_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6307__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6952_ _7551_/CLK _6952_/D fanout734/X VGND VGND VPWR VPWR _6952_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3520__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4959__A3 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5903_ _5948_/A1 _5903_/A1 hold42/X VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__mux2_1
X_6883_ _4169_/B2 _6883_/D _6833_/X VGND VGND VPWR VPWR _6883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5834_ _5834_/A0 _5969_/A1 _5838_/S VGND VGND VPWR VPWR _5834_/X sky130_fd_sc_hd__mux2_1
X_5765_ _5999_/A1 _5765_/A1 hold27/X VGND VGND VPWR VPWR _5765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6581__A2 _6425_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4989__C _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7504_ _7531_/CLK _7504_/D fanout743/X VGND VGND VPWR VPWR _7504_/Q sky130_fd_sc_hd__dfstp_4
X_4716_ _5260_/A _5079_/B VGND VGND VPWR VPWR _4716_/Y sky130_fd_sc_hd__nand2_4
X_5696_ _5696_/A0 hold487/X _5703_/S VGND VGND VPWR VPWR _5696_/X sky130_fd_sc_hd__mux2_1
X_7435_ _7435_/CLK _7435_/D fanout730/X VGND VGND VPWR VPWR _7435_/Q sky130_fd_sc_hd__dfrtp_4
X_4647_ _4646_/A _4646_/B _4643_/Y _4674_/A VGND VGND VPWR VPWR _4726_/A sky130_fd_sc_hd__a2bb2oi_4
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6333__A2 _6112_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5881__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7366_ _7478_/CLK _7366_/D fanout713/X VGND VGND VPWR VPWR _7366_/Q sky130_fd_sc_hd__dfrtp_4
Xhold720 hold720/A VGND VGND VPWR VPWR _7171_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4578_ _4984_/C _4578_/B VGND VGND VPWR VPWR _4675_/C sky130_fd_sc_hd__nor2_8
Xhold731 hold731/A VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold742 _5617_/X VGND VGND VPWR VPWR _7246_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold753 hold753/A VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_13_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6317_ _7047_/Q _6317_/B _6317_/C VGND VGND VPWR VPWR _6317_/X sky130_fd_sc_hd__and3_1
Xhold764 _4525_/X VGND VGND VPWR VPWR _7175_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout590_A hold487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3529_ _5938_/A _5938_/B _5938_/C VGND VGND VPWR VPWR _3529_/X sky130_fd_sc_hd__and3_4
X_7297_ _7329_/CLK _7297_/D fanout704/X VGND VGND VPWR VPWR _7297_/Q sky130_fd_sc_hd__dfrtp_4
Xhold775 hold775/A VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold786 _4205_/X VGND VGND VPWR VPWR _6920_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold797 hold797/A VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6248_ _7429_/Q _6112_/C _6074_/X _6120_/X _7341_/Q VGND VGND VPWR VPWR _6248_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2110 hold489/X VGND VGND VPWR VPWR _4230_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2121 _7658_/A VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5844__A1 _5853_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2132 hold326/X VGND VGND VPWR VPWR _4402_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6428__D _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2143 _7210_/Q VGND VGND VPWR VPWR hold393/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2154 _7342_/Q VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6179_ _7450_/Q _6144_/A _6116_/A _6274_/A3 _7514_/Q VGND VGND VPWR VPWR _6179_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2165 _7650_/A VGND VGND VPWR VPWR hold527/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1420 _4189_/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2176 hold533/X VGND VGND VPWR VPWR _4411_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1431 _6885_/Q VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1442 hold1442/A VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2187 hold565/X VGND VGND VPWR VPWR _4200_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1453 _7661_/A VGND VGND VPWR VPWR hold81/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2198 _5734_/X VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_57_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1464 hold1464/A VGND VGND VPWR VPWR _4209_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1475 _5891_/X VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1486 _4421_/X VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3870__A3 _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1497 hold53/X VGND VGND VPWR VPWR _7518_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3430__A _7402_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4280__A0 _3922_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__A_N _6429_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5375__A3 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5780__A0 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6324__A2 _6082_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5791__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4335__A1 _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6088__B2 _7463_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6627__A3 _6428_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5835__A1 _5997_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4638__A2 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__buf_4
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5966__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3880_ _7376_/Q _3498_/X _3658_/X _7113_/Q VGND VGND VPWR VPWR _3880_/X sky130_fd_sc_hd__a22o_1
XFILLER_188_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6563__A2 _6574_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2186_A _6917_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5550_ _5550_/A _5550_/B _5550_/C _5550_/D VGND VGND VPWR VPWR _5550_/Y sky130_fd_sc_hd__nand4_2
X_4501_ _5585_/A0 _4501_/A1 _4502_/S VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5481_ _5481_/A _5481_/B _5481_/C VGND VGND VPWR VPWR _5560_/A sky130_fd_sc_hd__and3_1
XANTENNA__4747__A_N _4879_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7220_ _4150_/A1 _7220_/D _6872_/X VGND VGND VPWR VPWR _7220_/Q sky130_fd_sc_hd__dfrtn_1
X_4432_ _4432_/A0 _5975_/A0 _4439_/S VGND VGND VPWR VPWR _4432_/X sky130_fd_sc_hd__mux2_1
XANTENNA_hold42_A hold42/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7151_ _7395_/CLK _7151_/D fanout737/X VGND VGND VPWR VPWR _7151_/Q sky130_fd_sc_hd__dfrtp_4
X_4363_ _4363_/A0 _5817_/A1 _4363_/S VGND VGND VPWR VPWR _4363_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3515__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6102_ _6102_/A _6102_/B _6102_/C _6102_/D VGND VGND VPWR VPWR _6122_/A sky130_fd_sc_hd__nor4_4
Xfanout507 _5216_/C VGND VGND VPWR VPWR _5339_/C sky130_fd_sc_hd__buf_6
Xfanout518 _4983_/C VGND VGND VPWR VPWR _5399_/C sky130_fd_sc_hd__buf_6
X_7082_ _7519_/CLK _7082_/D fanout742/X VGND VGND VPWR VPWR _7662_/A sky130_fd_sc_hd__dfrtp_1
Xfanout529 _4625_/Y VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__buf_6
X_4294_ _4302_/S _4294_/B VGND VGND VPWR VPWR _4294_/Y sky130_fd_sc_hd__nand2_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5826__A1 _5826_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6033_ _6099_/D _6028_/Y _6081_/C _6032_/B _6019_/A VGND VGND VPWR VPWR _6033_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_113_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4991__D _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7332__RESET_B fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__B2 _7485_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_3__f_mgmt_gpio_in[4]_A clkbuf_0_mgmt_gpio_in[4]/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ _7548_/CLK _6935_/D fanout731/X VGND VGND VPWR VPWR _6935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5876__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3604__A3 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6866_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6866_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout436_A _4491_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_849 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5817_ _5817_/A0 _5817_/A1 _5820_/S VGND VGND VPWR VPWR _5817_/X sky130_fd_sc_hd__mux2_1
X_6797_ _4427_/D _6794_/Y _6795_/Y _4427_/B _4430_/C VGND VGND VPWR VPWR _6797_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6554__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5762__A0 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5748_ _5748_/A0 hold20/X _5748_/S VGND VGND VPWR VPWR _5748_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5679_ hold375/X _5949_/A1 _5685_/S VGND VGND VPWR VPWR _5679_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7418_ _7548_/CLK _7418_/D fanout732/X VGND VGND VPWR VPWR _7418_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_163_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7349_ _7541_/CLK _7349_/D fanout713/X VGND VGND VPWR VPWR _7349_/Q sky130_fd_sc_hd__dfrtp_4
Xhold550 _5970_/X VGND VGND VPWR VPWR _7555_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold561 hold561/A VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold572 _5601_/X VGND VGND VPWR VPWR _7233_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_150_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3425__A _7442_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold583 hold583/A VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold1718_A _7360_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold594 hold594/A VGND VGND VPWR VPWR _7239_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3540__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold383_A _7464_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5817__A1 _5817_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5640__A _5640_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6490__A1 _7496_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6490__B2 _7560_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input136_A wb_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1250 _7208_/Q VGND VGND VPWR VPWR _3453_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1261 hold2907/X VGND VGND VPWR VPWR hold2908/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1272 hold2952/X VGND VGND VPWR VPWR _7179_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1283 hold3242/X VGND VGND VPWR VPWR hold3243/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1294 _4204_/X VGND VGND VPWR VPWR _6919_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5786__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4703__B _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6890__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_185_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4308__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5808__A1 _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5284__A2 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput170 wb_we_i VGND VGND VPWR VPWR _6824_/C sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3834__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _5339_/D _5029_/A _5034_/C VGND VGND VPWR VPWR _5047_/A sky130_fd_sc_hd__and3_2
XANTENNA__5696__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3932_ _7157_/Q _4539_/C _5632_/B _3617_/X _7229_/Q VGND VGND VPWR VPWR _3932_/X
+ sky130_fd_sc_hd__a32o_2
X_6720_ _7199_/Q _6463_/A _6574_/C _6463_/X _7164_/Q VGND VGND VPWR VPWR _6720_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6651_ _7036_/Q _6651_/B _6651_/C VGND VGND VPWR VPWR _6651_/X sky130_fd_sc_hd__and3_1
X_3863_ _3863_/A _5640_/A _4328_/A _5612_/B VGND VGND VPWR VPWR _3863_/X sky130_fd_sc_hd__and4_1
XFILLER_20_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6536__A2 _6042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5602_ hold116/X _5627_/A1 _5602_/S VGND VGND VPWR VPWR _5602_/X sky130_fd_sc_hd__mux2_1
X_6582_ _7404_/Q _6409_/X _6420_/B _7308_/Q _6581_/X VGND VGND VPWR VPWR _6582_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_164_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3794_ _3744_/X _3750_/X _3794_/C _3794_/D VGND VGND VPWR VPWR _3795_/B sky130_fd_sc_hd__and4bb_4
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5533_ _5533_/A _5533_/B VGND VGND VPWR VPWR _5533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_csclk clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR _7309_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3770__A2 _4352_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5464_ _5294_/Y _5422_/X _5463_/X VGND VGND VPWR VPWR _5464_/Y sky130_fd_sc_hd__o21ai_1
X_7203_ _7633_/CLK _7203_/D _6780_/B VGND VGND VPWR VPWR _7203_/Q sky130_fd_sc_hd__dfrtp_1
X_4415_ _4415_/A0 _4414_/X _4423_/S VGND VGND VPWR VPWR _4415_/X sky130_fd_sc_hd__mux2_1
X_5395_ wire674/X _4811_/D _5524_/A3 _5277_/X VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5511__A3 _5081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7134_ _7176_/CLK _7134_/D fanout724/X VGND VGND VPWR VPWR _7134_/Q sky130_fd_sc_hd__dfstp_4
X_4346_ _5640_/B _5596_/A _4346_/C _5640_/D VGND VGND VPWR VPWR _4351_/S sky130_fd_sc_hd__and4_2
XANTENNA__3522__A2 hold31/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7255_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7065_ _7181_/CLK _7065_/D fanout721/X VGND VGND VPWR VPWR _7065_/Q sky130_fd_sc_hd__dfrtp_4
Xfanout359 _3552_/X VGND VGND VPWR VPWR _4248_/S sky130_fd_sc_hd__buf_12
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4277_ _4425_/C _6780_/B VGND VGND VPWR VPWR _4289_/S sky130_fd_sc_hd__nand2_8
XFILLER_140_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout386_A _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6016_ _7585_/Q _7586_/Q _6017_/D _7587_/Q VGND VGND VPWR VPWR _6018_/B sky130_fd_sc_hd__a31o_1
XFILLER_101_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6472__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3825__A3 _4364_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout553_A _5673_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6224__A1 _7468_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6775__A2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout720_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3589__A2 _3501_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6918_ _7238_/CLK _6918_/D fanout690/X VGND VGND VPWR VPWR _6918_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4250__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__B _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3994__C1 _3992_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_803 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7181_/CLK sky130_fd_sc_hd__clkbuf_16
X_6849_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6849_/X sky130_fd_sc_hd__and2_1
XFILLER_23_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6527__A2 _6561_/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold1668_A _7465_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7562_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3761__A2 _5695_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6160__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5502__A3 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold380 hold380/A VGND VGND VPWR VPWR _7288_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold391 hold391/A VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3816__A3 _5619_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1080 hold2998/X VGND VGND VPWR VPWR hold1080/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 hold1091/A VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
XTAP_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6766__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6620__D1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6518__A2 _6420_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4529__A1 _4547_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5248__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3752__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_170_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6151__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ _4200_/A0 _5954_/A1 _4202_/S VGND VGND VPWR VPWR _4200_/X sky130_fd_sc_hd__mux2_1
X_5180_ _5180_/A _5180_/B _5216_/A VGND VGND VPWR VPWR _5180_/X sky130_fd_sc_hd__and3_1
XFILLER_123_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2709 hold809/X VGND VGND VPWR VPWR _4502_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4131_ _6896_/Q _4131_/B VGND VGND VPWR VPWR _4132_/A sky130_fd_sc_hd__nor2_2
X_4062_ _4062_/A _4062_/B VGND VGND VPWR VPWR _4062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3512__B _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__A3 _5623_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6206__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6757__A2 _6058_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4964_ _4963_/X _4960_/B _4855_/Y _4962_/Y VGND VGND VPWR VPWR _4964_/Y sky130_fd_sc_hd__o211ai_4
X_6703_ _6876_/Q _6466_/D _6459_/C _6421_/X _7008_/Q VGND VGND VPWR VPWR _6703_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3915_ input35/X _5695_/A _5612_/B _5704_/A _7320_/Q VGND VGND VPWR VPWR _3915_/X
+ sky130_fd_sc_hd__a32o_4
X_4895_ _4942_/A _5005_/A _5222_/B _4898_/C VGND VGND VPWR VPWR _4895_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__6509__A2 _6419_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5717__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6634_ _7334_/Q _6423_/X _6454_/X _7494_/Q _6633_/X VGND VGND VPWR VPWR _6634_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3991__A2 _5740_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3846_ _4076_/B _3552_/X _3652_/X _7149_/Q _3845_/X VGND VGND VPWR VPWR _3846_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_149_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3777_ _7282_/Q _3558_/X _3682_/X _7227_/Q _3776_/X VGND VGND VPWR VPWR _3782_/B
+ sky130_fd_sc_hd__a221o_4
X_6565_ _7307_/Q _6420_/B _6422_/X _7291_/Q VGND VGND VPWR VPWR _6565_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3743__A2 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5516_ _4705_/Y _4787_/Y _5516_/A3 _4798_/Y _4709_/Y VGND VGND VPWR VPWR _5516_/X
+ sky130_fd_sc_hd__o32a_1
X_6496_ _7280_/Q _6431_/Y _6623_/B1 VGND VGND VPWR VPWR _6496_/X sky130_fd_sc_hd__o21a_1
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _4889_/A _4726_/Y _4889_/B _5528_/A3 _5355_/D VGND VGND VPWR VPWR _5508_/A
+ sky130_fd_sc_hd__o41a_1
XFILLER_145_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5378_ _5480_/A1 _5509_/A3 _4741_/Y _5563_/A1 VGND VGND VPWR VPWR _5378_/X sky130_fd_sc_hd__a211o_1
XFILLER_160_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5902__B _5947_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7117_ _7519_/CLK _7117_/D fanout741/X VGND VGND VPWR VPWR _7117_/Q sky130_fd_sc_hd__dfrtp_4
X_4329_ _4329_/A0 _5582_/A0 _4333_/S VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout768_A _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6445__B2 _7295_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7048_ _7176_/CLK _7048_/D fanout722/X VGND VGND VPWR VPWR _7048_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6748__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5420__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5708__A0 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5068__C _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3982__A2 _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6381__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input64_A mgmt_gpio_in[35] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_821 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6684__A1 _7027_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7435__RESET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5812__B _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__A1 _7319_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6436__B2 _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout690 fanout691/X VGND VGND VPWR VPWR fanout690/X sky130_fd_sc_hd__buf_8
XTAP_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6739__A2 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _7523_/Q _5785_/B _4376_/B _3673_/X _7201_/Q VGND VGND VPWR VPWR _3700_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3973__A2 _5947_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4680_ _5158_/A _5248_/A _5248_/B VGND VGND VPWR VPWR _4830_/A sky130_fd_sc_hd__and3_1
XFILLER_187_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3631_ _4173_/A _4248_/S _3553_/X input40/X _3630_/X VGND VGND VPWR VPWR _3632_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5175__A1 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6372__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2266_A _6923_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6350_ _7199_/Q _6332_/B _6079_/X _6072_/X _7154_/Q VGND VGND VPWR VPWR _6350_/X
+ sky130_fd_sc_hd__a32o_1
X_3562_ _5590_/A _5596_/B _3562_/C VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__and3_2
XANTENNA__3725__A2 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5301_ _5494_/B2 _4730_/Y _4731_/Y _5138_/Y _5300_/X VGND VGND VPWR VPWR _5405_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__6124__B1 _6122_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6281_ _6266_/X _6268_/X _6280_/Y VGND VGND VPWR VPWR _6281_/X sky130_fd_sc_hd__a21bo_2
XFILLER_127_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3493_ _5803_/A _5590_/A _5640_/B VGND VGND VPWR VPWR _3493_/X sky130_fd_sc_hd__and3_2
Xhold3207 _4329_/X VGND VGND VPWR VPWR hold3207/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5232_ _4790_/C _4885_/X _4922_/B VGND VGND VPWR VPWR _5444_/D sky130_fd_sc_hd__a21oi_1
Xhold3218 _4383_/X VGND VGND VPWR VPWR hold3218/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold3229 hold3229/A VGND VGND VPWR VPWR _6927_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_170_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2506 _4354_/X VGND VGND VPWR VPWR hold918/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5722__B _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2517 _4181_/X VGND VGND VPWR VPWR hold486/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5163_ _5163_/A _5163_/B _5163_/C VGND VGND VPWR VPWR _5164_/B sky130_fd_sc_hd__nand3_1
Xhold2528 _5729_/X VGND VGND VPWR VPWR hold910/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2539 _4554_/X VGND VGND VPWR VPWR hold834/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1805 hold289/X VGND VGND VPWR VPWR _7247_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_4114_ _4096_/X _4114_/B VGND VGND VPWR VPWR _4115_/B sky130_fd_sc_hd__nand2b_1
Xhold1816 _5874_/S VGND VGND VPWR VPWR _5871_/S sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1827 _5886_/X VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5094_ _5094_/A _5096_/A VGND VGND VPWR VPWR _5473_/D sky130_fd_sc_hd__nand2_1
Xhold1838 hold108/X VGND VGND VPWR VPWR _5667_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1849 hold413/X VGND VGND VPWR VPWR _5652_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4045_ _6910_/Q _6908_/Q _4058_/A VGND VGND VPWR VPWR _4076_/C sky130_fd_sc_hd__and3_1
XANTENNA__5650__A2 hold365/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A0 _5996_/A1 _6000_/S VGND VGND VPWR VPWR _5996_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ _4948_/B _4948_/C _4947_/C _4954_/A VGND VGND VPWR VPWR _4947_/Y sky130_fd_sc_hd__nand4_4
XFILLER_177_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3964__A2 _3525_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7666_ _7666_/A VGND VGND VPWR VPWR _7666_/X sky130_fd_sc_hd__clkbuf_2
X_4878_ _5065_/A _4954_/C _5183_/C _4907_/B VGND VGND VPWR VPWR _4906_/D sky130_fd_sc_hd__nand4_1
X_6617_ _7565_/Q _6419_/C _6466_/X _7509_/Q _6601_/X VGND VGND VPWR VPWR _6617_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_193_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3829_ _7433_/Q _3525_/X _4485_/A _7144_/Q VGND VGND VPWR VPWR _3829_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6363__B1 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7597_ _7610_/CLK _7597_/D fanout693/X VGND VGND VPWR VPWR _7597_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_193_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6548_ _6547_/X _6572_/A2 _6573_/S VGND VGND VPWR VPWR _6548_/X sky130_fd_sc_hd__mux2_1
XFILLER_134_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6115__B1 _6379_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6479_ _7568_/Q _6424_/X _6474_/X _6478_/X _6430_/X VGND VGND VPWR VPWR _6479_/X
+ sky130_fd_sc_hd__a2111o_1
Xoutput260 _7224_/Q VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput271 _6914_/Q VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
XFILLER_160_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput282 _7240_/Q VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XANTENNA__5632__B _5632_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4141__A2 _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput293 _6911_/Q VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_102_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6447__C _6447_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3433__A _7378_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_785 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3955__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6354__B1 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire354 _6485_/Y VGND VGND VPWR VPWR _6495_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3707__A2 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output268_A _7231_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6657__A1 _7132_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6657__B2 _6988_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_590 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5969__S _5973_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4174__A _4174_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5850_ _5922_/A0 _5850_/A1 _5856_/S VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__mux2_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4801_ _4802_/A _4801_/B _4801_/C VGND VGND VPWR VPWR _4823_/B sky130_fd_sc_hd__and3_2
XANTENNA__6593__B1 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5781_ _5997_/A1 _5781_/A1 _5784_/S VGND VGND VPWR VPWR _5781_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7520_ _7562_/CLK _7520_/D fanout740/X VGND VGND VPWR VPWR _7520_/Q sky130_fd_sc_hd__dfstp_4
X_4732_ _4823_/D _4822_/D _4755_/A _5005_/A VGND VGND VPWR VPWR _4732_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3946__A2 _5965_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7451_ _7519_/CLK _7451_/D fanout741/X VGND VGND VPWR VPWR _7451_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6345__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4663_ _4667_/A _4667_/B _4831_/A VGND VGND VPWR VPWR _4861_/B sky130_fd_sc_hd__o21bai_4
XFILLER_159_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2550_A _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3518__A hold47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6402_ _6466_/A _6466_/B VGND VGND VPWR VPWR _6402_/Y sky130_fd_sc_hd__nor2_8
X_3614_ _7548_/Q _3637_/C hold90/A _5974_/A _7564_/Q VGND VGND VPWR VPWR _3614_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_190_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4594_ _4825_/A _5071_/B _5071_/C _4755_/A VGND VGND VPWR VPWR _4594_/Y sky130_fd_sc_hd__nor4_2
X_7382_ _7579_/CLK hold51/X fanout731/X VGND VGND VPWR VPWR _7382_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 _5737_/X VGND VGND VPWR VPWR _7348_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6360__A3 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold913 hold913/A VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3545_ _5590_/A _5722_/B _3562_/C VGND VGND VPWR VPWR _3545_/X sky130_fd_sc_hd__and3_4
Xhold924 hold924/A VGND VGND VPWR VPWR _7421_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6333_ _7194_/Q _6112_/B _6120_/B _6379_/B1 _7189_/Q VGND VGND VPWR VPWR _6333_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold935 hold935/A VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold946 _5809_/X VGND VGND VPWR VPWR _7412_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap665 fanout661/A VGND VGND VPWR VPWR _4778_/B sky130_fd_sc_hd__clkbuf_4
Xhold957 hold957/A VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold968 _4500_/X VGND VGND VPWR VPWR _7154_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6648__B2 _6431_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6264_ _7294_/Q _6144_/A _6270_/C1 _6074_/X _7302_/Q VGND VGND VPWR VPWR _6264_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_88_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3004 _5650_/A1 VGND VGND VPWR VPWR _5633_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3476_ _3511_/C _3476_/B VGND VGND VPWR VPWR _3477_/B sky130_fd_sc_hd__nand2b_2
Xhold3015 _7567_/Q VGND VGND VPWR VPWR hold3015/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3026 _7551_/Q VGND VGND VPWR VPWR hold3026/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3037 _7575_/Q VGND VGND VPWR VPWR hold3037/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_5215_ _4622_/Y _4709_/Y _4726_/Y _5214_/X VGND VGND VPWR VPWR _5223_/A sky130_fd_sc_hd__o31a_1
Xhold2303 hold539/X VGND VGND VPWR VPWR _5997_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5320__A1 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3048 _7262_/Q VGND VGND VPWR VPWR hold999/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6195_ _7499_/Q _6075_/A _6388_/A3 _6116_/X _7315_/Q VGND VGND VPWR VPWR _6195_/X
+ sky130_fd_sc_hd__a32o_1
Xhold2314 _5780_/X VGND VGND VPWR VPWR hold676/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3059 hold3059/A VGND VGND VPWR VPWR hold3059/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2325 _5718_/X VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2336 hold803/X VGND VGND VPWR VPWR _5692_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1602 hold68/X VGND VGND VPWR VPWR _5927_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2347 _6968_/Q VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5146_ _5404_/C _5410_/B _4977_/X _4776_/A VGND VGND VPWR VPWR _5308_/A sky130_fd_sc_hd__a31o_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1613 _5854_/X VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2358 _6953_/Q VGND VGND VPWR VPWR hold545/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2369 _5834_/X VGND VGND VPWR VPWR hold686/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1624 _7549_/Q VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3882__A1 _7352_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1635 hold215/X VGND VGND VPWR VPWR _7377_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5879__S _5883_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3882__B2 _7042_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1646 hold264/X VGND VGND VPWR VPWR _7260_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5077_ _5260_/C _5077_/B VGND VGND VPWR VPWR _5077_/Y sky130_fd_sc_hd__nand2_4
Xhold1657 _5724_/X VGND VGND VPWR VPWR hold402/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1668 _7465_/Q VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1679 hold188/X VGND VGND VPWR VPWR _4253_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6820__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4028_ _4028_/A0 _4027_/Y _4040_/A VGND VGND VPWR VPWR _6905_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6820__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4515__C _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6179__A3 _6116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5979_ _5979_/A0 _5979_/A1 _5982_/S VGND VGND VPWR VPWR _5979_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3937__A2 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7649_ _7649_/A VGND VGND VPWR VPWR _7649_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6336__B1 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3428__A _7418_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_176_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1915_A _7363_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6639__A1 _7350_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6639__B2 _7414_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input166_A wb_sel_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6103__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4259__A _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2870 hold2870/A VGND VGND VPWR VPWR _5924_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5789__S hold48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input27_A mask_rev_in[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2881 _5942_/X VGND VGND VPWR VPWR hold2881/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2892 hold2892/A VGND VGND VPWR VPWR _5906_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6811__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6811__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3625__B2 _7524_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_141_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4968__A4 _4679_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5378__A1 _5480_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6575__B1 _6462_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4722__A _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5393__A4 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_user_clock user_clock VGND VGND VPWR VPWR clkbuf_0_user_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6342__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5029_/A _5038_/C _5216_/A VGND VGND VPWR VPWR _5026_/B sky130_fd_sc_hd__and3_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5699__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6802__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6802__B2 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6951_ _7551_/CLK _6951_/D fanout734/X VGND VGND VPWR VPWR _6951_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4616__B _4645_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3520__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5902_ hold41/X _5947_/C VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__nand2_8
X_6882_ _7075_/CLK _6882_/D _6832_/X VGND VGND VPWR VPWR _6882_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5369__A1 _4601_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5833_ _5833_/A0 _5995_/A1 _5838_/S VGND VGND VPWR VPWR _5833_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6566__B1 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3919__A2 _5686_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5764_ _5953_/A1 _5764_/A1 hold27/X VGND VGND VPWR VPWR _5764_/X sky130_fd_sc_hd__mux2_1
X_7503_ _7519_/CLK _7503_/D fanout741/X VGND VGND VPWR VPWR _7503_/Q sky130_fd_sc_hd__dfstp_2
X_4715_ _4786_/D _4909_/D _4772_/B _4767_/A VGND VGND VPWR VPWR _4715_/Y sky130_fd_sc_hd__nor4b_2
XFILLER_187_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6318__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5695_ _5695_/A _5731_/B _5947_/C VGND VGND VPWR VPWR _5703_/S sky130_fd_sc_hd__and3_4
XANTENNA__7191__RESET_B _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_190_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7434_ _7548_/CLK _7434_/D fanout731/X VGND VGND VPWR VPWR _7434_/Q sky130_fd_sc_hd__dfrtp_4
X_4646_ _4646_/A _4646_/B VGND VGND VPWR VPWR _4646_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__6333__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold710 _4399_/X VGND VGND VPWR VPWR _7065_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_4577_ _4831_/A _4767_/A _4909_/D VGND VGND VPWR VPWR _4578_/B sky130_fd_sc_hd__nand3_4
XFILLER_190_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7365_ _7365_/CLK _7365_/D fanout713/X VGND VGND VPWR VPWR _7365_/Q sky130_fd_sc_hd__dfrtp_4
Xhold721 hold721/A VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold732 hold732/A VGND VGND VPWR VPWR _7131_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold743 hold743/A VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold754 hold754/A VGND VGND VPWR VPWR _7121_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6316_ _6875_/Q _6112_/X _6121_/X _6989_/Q _6315_/X VGND VGND VPWR VPWR _6316_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold765 hold765/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3528_ _7510_/Q _5695_/A _5947_/B _3527_/X _6918_/Q VGND VGND VPWR VPWR _3528_/X
+ sky130_fd_sc_hd__a32o_4
X_7296_ _7329_/CLK _7296_/D fanout704/X VGND VGND VPWR VPWR _7296_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold776 _4363_/X VGND VGND VPWR VPWR _7035_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold787 hold787/A VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold798 hold798/A VGND VGND VPWR VPWR _7540_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6247_ _7317_/Q _6116_/X _6121_/X _7309_/Q _6246_/X VGND VGND VPWR VPWR _6257_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3459_ _3459_/A hold46/X hold30/X VGND VGND VPWR VPWR _3459_/X sky130_fd_sc_hd__and3_4
Xhold2100 hold35/X VGND VGND VPWR VPWR _5838_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout583_A _5894_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2111 _4230_/X VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2122 hold511/X VGND VGND VPWR VPWR _4413_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2133 _4402_/X VGND VGND VPWR VPWR hold327/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2144 hold393/X VGND VGND VPWR VPWR _5583_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_162_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1410 _4185_/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6178_ _6144_/C _6172_/X _6175_/X _6177_/X VGND VGND VPWR VPWR _6178_/X sky130_fd_sc_hd__a211o_4
XFILLER_130_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2155 hold54/X VGND VGND VPWR VPWR _5730_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2166 hold527/X VGND VGND VPWR VPWR _4241_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1421 hold2/X VGND VGND VPWR VPWR _5673_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2177 _4411_/X VGND VGND VPWR VPWR hold534/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1432 hold12/X VGND VGND VPWR VPWR _4187_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1443 _7098_/Q VGND VGND VPWR VPWR hold1443/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2188 _6918_/Q VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5129_ _5410_/A _5059_/B _5399_/C _5047_/A VGND VGND VPWR VPWR _5317_/A sky130_fd_sc_hd__a31o_1
Xhold1454 hold81/X VGND VGND VPWR VPWR _4419_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2199 _7473_/Q VGND VGND VPWR VPWR hold645/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1465 _4209_/X VGND VGND VPWR VPWR hold127/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1476 _7516_/Q VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1487 hold71/X VGND VGND VPWR VPWR _7082_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1498 _7240_/Q VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6557__B1 _6434_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6460__C _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7645__CLK _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_580 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_hold3079_A _7511_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6088__A2 _6085_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3846__A1 _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5599__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5220__B1 _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6563__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5771__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4500_ _5914_/A1 _4500_/A1 _4502_/S VGND VGND VPWR VPWR _4500_/X sky130_fd_sc_hd__mux2_1
X_5480_ _5480_/A1 _4826_/Y _4832_/Y _4846_/Y _5480_/B2 VGND VGND VPWR VPWR _5481_/C
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6315__A3 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 _3488_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4431_ _4431_/A _5992_/C _5956_/C VGND VGND VPWR VPWR _4439_/S sky130_fd_sc_hd__and3_4
XANTENNA__6720__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3534__B1 _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7150_ _7561_/CLK _7150_/D fanout738/X VGND VGND VPWR VPWR _7150_/Q sky130_fd_sc_hd__dfrtp_4
X_4362_ _4362_/A0 _5585_/A0 _4363_/S VGND VGND VPWR VPWR _4362_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3515__B _3598_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6101_ _7351_/Q _6099_/X _6100_/X _7471_/Q _6098_/X VGND VGND VPWR VPWR _6102_/D
+ sky130_fd_sc_hd__a221o_1
X_7081_ _7519_/CLK hold82/X fanout742/X VGND VGND VPWR VPWR _7661_/A sky130_fd_sc_hd__dfrtp_1
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout508 _4946_/Y VGND VGND VPWR VPWR _5516_/A3 sky130_fd_sc_hd__buf_8
X_4293_ _3922_/Y _4293_/A1 _4302_/S VGND VGND VPWR VPWR _6981_/D sky130_fd_sc_hd__mux2_1
XFILLER_140_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout519 _4743_/Y VGND VGND VPWR VPWR _5061_/B sky130_fd_sc_hd__buf_8
Xclkbuf_0__1111_ _3733_/X VGND VGND VPWR VPWR clkbuf_0__1111_/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__4629__A3 _5494_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6032_ _6081_/C _6032_/B VGND VGND VPWR VPWR _6032_/Y sky130_fd_sc_hd__nor2_8
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3531__A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4346__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6251__A2 _6070_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5054__A3 _5049_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6934_ _7551_/CLK _6934_/D fanout735/X VGND VGND VPWR VPWR _6934_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4262__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6865_ _6873_/A _6869_/B VGND VGND VPWR VPWR _6865_/X sky130_fd_sc_hd__and2_1
XANTENNA__6539__B1 _6435_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5816_ _5816_/A0 _5969_/A1 _5820_/S VGND VGND VPWR VPWR _5816_/X sky130_fd_sc_hd__mux2_1
X_6796_ _6824_/C _6825_/A3 _4427_/C VGND VGND VPWR VPWR _6798_/B sky130_fd_sc_hd__a21bo_1
XFILLER_10_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_A _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5747_ _5747_/A0 _5999_/A1 _5748_/S VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7673__A _7673_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_191_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5678_ _5678_/A0 _5894_/A0 _5685_/S VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7417_ _7497_/CLK _7417_/D fanout709/X VGND VGND VPWR VPWR _7417_/Q sky130_fd_sc_hd__dfrtp_4
X_4629_ _4814_/C _4568_/Y _5494_/B2 _4627_/Y VGND VGND VPWR VPWR _4768_/B sky130_fd_sc_hd__o31a_4
XANTENNA__6711__B1 _6424_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4301__S _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold540 hold540/A VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7348_ _7478_/CLK _7348_/D _4079_/A VGND VGND VPWR VPWR _7348_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold551 hold551/A VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold562 _4210_/X VGND VGND VPWR VPWR _6925_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold573 hold573/A VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold584 hold584/A VGND VGND VPWR VPWR _7371_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold595 hold595/A VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7279_ _7329_/CLK _7279_/D fanout703/X VGND VGND VPWR VPWR _7279_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_103_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5640__B _5640_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6490__A2 _6600_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1240 hold3088/X VGND VGND VPWR VPWR hold3089/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3441__A _7314_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1251 _3453_/X VGND VGND VPWR VPWR _3475_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1262 hold2909/X VGND VGND VPWR VPWR _7189_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1273 hold2955/X VGND VGND VPWR VPWR hold2956/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input129_A wb_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1284 hold3244/X VGND VGND VPWR VPWR _7407_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 hold3250/X VGND VGND VPWR VPWR hold3251/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6242__A2 _6274_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4253__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_45 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input94_A uart_enabled VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_167_850 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5753__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3616__A _7348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_794 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6481__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR _6818_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6218__C1 _6136_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6769__B1 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6233__A2 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4244__A1 _5881_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4980_ _4984_/B _4984_/A _4660_/Y _4690_/Y VGND VGND VPWR VPWR _4980_/X sky130_fd_sc_hd__a211o_1
XFILLER_189_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3931_ _7162_/Q _3931_/B _5612_/C _4491_/C VGND VGND VPWR VPWR _3931_/X sky130_fd_sc_hd__and4_1
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_csclk_A clkbuf_3_2_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2296_A _7370_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_189_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6650_ _6649_/X _6650_/A1 _6777_/S VGND VGND VPWR VPWR _7622_/D sky130_fd_sc_hd__mux2_1
X_3862_ _7236_/Q _5619_/A _5632_/B VGND VGND VPWR VPWR _3862_/X sky130_fd_sc_hd__and3_4
XFILLER_20_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5601_ _5601_/A0 _5736_/A1 _5602_/S VGND VGND VPWR VPWR _5601_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5744__A1 _5969_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6581_ _7340_/Q _6425_/X _6454_/X _7492_/Q _6580_/X VGND VGND VPWR VPWR _6581_/X
+ sky130_fd_sc_hd__a221o_1
X_3793_ _3764_/X _3773_/X _3793_/C _3793_/D VGND VGND VPWR VPWR _3794_/D sky130_fd_sc_hd__and4bb_4
XFILLER_158_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5532_ _5532_/A _5532_/B _5532_/C _5532_/D VGND VGND VPWR VPWR _5533_/B sky130_fd_sc_hd__and4_1
XFILLER_145_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_csclk _7416_/CLK VGND VGND VPWR VPWR _7210_/CLK sky130_fd_sc_hd__clkbuf_16
X_5463_ _5462_/X _5460_/X _5442_/X _5441_/X VGND VGND VPWR VPWR _5463_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3770__A3 _4352_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2630_A _6878_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3526__A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7202_ _7633_/CLK _7202_/D _6780_/B VGND VGND VPWR VPWR _7202_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4414_ _4444_/A0 _5996_/A1 _4422_/S VGND VGND VPWR VPWR _4414_/X sky130_fd_sc_hd__mux2_1
X_5394_ _5394_/A _5476_/B _5394_/C VGND VGND VPWR VPWR _5394_/Y sky130_fd_sc_hd__nand3_1
XFILLER_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7133_ _7184_/CLK _7133_/D fanout722/X VGND VGND VPWR VPWR _7133_/Q sky130_fd_sc_hd__dfrtp_4
X_4345_ _4544_/A1 _4345_/A1 _4345_/S VGND VGND VPWR VPWR _4345_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7064_ _7213_/CLK _7064_/D fanout701/X VGND VGND VPWR VPWR _7064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ _4276_/A0 _5817_/A1 _4276_/S VGND VGND VPWR VPWR _4276_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6908__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6015_ _6018_/A _6015_/B _6015_/C VGND VGND VPWR VPWR _7586_/D sky130_fd_sc_hd__and3_1
XFILLER_55_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4076__B _4076_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6224__A2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout546_A hold1428/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ _7238_/CLK _6917_/D fanout690/X VGND VGND VPWR VPWR _6917_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6848_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6848_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout713_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_815 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6527__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5735__A1 _5951_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold124_A _3485_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6779_ _7108_/D _4115_/B _6778_/Y _6779_/B2 VGND VGND VPWR VPWR _6779_/X sky130_fd_sc_hd__a22o_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_831 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3761__A3 _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3436__A _7354_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold370 hold370/A VGND VGND VPWR VPWR _7320_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold381 hold381/A VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3513__A3 _5965_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold392 hold392/A VGND VGND VPWR VPWR _7400_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5671__A0 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4474__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold3111_A _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 hold2977/X VGND VGND VPWR VPWR hold1070/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1081 hold1081/A VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XTAP_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1092 hold2964/X VGND VGND VPWR VPWR hold2965/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4887__A_N _4840_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5726__A1 _5726_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output298_A _7247_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4130_ _4130_/A VGND VGND VPWR VPWR _4130_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4061_ _4058_/A _3856_/A _4057_/S _4067_/C VGND VGND VPWR VPWR _4062_/B sky130_fd_sc_hd__a211o_2
XANTENNA__4465__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3512__C _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6206__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4217__A1 _5993_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4624__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4963_ _4571_/Y _5073_/B _4843_/A VGND VGND VPWR VPWR _4963_/X sky130_fd_sc_hd__a21o_2
X_6702_ _7174_/Q _6747_/B _6747_/C VGND VGND VPWR VPWR _6702_/X sky130_fd_sc_hd__and3_1
X_3914_ _7552_/Q _5965_/A _5965_/B _3501_/X _7576_/Q VGND VGND VPWR VPWR _3914_/X
+ sky130_fd_sc_hd__a32o_1
X_4894_ _4997_/B _4907_/B _5049_/C _4940_/D VGND VGND VPWR VPWR _4894_/Y sky130_fd_sc_hd__nand4_2
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6633_ _7374_/Q _6459_/B _6769_/A3 _6422_/X _7294_/Q VGND VGND VPWR VPWR _6633_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_149_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3845_ input54/X _4431_/A _5614_/B _5974_/A _7561_/Q VGND VGND VPWR VPWR _3845_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3991__A3 _5983_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3728__B1 _5974_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6331__S _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6564_ _7299_/Q _6420_/A _6454_/X _7491_/Q _6563_/X VGND VGND VPWR VPWR _6569_/B
+ sky130_fd_sc_hd__a221o_1
X_3776_ _6965_/Q _5632_/B _5640_/C _3657_/X _6960_/Q VGND VGND VPWR VPWR _3776_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5515_ _5294_/C _5294_/A _5294_/B _5493_/Y _5514_/X VGND VGND VPWR VPWR _5515_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_118_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6495_ _6479_/X _6495_/B _6495_/C VGND VGND VPWR VPWR _6495_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_105_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5446_ _4737_/Y _5065_/Y _5355_/B _5223_/A _4897_/X VGND VGND VPWR VPWR _5448_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__6693__A2 _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5377_ _5255_/X _5509_/A3 _5480_/A1 _4717_/Y VGND VGND VPWR VPWR _5384_/C sky130_fd_sc_hd__a31o_1
XANTENNA_fanout496_A _6042_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3900__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7116_ _7186_/CLK _7116_/D fanout722/X VGND VGND VPWR VPWR _7116_/Q sky130_fd_sc_hd__dfrtp_4
X_4328_ _4328_/A _4388_/B _4346_/C _5619_/C VGND VGND VPWR VPWR _4333_/S sky130_fd_sc_hd__and4_4
XFILLER_113_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input1_A debug_mode VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6445__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7047_ _7471_/CLK _7047_/D fanout729/X VGND VGND VPWR VPWR _7047_/Q sky130_fd_sc_hd__dfrtp_4
X_4259_ _5640_/B _5596_/A _5640_/C _5640_/D VGND VGND VPWR VPWR _4264_/S sky130_fd_sc_hd__and4_2
XANTENNA__4456__A1 _5876_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6880__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5653__A0 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4208__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3982__A3 _5614_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire536 wire536/A VGND VGND VPWR VPWR _4428_/B sky130_fd_sc_hd__buf_4
XANTENNA__5184__A2 _5528_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4392__A0 _5647_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input57_A mgmt_gpio_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6684__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4709__B _4844_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6436__A2 _6421_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__7475__RESET_B fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4447__A1 _4447_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5644__A0 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout691 fanout750/X VGND VGND VPWR VPWR fanout691/X sky130_fd_sc_hd__buf_6
XFILLER_92_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output213_A _4156_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7264_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3973__A3 _4539_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3630_ _7380_/Q _5803_/A _5695_/A _3503_/X input31/X VGND VGND VPWR VPWR _3630_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3561_ _5612_/A _5590_/A _5731_/B VGND VGND VPWR VPWR _5713_/A sky130_fd_sc_hd__and3_4
XANTENNA__3725__A3 _4265_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_143_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _4625_/Y _5480_/B2 _4687_/Y _4605_/Y VGND VGND VPWR VPWR _5300_/X sky130_fd_sc_hd__a211o_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold2259_A _7354_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6280_ _6280_/A _6280_/B _6280_/C _6280_/D VGND VGND VPWR VPWR _6280_/Y sky130_fd_sc_hd__nor4_1
X_3492_ _3504_/A _3504_/B _3682_/A VGND VGND VPWR VPWR _3492_/X sky130_fd_sc_hd__and3_4
XANTENNA__3507__C _4509_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5231_ _5231_/A _5231_/B _5231_/C VGND VGND VPWR VPWR _5235_/A sky130_fd_sc_hd__nor3_1
Xhold3208 _7066_/Q VGND VGND VPWR VPWR hold3208/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_130_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__7109__CLK _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3219 _6976_/Q VGND VGND VPWR VPWR _4285_/B sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2507 _7356_/Q VGND VGND VPWR VPWR hold961/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2518 hold486/X VGND VGND VPWR VPWR hold2518/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_69_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5162_ _4748_/Y _4888_/Y _4826_/Y _4814_/Y VGND VGND VPWR VPWR _5491_/C sky130_fd_sc_hd__a211o_1
Xhold2529 _7441_/Q VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_12_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7212_/CLK sky130_fd_sc_hd__clkbuf_16
X_4113_ _6880_/Q _4047_/S _3400_/Y _4113_/B1 VGND VGND VPWR VPWR _4113_/X sky130_fd_sc_hd__a31o_1
Xhold1806 _6960_/Q VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5093_ _4707_/Y _5516_/A3 _5092_/Y VGND VGND VPWR VPWR _5093_/Y sky130_fd_sc_hd__o21ai_1
Xhold1817 _5868_/X VGND VGND VPWR VPWR hold384/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4438__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1828 _7195_/Q VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5635__A0 _5635_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1839 _5667_/X VGND VGND VPWR VPWR hold109/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_4044_ _4044_/A1 _4040_/D _4014_/B _4043_/X VGND VGND VPWR VPWR _6900_/D sky130_fd_sc_hd__a31o_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6834__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5650__A3 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_csclk clkbuf_3_7_0_csclk/X VGND VGND VPWR VPWR _7574_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_52_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5995_ _5995_/A0 _5995_/A1 _6000_/S VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__mux2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4946_ _5091_/A _5072_/B VGND VGND VPWR VPWR _4946_/Y sky130_fd_sc_hd__nand2_4
X_7665_ _7665_/A VGND VGND VPWR VPWR _7665_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4877_ _4877_/A _4970_/C VGND VGND VPWR VPWR _5185_/C sky130_fd_sc_hd__nand2_4
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6616_ _7445_/Q _6574_/B _6574_/C _6443_/X _7453_/Q VGND VGND VPWR VPWR _6616_/X
+ sky130_fd_sc_hd__a32o_1
X_3828_ _3828_/A _3828_/B _3828_/C _3828_/D VGND VGND VPWR VPWR _3854_/A sky130_fd_sc_hd__nor4_1
X_7596_ _7610_/CLK _7596_/D fanout693/X VGND VGND VPWR VPWR _7596_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5020__D1 _5180_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6547_ _6649_/S _7617_/Q _6545_/Y _6546_/X VGND VGND VPWR VPWR _6547_/X sky130_fd_sc_hd__a22o_1
XFILLER_118_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3759_ _3759_/A _3759_/B _3759_/C _3759_/D VGND VGND VPWR VPWR _3794_/C sky130_fd_sc_hd__nor4_2
XANTENNA__6115__A1 _7447_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6115__B2 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6478_ _7400_/Q _6409_/X _6476_/X _6477_/X VGND VGND VPWR VPWR _6478_/X sky130_fd_sc_hd__a211o_1
XFILLER_106_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6666__A2 _6408_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5429_ _5113_/A _5089_/D _5049_/C _5059_/A VGND VGND VPWR VPWR _5429_/X sky130_fd_sc_hd__o31a_1
Xoutput250 _4130_/A VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput261 _7225_/Q VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
Xoutput272 _6915_/Q VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput283 _7241_/Q VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
Xoutput294 _6912_/Q VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold1895_A _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input111_A wb_adr_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5079__C _5248_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_797 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5157__A2 _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire344 _3888_/Y VGND VGND VPWR VPWR _3922_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3707__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire377 _4594_/Y VGND VGND VPWR VPWR _4836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6657__A2 _6409_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5865__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4455__A _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6092__D _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _4800_/A _4800_/B _4800_/C VGND VGND VPWR VPWR _4800_/Y sky130_fd_sc_hd__nor3_1
X_5780_ _5969_/A1 _5780_/A1 _5784_/S VGND VGND VPWR VPWR _5780_/X sky130_fd_sc_hd__mux2_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5396__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _5138_/A _4822_/D VGND VGND VPWR VPWR _4731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_175_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3946__A3 _3562_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7450_ _7519_/CLK _7450_/D fanout742/X VGND VGND VPWR VPWR _7450_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6345__A1 _7048_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4662_ _4984_/A _4984_/B _4660_/Y VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__5002__D1 _5158_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6401_ _6400_/X _6401_/A1 _6777_/S VGND VGND VPWR VPWR _6401_/X sky130_fd_sc_hd__mux2_1
X_3613_ _7556_/Q _3508_/X _5920_/A _7516_/Q _3612_/X VGND VGND VPWR VPWR _3623_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3518__B _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7381_ _7421_/CLK _7381_/D fanout716/X VGND VGND VPWR VPWR _7381_/Q sky130_fd_sc_hd__dfrtp_4
X_4593_ _4593_/A _4825_/A VGND VGND VPWR VPWR _4593_/Y sky130_fd_sc_hd__nand2_1
XFILLER_190_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold903 hold903/A VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6332_ _7068_/Q _6332_/B _6332_/C VGND VGND VPWR VPWR _6332_/X sky130_fd_sc_hd__and3_1
Xhold914 hold914/A VGND VGND VPWR VPWR _7129_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold925 hold925/A VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3544_ hold40/A hold32/A _5596_/B VGND VGND VPWR VPWR _3544_/X sky130_fd_sc_hd__and3_4
Xhold936 hold936/A VGND VGND VPWR VPWR _7047_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold947 hold947/A VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap666 _4704_/Y VGND VGND VPWR VPWR fanout661/A sky130_fd_sc_hd__clkbuf_2
Xhold958 hold958/A VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6263_ _7318_/Q _6097_/B _6116_/A _6262_/X VGND VGND VPWR VPWR _6263_/X sky130_fd_sc_hd__a31o_1
XFILLER_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold969 hold969/A VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3475_ _4181_/S _3475_/A2 _3475_/B1 VGND VGND VPWR VPWR _3475_/X sky130_fd_sc_hd__o21a_1
Xhold3005 _5633_/X VGND VGND VPWR VPWR hold3005/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3016 hold3016/A VGND VGND VPWR VPWR _5984_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5856__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3027 hold3027/A VGND VGND VPWR VPWR _5966_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3038 hold3038/A VGND VGND VPWR VPWR _5993_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2808_A _7185_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5214_ _4622_/Y _4726_/Y _4946_/Y _4898_/Y VGND VGND VPWR VPWR _5214_/X sky130_fd_sc_hd__o31a_1
X_6194_ _7323_/Q _6082_/X _6120_/X _7339_/Q _6193_/X VGND VGND VPWR VPWR _6212_/A
+ sky130_fd_sc_hd__a221o_1
Xhold2304 _5997_/X VGND VGND VPWR VPWR hold540/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3049 hold999/X VGND VGND VPWR VPWR _5639_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2315 _7349_/Q VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2326 _7547_/Q VGND VGND VPWR VPWR hold535/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2337 _5692_/X VGND VGND VPWR VPWR hold804/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1603 _5927_/X VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2348 hold817/X VGND VGND VPWR VPWR _4273_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5145_ _5145_/A _5145_/B _5145_/C VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__nand3_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1614 hold227/X VGND VGND VPWR VPWR _7452_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2359 hold545/X VGND VGND VPWR VPWR _4255_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1625 hold110/X VGND VGND VPWR VPWR _5963_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1636 _7469_/Q VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1647 _7232_/Q VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5076_ _5387_/C _5070_/X _5075_/Y VGND VGND VPWR VPWR _5084_/A sky130_fd_sc_hd__a21oi_1
Xhold1658 hold402/X VGND VGND VPWR VPWR _7336_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1669 hold208/X VGND VGND VPWR VPWR _5869_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_4027_ _4025_/A _4017_/B _4026_/Y _3447_/Y VGND VGND VPWR VPWR _4027_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout361_A _4527_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3634__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5895__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4515__D _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6584__A1 _7593_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5978_ _5978_/A0 _5978_/A1 _5982_/S VGND VGND VPWR VPWR _5978_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4929_ _4933_/A _5038_/C _5342_/B VGND VGND VPWR VPWR _4930_/C sky130_fd_sc_hd__nand3_1
XANTENNA__3937__A3 _3563_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold1476_A _7516_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7648_ _7648_/A VGND VGND VPWR VPWR _7648_/X sky130_fd_sc_hd__buf_2
XANTENNA__6336__A1 _6969_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6336__B2 _7033_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7579_ _7579_/CLK _7579_/D fanout732/X VGND VGND VPWR VPWR _7579_/Q sky130_fd_sc_hd__dfrtp_4
Xmgmt_gpio_9_buff_inst _4150_/X VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_8
XFILLER_106_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6639__A2 _6452_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__7067__RESET_B _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6879__CLK_N _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input159_A wb_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__B _5596_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2860 _7506_/Q VGND VGND VPWR VPWR hold2860/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2871 _5924_/X VGND VGND VPWR VPWR hold2871/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2882 _6921_/Q VGND VGND VPWR VPWR hold2882/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5075__A1 _4605_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2893 _5906_/X VGND VGND VPWR VPWR hold2893/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6272__B1 _6112_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3625__A2 _5857_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5378__A2 _5509_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4722__B _5399_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_781 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6950_ _7575_/CLK _6950_/D fanout735/X VGND VGND VPWR VPWR _6950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3520__C _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5901_ _6000_/A1 _5901_/A1 _5901_/S VGND VGND VPWR VPWR _5901_/X sky130_fd_sc_hd__mux2_1
X_6881_ _6881_/CLK _6881_/D _4079_/X VGND VGND VPWR VPWR _6881_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5832_ _5832_/A0 _5985_/A1 _5838_/S VGND VGND VPWR VPWR _5832_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5369__A2 _4956_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_179_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6566__B2 _7539_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5763_ _5997_/A1 _5763_/A1 hold27/X VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__mux2_1
X_7502_ _7573_/CLK hold43/X fanout736/X VGND VGND VPWR VPWR _7502_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3529__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4714_ _4786_/D _4767_/A VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__and2b_4
XANTENNA_hold2758_A _7311_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5694_ _5955_/A1 _5694_/A1 _5694_/S VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__mux2_1
XANTENNA__7488__SET_B fanout719/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_147_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7433_ _7472_/CLK _7433_/D fanout719/X VGND VGND VPWR VPWR _7433_/Q sky130_fd_sc_hd__dfrtp_4
X_4645_ _4675_/B _5089_/B _4675_/A _4645_/D VGND VGND VPWR VPWR _4646_/B sky130_fd_sc_hd__nand4_4
XFILLER_190_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold700 hold700/A VGND VGND VPWR VPWR _7022_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7364_ _7478_/CLK _7364_/D fanout713/X VGND VGND VPWR VPWR _7364_/Q sky130_fd_sc_hd__dfrtp_4
Xhold711 hold711/A VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4576_ _4615_/A _4668_/C VGND VGND VPWR VPWR _4861_/A sky130_fd_sc_hd__nand2_2
Xhold722 hold722/A VGND VGND VPWR VPWR _7181_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap430 _5012_/A VGND VGND VPWR VPWR _5328_/A sky130_fd_sc_hd__buf_6
Xhold733 hold733/A VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold744 _4261_/X VGND VGND VPWR VPWR _6958_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6315_ _7057_/Q _6317_/B _6388_/A3 _6075_/X _7163_/Q VGND VGND VPWR VPWR _6315_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3527_ _5590_/A _5640_/B _3598_/B VGND VGND VPWR VPWR _3527_/X sky130_fd_sc_hd__and3_4
Xhold755 hold755/A VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7295_ _7360_/CLK _7295_/D fanout703/X VGND VGND VPWR VPWR _7295_/Q sky130_fd_sc_hd__dfstp_2
Xhold766 hold766/A VGND VGND VPWR VPWR _7223_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold788 hold788/A VGND VGND VPWR VPWR _7419_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6246_ _7517_/Q _6112_/C _6274_/A3 _6085_/X _7501_/Q VGND VGND VPWR VPWR _6246_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4079__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3458_ _4181_/S _3458_/A2 hold248/X VGND VGND VPWR VPWR _3485_/C sky130_fd_sc_hd__a21oi_1
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2101 _5838_/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2112 _7007_/Q VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4501__A0 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2123 _4413_/X VGND VGND VPWR VPWR hold512/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2134 _7663_/A VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_6177_ _7314_/Q _6116_/X _6119_/X _7402_/Q _6176_/X VGND VGND VPWR VPWR _6177_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1400 _7639_/Q VGND VGND VPWR VPWR _4185_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2145 _5583_/X VGND VGND VPWR VPWR hold394/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_fanout576_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1411 hold5/X VGND VGND VPWR VPWR _5635_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2156 _5730_/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2167 _4241_/X VGND VGND VPWR VPWR hold528/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1422 _5673_/X VGND VGND VPWR VPWR hold1422/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5128_ _4695_/Y _4732_/Y _5531_/D _5531_/C VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__o211a_1
Xhold1433 _4187_/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2178 _7659_/A VGND VGND VPWR VPWR hold509/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1444 hold1444/A VGND VGND VPWR VPWR _4446_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2189 hold525/X VGND VGND VPWR VPWR _4202_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1455 _4419_/X VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__B1 _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1466 _7573_/Q VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4095__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1477 hold240/X VGND VGND VPWR VPWR _5926_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout743_A fanout749/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5059_ _5059_/A _5059_/B _5282_/C VGND VGND VPWR VPWR _5060_/A sky130_fd_sc_hd__and3_2
Xhold1488 _7533_/Q VGND VGND VPWR VPWR hold1488/X sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 hold168/X VGND VGND VPWR VPWR _5609_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_44_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4823__A _5295_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6557__B2 _7467_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3439__A _7330_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6309__A1 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5296__B2 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6493__B1 _6468_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3846__A2 _3552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6245__B1 _6081_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2690 _4338_/X VGND VGND VPWR VPWR hold870/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6651__C _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4430_ _7105_/D _4430_/B _4430_/C _4430_/D VGND VGND VPWR VPWR _7084_/D sky130_fd_sc_hd__nand4b_1
XANTENNA_2 _3528_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6720__A1 _7199_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4361_ _4361_/A0 _5788_/A1 _4363_/S VGND VGND VPWR VPWR _4361_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ _6119_/B _6116_/C _6332_/B _6119_/A VGND VGND VPWR VPWR _6100_/X sky130_fd_sc_hd__and4b_4
X_7080_ _7197_/CLK _7080_/D fanout741/X VGND VGND VPWR VPWR _7660_/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__3515__C _4388_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout509 _5203_/B VGND VGND VPWR VPWR _5183_/B sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_52_csclk_A _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4292_ _4302_/S _3996_/B _4291_/Y VGND VGND VPWR VPWR _6980_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__5287__A1 _5061_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6484__B1 _6454_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6031_ _6099_/D _6116_/C VGND VGND VPWR VPWR _6032_/B sky130_fd_sc_hd__nand2_4
XFILLER_140_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3531__B _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6787__A1 _6792_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__C _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6933_ _7551_/CLK _6933_/D fanout734/X VGND VGND VPWR VPWR _6933_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6864_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6864_/X sky130_fd_sc_hd__and2_1
XANTENNA__6539__A1 _7546_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6539__B2 _7514_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5815_ _5815_/A0 _5815_/A1 _5820_/S VGND VGND VPWR VPWR _5815_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6795_ _6824_/C _6795_/B VGND VGND VPWR VPWR _6795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_167_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5746_ _5746_/A0 _5953_/A1 _5748_/S VGND VGND VPWR VPWR _5746_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3773__A1 _7490_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5677_ _5749_/B _5731_/B _5947_/C VGND VGND VPWR VPWR _5685_/S sky130_fd_sc_hd__and3_4
XFILLER_157_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7416_ _7416_/CLK _7416_/D fanout719/X VGND VGND VPWR VPWR _7416_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_135_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4628_ _4747_/B _4786_/D _4909_/D VGND VGND VPWR VPWR _4628_/Y sky130_fd_sc_hd__nand3_1
Xhold530 hold530/A VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7347_ _7360_/CLK _7347_/D fanout707/X VGND VGND VPWR VPWR _7347_/Q sky130_fd_sc_hd__dfrtp_4
X_4559_ _4086_/Y _5115_/A _4558_/X VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__a21o_4
Xhold541 hold541/A VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold552 _4196_/X VGND VGND VPWR VPWR _6915_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold563 hold563/A VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold574 hold574/A VGND VGND VPWR VPWR _6945_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold585 hold585/A VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7278_ _7314_/CLK _7278_/D _4079_/A VGND VGND VPWR VPWR _7278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold596 hold596/A VGND VGND VPWR VPWR _7409_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6475__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6229_ _7524_/Q _6119_/A _6119_/B _6136_/B _6119_/D VGND VGND VPWR VPWR _6229_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_58_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6490__A3 _6651_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1230 hold2934/X VGND VGND VPWR VPWR hold2935/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1241 _4409_/X VGND VGND VPWR VPWR _7076_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6227__B1 _6388_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1252 _3500_/B VGND VGND VPWR VPWR _3476_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1263 hold2968/X VGND VGND VPWR VPWR hold2969/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1274 hold2957/X VGND VGND VPWR VPWR _7194_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1285 hold3203/X VGND VGND VPWR VPWR hold3204/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1296 hold3252/X VGND VGND VPWR VPWR _7495_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A spimemio_flash_io1_do VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5505__A2 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4666__A_N _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3616__B _5731_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_142_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output243_A _4152_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3819__A2 hold41/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6481__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR _6805_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR _6821_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6218__B1 _6116_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3930_ _3930_/A _5640_/A _4328_/A _5612_/B VGND VGND VPWR VPWR _3930_/X sky130_fd_sc_hd__and4_1
XFILLER_32_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ _7264_/Q _5640_/A _5640_/B _5640_/C VGND VGND VPWR VPWR _3861_/X sky130_fd_sc_hd__and4_1
XANTENNA__5993__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5600_ _5600_/A0 _5625_/A1 _5602_/S VGND VGND VPWR VPWR _5600_/X sky130_fd_sc_hd__mux2_1
X_6580_ _7292_/Q _6422_/X _6457_/X _7476_/Q _6579_/X VGND VGND VPWR VPWR _6580_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3792_ _3792_/A _3792_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3793_/D sky130_fd_sc_hd__nor4_1
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3755__A1 _4168_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5531_ _5531_/A _5531_/B _5531_/C _5531_/D VGND VGND VPWR VPWR _5532_/D sky130_fd_sc_hd__and4_1
XANTENNA__4910__B _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2456_A _7043_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5462_ _4622_/Y _4654_/Y _4880_/Y _5461_/X _4854_/X VGND VGND VPWR VPWR _5462_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_145_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7201_ _7201_/CLK _7201_/D fanout728/X VGND VGND VPWR VPWR _7201_/Q sky130_fd_sc_hd__dfrtp_4
X_4413_ _4413_/A0 _4412_/X _4423_/S VGND VGND VPWR VPWR _4413_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3526__B _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5393_ _5222_/A _4810_/C _5061_/B _5453_/C _5100_/X VGND VGND VPWR VPWR _5393_/X
+ sky130_fd_sc_hd__o41a_1
X_7132_ _7176_/CLK _7132_/D fanout722/X VGND VGND VPWR VPWR _7132_/Q sky130_fd_sc_hd__dfrtp_4
X_4344_ _5647_/A0 _4344_/A1 _4345_/S VGND VGND VPWR VPWR _4344_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6837__B _6839_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7063_ _7266_/CLK _7063_/D fanout692/X VGND VGND VPWR VPWR _7063_/Q sky130_fd_sc_hd__dfstp_2
X_4275_ _4275_/A0 _5585_/A0 _4276_/S VGND VGND VPWR VPWR _4275_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3542__A _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _7585_/Q _6017_/D _7586_/Q VGND VGND VPWR VPWR _6015_/C sky130_fd_sc_hd__a21o_1
XANTENNA__5680__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6209__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6853__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3691__B1 _5794_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6916_ _7264_/CLK _6916_/D fanout690/X VGND VGND VPWR VPWR _6916_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA_fanout441_A _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout539_A hold1494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6847_ _6864_/A _6873_/B VGND VGND VPWR VPWR _6847_/X sky130_fd_sc_hd__and2_1
XFILLER_23_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_827 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout706_A fanout720/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6778_ _7101_/Q _7102_/Q _7105_/Q _7105_/D _4115_/B VGND VGND VPWR VPWR _6778_/Y
+ sky130_fd_sc_hd__o41ai_1
XFILLER_167_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3746__A1 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5729_ _5729_/A0 _5954_/A1 _5730_/S VGND VGND VPWR VPWR _5729_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3746__B2 _7125_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4820__B _4856_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_843 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4312__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6145__C1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6696__B1 _6422_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6160__A2 _6074_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold360 hold360/A VGND VGND VPWR VPWR _7282_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6747__B _6747_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold382 hold382/A VGND VGND VPWR VPWR _7568_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold393 hold393/A VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__B1 _6446_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6466__C _6466_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input141_A wb_dat_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1060 hold3113/X VGND VGND VPWR VPWR hold3114/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 hold1071/A VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XTAP_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 hold3025/X VGND VGND VPWR VPWR hold1082/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1093 hold1093/A VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
XTAP_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_813 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6687__B1 _6457_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4618__B1_N _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4162__A1 _4164_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4060_ _4058_/A _4001_/Y _4008_/Y _4059_/X VGND VGND VPWR VPWR _4067_/C sky130_fd_sc_hd__a31oi_4
XANTENNA__4177__B _4177_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5662__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold2204_A _6926_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5414__A1 _5113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6611__B1 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4962_ _4962_/A _4962_/B VGND VGND VPWR VPWR _4962_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4624__C _5399_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6701_ _6700_/X _6726_/A1 _6777_/S VGND VGND VPWR VPWR _7624_/D sky130_fd_sc_hd__mux2_1
X_3913_ _3913_/A _3913_/B _3913_/C _3913_/D VGND VGND VPWR VPWR _3921_/C sky130_fd_sc_hd__nor4_1
X_4893_ _5183_/A _5049_/C VGND VGND VPWR VPWR _4893_/Y sky130_fd_sc_hd__nand2_1
X_6632_ _7558_/Q _6408_/A _6419_/D _7318_/Q VGND VGND VPWR VPWR _6632_/X sky130_fd_sc_hd__a22o_1
X_3844_ _7513_/Q _5920_/A _3838_/X _3840_/X _3843_/X VGND VGND VPWR VPWR _3844_/Y
+ sky130_fd_sc_hd__a2111oi_4
XANTENNA__3728__A1 _7141_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6563_ _7475_/Q _6574_/B _6441_/X _6425_/X _7339_/Q VGND VGND VPWR VPWR _6563_/X
+ sky130_fd_sc_hd__a32o_1
X_3775_ _7402_/Q _5794_/A _3564_/X _7362_/Q _3774_/X VGND VGND VPWR VPWR _3782_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6390__A2 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3537__A _3682_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5514_ _5462_/X _5513_/X _5505_/X _5550_/C VGND VGND VPWR VPWR _5514_/X sky130_fd_sc_hd__a22o_1
X_6494_ _6494_/A _6494_/B _6494_/C _6494_/D VGND VGND VPWR VPWR _6495_/C sky130_fd_sc_hd__nor4_2
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6678__B1 _6423_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5445_ _4600_/Y _5453_/C _5213_/B _5387_/D VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__o211a_1
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4153__A1 _7221_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5376_ _5480_/A1 _5509_/A3 _5255_/X _4774_/Y VGND VGND VPWR VPWR _5384_/B sky130_fd_sc_hd__a31o_1
XANTENNA__6693__A3 _6441_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7115_ _7186_/CLK _7115_/D _6839_/A VGND VGND VPWR VPWR _7115_/Q sky130_fd_sc_hd__dfrtp_4
X_4327_ _4544_/A1 _4327_/A1 _4327_/S VGND VGND VPWR VPWR _4327_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout391_A _3514_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7046_ _7184_/CLK _7046_/D fanout722/X VGND VGND VPWR VPWR _7046_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_86_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4258_ _4258_/A0 _5991_/A1 _4258_/S VGND VGND VPWR VPWR _4258_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5898__S _5901_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4189_ _4189_/A0 _4189_/A1 _4429_/B VGND VGND VPWR VPWR _4189_/X sky130_fd_sc_hd__mux2_4
XFILLER_28_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4815__B _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6602__B1 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5169__B1 _4692_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4831__A _4831_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3719__A1 _7146_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5184__A3 _5046_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6381__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_155_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6669__B1 _6467_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6684__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5892__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4278__A _4289_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout692 fanout694/X VGND VGND VPWR VPWR fanout692/X sky130_fd_sc_hd__buf_8
XFILLER_92_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk _7416_/CLK VGND VGND VPWR VPWR _7213_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4217__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_160_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A1 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3560_ _7390_/Q _5776_/A _5704_/A _7326_/Q _3559_/X VGND VGND VPWR VPWR _3560_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6124__A2 _6777_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3491_ input28/X _3488_/X _3490_/X input19/X _3487_/X VGND VGND VPWR VPWR _3491_/X
+ sky130_fd_sc_hd__a221o_4
X_5230_ _5213_/A _4924_/B _4943_/B _5102_/B _5091_/C VGND VGND VPWR VPWR _5231_/C
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3209 hold3209/A VGND VGND VPWR VPWR _4401_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5883__A1 _5955_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5161_ _4748_/Y _5528_/A3 _4826_/Y _4814_/Y VGND VGND VPWR VPWR _5163_/C sky130_fd_sc_hd__a211o_1
XANTENNA__5722__D _5893_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2508 hold961/X VGND VGND VPWR VPWR _5746_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2519 _5669_/X VGND VGND VPWR VPWR hold488/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4112_ _6929_/Q _3409_/Y _4099_/Y _4112_/B2 VGND VGND VPWR VPWR _4112_/X sky130_fd_sc_hd__a22o_1
Xhold1807 hold242/X VGND VGND VPWR VPWR _4263_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5092_ _5387_/C _5091_/X _5067_/X _5090_/Y VGND VGND VPWR VPWR _5092_/Y sky130_fd_sc_hd__a211oi_1
Xhold1818 hold384/X VGND VGND VPWR VPWR _7464_/D sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1829 hold290/X VGND VGND VPWR VPWR _4549_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4043_ _3399_/Y _4025_/A _3465_/Y _4040_/A VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4127__S _6896_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5994_ _5994_/A0 _5994_/A1 _6000_/S VGND VGND VPWR VPWR _5994_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6060__B2 _6067_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4945_ _4945_/A _4960_/A VGND VGND VPWR VPWR _5248_/C sky130_fd_sc_hd__nor2_8
X_7664_ _7664_/A VGND VGND VPWR VPWR _7664_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4876_ _4861_/A _4861_/B _4974_/C _4974_/D VGND VGND VPWR VPWR _4876_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6615_ _7333_/Q _6423_/X _6606_/X _6610_/X _6614_/X VGND VGND VPWR VPWR _6615_/X
+ sky130_fd_sc_hd__a2111o_1
X_3827_ _7038_/Q _4364_/A _5623_/B _3824_/X _3826_/X VGND VGND VPWR VPWR _3828_/D
+ sky130_fd_sc_hd__a311o_1
X_7595_ _7610_/CLK _7595_/D fanout692/X VGND VGND VPWR VPWR _7595_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4370__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6363__A2 _6121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5020__C1 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6546_ _7282_/Q _6431_/Y _6623_/B1 VGND VGND VPWR VPWR _6546_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5185__C _5185_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout404_A _3590_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3758_ _7306_/Q _5686_/A _4467_/A _7130_/Q _3757_/X VGND VGND VPWR VPWR _3759_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6115__A2 _6144_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6477_ _7512_/Q _6435_/X _6466_/X _7504_/Q VGND VGND VPWR VPWR _6477_/X sky130_fd_sc_hd__a22o_1
XFILLER_106_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3689_ _7435_/Q _3525_/X _3651_/X _7050_/Q _3688_/X VGND VGND VPWR VPWR _3689_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5428_ _5183_/B _5216_/A _5328_/X _5427_/X VGND VGND VPWR VPWR _5435_/D sky130_fd_sc_hd__a31o_2
Xoutput240 _7650_/X VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
Xoutput251 _4130_/Y VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
XFILLER_121_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput262 _7226_/Q VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
XFILLER_160_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5874__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput273 _6916_/Q VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
XFILLER_114_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5359_ _4915_/C _5346_/X _5228_/A VGND VGND VPWR VPWR _5573_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 _7242_/Q VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xoutput295 _7244_/Q VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5626__A1 _5815_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7029_ _7035_/CLK _7029_/D fanout723/X VGND VGND VPWR VPWR _7029_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4826__A _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4545__B _4551_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input104_A wb_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold3171_A _7001_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire345 _3844_/Y VGND VGND VPWR VPWR _3854_/C sky130_fd_sc_hd__clkbuf_2
Xwire378 _4145_/Y VGND VGND VPWR VPWR wire378/X sky130_fd_sc_hd__buf_6
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5617__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5093__A2 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6290__A1 _7187_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6593__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4730_ _4772_/A _4802_/A _4730_/C VGND VGND VPWR VPWR _4730_/Y sky130_fd_sc_hd__nand3b_4
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _5058_/D _4888_/B _4888_/C _4805_/B VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__a31o_4
XANTENNA__5002__C1 _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_174_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6400_ _6930_/Q _6400_/A2 _6398_/X _6399_/X VGND VGND VPWR VPWR _6400_/X sky130_fd_sc_hd__a22o_1
X_3612_ _7240_/Q _3485_/X _5632_/B _3525_/X _7436_/Q VGND VGND VPWR VPWR _3612_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4356__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7380_ _7478_/CLK _7380_/D fanout716/X VGND VGND VPWR VPWR _7380_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3518__C _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4592_ _5115_/B _4591_/B _4675_/A _4675_/B _4586_/C VGND VGND VPWR VPWR _4592_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold904 hold904/A VGND VGND VPWR VPWR _7316_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6331_ _6330_/X _6354_/A2 _6777_/S VGND VGND VPWR VPWR _7611_/D sky130_fd_sc_hd__mux2_1
XFILLER_127_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3543_ _5640_/A _5596_/B _5731_/B VGND VGND VPWR VPWR _5668_/A sky130_fd_sc_hd__and3_4
Xhold915 hold915/A VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold926 hold926/A VGND VGND VPWR VPWR _7388_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold937 hold937/A VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4410__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold948 _5645_/X VGND VGND VPWR VPWR _7266_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap656 _4831_/Y VGND VGND VPWR VPWR _5549_/A3 sky130_fd_sc_hd__clkbuf_2
X_6262_ _7382_/Q _6089_/X _6276_/A3 _7366_/Q VGND VGND VPWR VPWR _6262_/X sky130_fd_sc_hd__a22o_1
Xhold959 hold959/A VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap667 _4706_/A VGND VGND VPWR VPWR _5152_/B2 sky130_fd_sc_hd__clkbuf_2
X_3474_ _3505_/A hold38/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__nor2_1
Xhold3006 _7543_/Q VGND VGND VPWR VPWR hold3006/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_131_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5213_ _5213_/A _5213_/B _5213_/C _5342_/B VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__and4_1
XFILLER_170_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3017 _7634_/Q VGND VGND VPWR VPWR _6790_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3028 _7636_/Q VGND VGND VPWR VPWR _6792_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
X_6193_ _7491_/Q _6075_/A _6276_/A3 _6110_/X _7435_/Q VGND VGND VPWR VPWR _6193_/X
+ sky130_fd_sc_hd__a32o_1
Xhold3039 _5993_/X VGND VGND VPWR VPWR hold3039/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2305 hold540/X VGND VGND VPWR VPWR _7579_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2316 hold781/X VGND VGND VPWR VPWR _5738_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_clkbuf_0_wb_clk_i_A wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2327 hold535/X VGND VGND VPWR VPWR _5961_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5144_ _4687_/Y _4713_/X _4821_/Y _4723_/Y _4716_/Y VGND VGND VPWR VPWR _5145_/C
+ sky130_fd_sc_hd__o32a_1
Xhold2338 _7060_/Q VGND VGND VPWR VPWR hold605/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1604 _7238_/Q VGND VGND VPWR VPWR hold128/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2349 _4273_/X VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5608__A1 _5736_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1615 _7566_/Q VGND VGND VPWR VPWR hold79/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1626 _5963_/X VGND VGND VPWR VPWR hold111/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3882__A3 _5956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1637 hold162/X VGND VGND VPWR VPWR _5873_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
X_5075_ _4605_/Y _4705_/Y _5480_/B2 _5072_/Y _5074_/Y VGND VGND VPWR VPWR _5075_/Y
+ sky130_fd_sc_hd__o311ai_1
Xhold1648 hold132/X VGND VGND VPWR VPWR _5600_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1659 _7401_/Q VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3550__A _5992_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4026_ _6904_/Q _4025_/B _6905_/Q VGND VGND VPWR VPWR _4026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5977_ _5986_/A1 _5977_/A1 _5982_/S VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_csclk_A clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4928_ _4933_/B _4928_/B VGND VGND VPWR VPWR _4930_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout619_A _7592_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6336__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4859_ _5248_/B _5453_/A _4939_/C VGND VGND VPWR VPWR _4949_/A sky130_fd_sc_hd__and3_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_796 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4347__A1 _5948_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1469_A _7556_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5544__B1 _5248_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7578_ _7578_/CLK _7578_/D fanout745/X VGND VGND VPWR VPWR _7578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6529_ _7578_/Q _6427_/X _6524_/X _6528_/X _6430_/X VGND VGND VPWR VPWR _6529_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_106_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold1636_A _7469_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4320__S _4321_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5847__A1 _5991_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2850 _7023_/Q VGND VGND VPWR VPWR hold2850/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2861 hold2861/A VGND VGND VPWR VPWR _5915_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xclkbuf_leaf_73_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _7263_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold2872 _7667_/A VGND VGND VPWR VPWR hold2872/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2883 hold2883/A VGND VGND VPWR VPWR _4206_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2894 _7458_/Q VGND VGND VPWR VPWR hold2894/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6575__A2 _6413_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6893__CLK _4127_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4291__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7176_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4338__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output273_A _6916_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_171_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_csclk clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR _7528_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5838__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_180_793 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7399__CLK _7399_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__B1 _3846_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_744 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5996__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5900_ _5999_/A1 _5900_/A1 _5901_/S VGND VGND VPWR VPWR _5900_/X sky130_fd_sc_hd__mux2_1
X_6880_ _7075_/CLK _6880_/D _6831_/X VGND VGND VPWR VPWR _6880_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5831_ _5831_/A0 _5993_/A1 _5838_/S VGND VGND VPWR VPWR _5831_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6566__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5369__A3 _4956_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5762_ _5969_/A1 _5762_/A1 hold27/X VGND VGND VPWR VPWR _5762_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7501_ _7541_/CLK _7501_/D fanout713/X VGND VGND VPWR VPWR _7501_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3529__B _5938_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4713_ _4733_/A _4733_/B _4801_/C _4712_/Y VGND VGND VPWR VPWR _4713_/X sky130_fd_sc_hd__a211o_2
X_5693_ _5972_/A1 _5693_/A1 _5694_/S VGND VGND VPWR VPWR _5693_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _4675_/A _4675_/B _4643_/C _4645_/D _5089_/B VGND VGND VPWR VPWR _4644_/Y
+ sky130_fd_sc_hd__a41oi_4
X_7432_ _7435_/CLK _7432_/D fanout730/X VGND VGND VPWR VPWR _7432_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_147_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4575_ _4879_/D _4887_/B _4945_/A _4772_/B VGND VGND VPWR VPWR _4984_/C sky130_fd_sc_hd__nand4_4
X_7363_ _7539_/CLK _7363_/D fanout708/X VGND VGND VPWR VPWR _7363_/Q sky130_fd_sc_hd__dfrtp_4
Xhold701 hold701/A VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold712 hold712/A VGND VGND VPWR VPWR _7451_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3545__A _5590_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold723 hold723/A VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold734 hold734/A VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6314_ _7062_/Q _6032_/Y _6313_/X _6082_/C VGND VGND VPWR VPWR _6314_/X sky130_fd_sc_hd__a211o_1
X_3526_ _3682_/A _4455_/A _5938_/C VGND VGND VPWR VPWR _3526_/X sky130_fd_sc_hd__and3_4
Xhold745 hold745/A VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlymetal6s2s_1
X_7294_ _7334_/CLK _7294_/D fanout710/X VGND VGND VPWR VPWR _7294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold756 hold756/A VGND VGND VPWR VPWR _7196_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold767 hold767/A VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5829__A1 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold778 hold778/A VGND VGND VPWR VPWR _6970_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6245_ _7477_/Q _6032_/Y _6081_/X _7453_/Q _6244_/X VGND VGND VPWR VPWR _6245_/X
+ sky130_fd_sc_hd__a221o_1
Xhold789 hold789/A VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3457_ _4181_/S _3458_/A2 _3456_/X VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2102 _6934_/Q VGND VGND VPWR VPWR hold529/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2113 hold328/X VGND VGND VPWR VPWR _4330_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2124 hold512/X VGND VGND VPWR VPWR _7078_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_6176_ _7370_/Q _3444_/Y _6388_/A3 _6070_/X _7346_/Q VGND VGND VPWR VPWR _6176_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2135 hold483/X VGND VGND VPWR VPWR _4423_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1401 hold1952/X VGND VGND VPWR VPWR hold1953/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2146 _7037_/Q VGND VGND VPWR VPWR hold405/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1412 _4443_/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2157 hold55/X VGND VGND VPWR VPWR _7342_/D sky130_fd_sc_hd__clkdlybuf4s50_2
X_5127_ _5127_/A _5295_/B _5138_/D VGND VGND VPWR VPWR _5164_/A sky130_fd_sc_hd__and3_1
Xhold2168 _6942_/Q VGND VGND VPWR VPWR hold599/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1423 hold1423/A VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__A _4455_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2179 hold509/X VGND VGND VPWR VPWR _4415_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1434 hold13/X VGND VGND VPWR VPWR _5726_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1445 _4446_/X VGND VGND VPWR VPWR hold1445/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout569_A _5968_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1456 _7492_/Q VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__B2 _6087_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5058_ _4856_/A _5282_/A _5058_/C _5058_/D VGND VGND VPWR VPWR _5060_/B sky130_fd_sc_hd__and4b_1
Xhold1467 hold72/X VGND VGND VPWR VPWR _5990_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1478 _5926_/X VGND VGND VPWR VPWR hold241/A sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1489 hold1489/A VGND VGND VPWR VPWR _5945_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _6910_/Q _6909_/Q _6908_/Q VGND VGND VPWR VPWR _4123_/B sky130_fd_sc_hd__and3_2
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout736_A fanout750/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6557__A2 _6419_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5000__A _5029_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6309__A2 _6384_/A4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3791__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6190__B1 _6178_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_771 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6493__B2 _7408_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3370 _4050_/X VGND VGND VPWR VPWR _6897_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input32_A mask_rev_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2680 _7421_/Q VGND VGND VPWR VPWR hold923/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2691 _7405_/Q VGND VGND VPWR VPWR hold895/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1990 hold465/X VGND VGND VPWR VPWR _4481_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4225__S _4231_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7071__CLK _7075_/CLK VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_3 _3614_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6720__A2 _6463_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3534__A2 _3529_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ _4360_/A0 _4547_/A0 _4363_/S VGND VGND VPWR VPWR _4360_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_792 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4291_ _4302_/S _4291_/B VGND VGND VPWR VPWR _4291_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6030_ _6081_/C _6019_/Y _6029_/X VGND VGND VPWR VPWR _7590_/D sky130_fd_sc_hd__a21o_1
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5287__A2 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6787__A2 _3795_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6932_ _7601_/CLK _6932_/D fanout692/X VGND VGND VPWR VPWR _6932_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4924__A _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6863_ _6869_/A _6869_/B VGND VGND VPWR VPWR _6863_/X sky130_fd_sc_hd__and2_1
XANTENNA__6539__A2 _6419_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5814_ _5814_/A0 hold198/X _5820_/S VGND VGND VPWR VPWR _5814_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6794_ _6824_/B _6824_/C VGND VGND VPWR VPWR _6794_/Y sky130_fd_sc_hd__nand2_1
XFILLER_179_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5745_ _5745_/A0 _5979_/A0 _5748_/S VGND VGND VPWR VPWR _5745_/X sky130_fd_sc_hd__mux2_1
X_5676_ _5955_/A1 _5676_/A1 _5676_/S VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7415_ _7471_/CLK _7415_/D fanout729/X VGND VGND VPWR VPWR _7415_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__6172__B1 _6267_/B1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4627_ _4667_/A _5494_/B2 _4831_/A VGND VGND VPWR VPWR _4627_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_135_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6711__A2 _6408_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4558_ _4825_/A _4674_/A _5071_/B _5071_/C VGND VGND VPWR VPWR _4558_/X sky130_fd_sc_hd__and4_2
X_7346_ _7365_/CLK _7346_/D _4079_/A VGND VGND VPWR VPWR _7346_/Q sky130_fd_sc_hd__dfrtp_4
Xhold531 hold531/A VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold542 hold542/A VGND VGND VPWR VPWR _7311_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_190_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold553 hold553/A VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold564 hold564/A VGND VGND VPWR VPWR _7334_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold575 hold575/A VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3509_ _7358_/Q _5803_/A _5956_/B _3508_/X _7558_/Q VGND VGND VPWR VPWR _3509_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold586 hold586/A VGND VGND VPWR VPWR _7497_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7277_ _7306_/CLK _7277_/D fanout714/X VGND VGND VPWR VPWR _7277_/Q sky130_fd_sc_hd__dfrtp_1
X_4489_ _5625_/A1 _4489_/A1 _4490_/S VGND VGND VPWR VPWR _4489_/X sky130_fd_sc_hd__mux2_1
Xhold597 hold597/A VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6475__A1 _7448_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6228_ _7388_/Q _6274_/A3 _6112_/C _6227_/X _6226_/X VGND VGND VPWR VPWR _6228_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4486__A0 _5732_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _7385_/Q _6119_/A _6119_/B _6112_/B _6112_/C VGND VGND VPWR VPWR _6159_/X
+ sky130_fd_sc_hd__a41o_1
Xhold1220 hold2912/X VGND VGND VPWR VPWR hold2913/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5640__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1231 hold2936/X VGND VGND VPWR VPWR _7490_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1242 hold2900/X VGND VGND VPWR VPWR hold2901/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1253 _3477_/B VGND VGND VPWR VPWR _3496_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1264 hold2970/X VGND VGND VPWR VPWR _7068_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1275 hold3235/X VGND VGND VPWR VPWR hold3236/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1286 _4260_/X VGND VGND VPWR VPWR _6957_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1297 hold3253/X VGND VGND VPWR VPWR hold3254/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold1968_A _7307_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__A2 _3490_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4961__A1 _4970_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_182_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6163__B1 _6089_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_154_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5910__A0 hold20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR _6802_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR _6808_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR _6799_/B1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6769__A2 _6459_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5977__A0 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3860_ _7183_/Q hold32/A _5830_/C _3860_/D VGND VGND VPWR VPWR _3860_/X sky130_fd_sc_hd__and4_1
XFILLER_189_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3791_ _7054_/Q _3931_/B _3738_/B _3788_/X _3790_/X VGND VGND VPWR VPWR _3792_/D
+ sky130_fd_sc_hd__a311o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _4956_/A _4834_/Y _5294_/C _5163_/C _5294_/B VGND VGND VPWR VPWR _5532_/C
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__3755__A2 _3552_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4910__C _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5461_ _4965_/X _5461_/B VGND VGND VPWR VPWR _5461_/X sky130_fd_sc_hd__and2b_1
XANTENNA__6154__B1 _6110_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_184_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4412_ hold7/X _5986_/A1 _4422_/S VGND VGND VPWR VPWR _4412_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7200_ _7201_/CLK _7200_/D fanout728/X VGND VGND VPWR VPWR _7200_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5901__A0 _6000_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3526__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_145_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5392_ _5255_/X _4844_/Y _4703_/Y _4806_/Y _5561_/A1 VGND VGND VPWR VPWR _5394_/C
+ sky130_fd_sc_hd__a311o_1
XANTENNA_hold40_A hold40/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4343_ _4548_/A0 _4343_/A1 _4345_/S VGND VGND VPWR VPWR _4343_/X sky130_fd_sc_hd__mux2_1
X_7131_ _7561_/CLK _7131_/D fanout737/X VGND VGND VPWR VPWR _7131_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7062_ _7191_/CLK _7062_/D fanout701/X VGND VGND VPWR VPWR _7062_/Q sky130_fd_sc_hd__dfrtp_4
X_4274_ _4274_/A0 _5788_/A1 _4276_/S VGND VGND VPWR VPWR _4274_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6013_ _7585_/Q _7586_/Q _6017_/D VGND VGND VPWR VPWR _6015_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3542__B _5612_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3691__A1 _7299_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5432__A2 _4821_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6915_ _7264_/CLK _6915_/D fanout690/X VGND VGND VPWR VPWR _6915_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__3994__A2 _3486_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6846_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6846_/X sky130_fd_sc_hd__and2_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout434_A hold90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_168_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6393__B1 _6092_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6777_ _6776_/X _6777_/A1 _6777_/S VGND VGND VPWR VPWR _7627_/D sky130_fd_sc_hd__mux2_1
X_3989_ input93/X _5640_/A _5722_/B _5612_/B _3930_/X VGND VGND VPWR VPWR _3989_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout601_A _4101_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5728_ _5728_/A0 _5881_/A1 _5730_/S VGND VGND VPWR VPWR _5728_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4820__C _5072_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5659_ _5731_/A _5659_/B _5947_/C VGND VGND VPWR VPWR _5667_/S sky130_fd_sc_hd__and3_4
XFILLER_136_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6696__A1 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold350 hold350/A VGND VGND VPWR VPWR _7376_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7329_ _7329_/CLK _7329_/D fanout704/X VGND VGND VPWR VPWR _7329_/Q sky130_fd_sc_hd__dfrtp_4
Xhold361 hold361/A VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4829__A _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold372 hold372/A VGND VGND VPWR VPWR _7362_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__A1 _7439_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6747__C _6747_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold383 _7464_/Q VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6448__B2 _7519_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold394 hold394/A VGND VGND VPWR VPWR _7210_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input134_A wb_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 _5651_/X VGND VGND VPWR VPWR _7271_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1061 _4522_/X VGND VGND VPWR VPWR _7172_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1072 hold2996/X VGND VGND VPWR VPWR hold1072/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1083 hold1083/A VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 hold3165/X VGND VGND VPWR VPWR hold3166/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A2 _3933_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6384__B1 _6082_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_186_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_825 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6439__A1 _7399_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5139__A_N _5013_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5414__A2 _5404_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4961_ _4970_/C _4953_/X _5252_/B _4959_/X VGND VGND VPWR VPWR _4962_/B sky130_fd_sc_hd__a211oi_1
XFILLER_45_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6700_ _6751_/S _6700_/A2 _6698_/Y _6699_/X VGND VGND VPWR VPWR _6700_/X sky130_fd_sc_hd__a22o_1
X_3912_ _7344_/Q _3545_/X _3562_/X _7296_/Q _3911_/X VGND VGND VPWR VPWR _3913_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_177_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3976__A2 _5659_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4892_ _4909_/C _4909_/D _4909_/A VGND VGND VPWR VPWR _4940_/D sky130_fd_sc_hd__and3_4
XFILLER_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6631_ _7582_/Q _6427_/X _6626_/X _6630_/X _6430_/X VGND VGND VPWR VPWR _6631_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_177_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3843_ _7481_/Q _3535_/X _3661_/X _7033_/Q _3842_/X VGND VGND VPWR VPWR _3843_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4921__B _4997_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4413__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3774_ _7251_/Q _5659_/B _4364_/B _3648_/X _7039_/Q VGND VGND VPWR VPWR _3774_/X
+ sky130_fd_sc_hd__a32o_2
X_6562_ _7315_/Q _6419_/D _6451_/X _7483_/Q _6561_/X VGND VGND VPWR VPWR _6569_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3537__B hold32/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5513_ _4811_/D _4953_/X _5366_/X _5512_/Y VGND VGND VPWR VPWR _5513_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6127__B1 _6120_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_157_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6493_ _7424_/Q _6463_/X _6468_/X _7408_/Q _6492_/X VGND VGND VPWR VPWR _6494_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_145_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6678__A1 _7037_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6678__B2 _7012_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ _5444_/A _5444_/B _5444_/C _5444_/D VGND VGND VPWR VPWR _5510_/B sky130_fd_sc_hd__and4_1
XFILLER_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5350__A1 _5089_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5375_ _5480_/A1 _5255_/X _5509_/A3 _4707_/Y VGND VGND VPWR VPWR _5473_/C sky130_fd_sc_hd__a31o_1
XANTENNA__3553__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7114_ _7186_/CLK _7114_/D fanout725/X VGND VGND VPWR VPWR _7114_/Q sky130_fd_sc_hd__dfstp_4
X_4326_ _5647_/A0 _4326_/A1 _4327_/S VGND VGND VPWR VPWR _4326_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7045_ _7201_/CLK _7045_/D _6839_/A VGND VGND VPWR VPWR _7045_/Q sky130_fd_sc_hd__dfrtp_4
X_4257_ _4257_/A0 _5990_/A1 _4258_/S VGND VGND VPWR VPWR _4257_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout384_A _3576_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4188_ _4188_/A0 _5585_/A0 _4190_/S VGND VGND VPWR VPWR _4188_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout551_A _5952_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6063__C1 _4117_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5199__B _5342_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__A2 _3931_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6829_ wire536/A _6827_/Y _6828_/X _6826_/X VGND VGND VPWR VPWR _6829_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5169__B2 _4814_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6366__B1 _6079_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4831__B _4860_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_183_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3719__A2 _4364_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire516 _4825_/Y VGND VGND VPWR VPWR wire516/X sky130_fd_sc_hd__clkbuf_2
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6381__A3 _6144_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6669__A1 _7122_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6669__B2 _7152_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5341__A1 _5180_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 hold180/A VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold191 hold191/A VGND VGND VPWR VPWR _7087_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_120_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout682 _4840_/D VGND VGND VPWR VPWR _4856_/A sky130_fd_sc_hd__buf_12
Xfanout693 fanout694/X VGND VGND VPWR VPWR fanout693/X sky130_fd_sc_hd__buf_8
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4852__B1 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4294__A _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A2 _5785_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4741__B _4814_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__B1 _6119_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_187_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6372__A3 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3591__B1 _5704_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3490_ _4328_/A _5612_/B _5612_/C VGND VGND VPWR VPWR _3490_/X sky130_fd_sc_hd__and3_4
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ _5317_/A _5160_/B _5160_/C _5160_/D VGND VGND VPWR VPWR _5163_/B sky130_fd_sc_hd__nor4_1
Xhold2509 _5746_/X VGND VGND VPWR VPWR hold962/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5999__S _6000_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4111_ _4427_/D _4084_/X _4425_/C VGND VGND VPWR VPWR _7111_/D sky130_fd_sc_hd__a21o_1
XFILLER_69_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _5091_/A _5399_/A _5091_/C VGND VGND VPWR VPWR _5091_/X sky130_fd_sc_hd__and3_1
Xhold1808 _4263_/X VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_110_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1819 _7059_/Q VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ _4042_/A _4042_/B VGND VGND VPWR VPWR _6901_/D sky130_fd_sc_hd__nor2_1
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4408__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6596__B1 _6067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5993_ _5993_/A0 _5993_/A1 _6000_/S VGND VGND VPWR VPWR _5993_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3949__A2 _4346_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4944_ _4944_/A _4944_/B _4944_/C VGND VGND VPWR VPWR _4949_/C sky130_fd_sc_hd__nand3_1
XFILLER_33_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7663_ _7663_/A VGND VGND VPWR VPWR _7663_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6348__B1 _6100_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4875_ _5328_/A _5328_/B _5183_/B VGND VGND VPWR VPWR _5038_/C sky130_fd_sc_hd__and3_4
XFILLER_149_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3548__A _4551_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6614_ _7541_/Q _6427_/A _6466_/C _6468_/C _6613_/X VGND VGND VPWR VPWR _6614_/X
+ sky130_fd_sc_hd__a41o_1
X_3826_ _7345_/Q _3545_/X _3649_/X _7068_/Q _3825_/X VGND VGND VPWR VPWR _3826_/X
+ sky130_fd_sc_hd__a221o_1
X_7594_ _7594_/CLK _7594_/D fanout694/X VGND VGND VPWR VPWR _7594_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6545_ _6529_/X _6545_/B _6545_/C VGND VGND VPWR VPWR _6545_/Y sky130_fd_sc_hd__nand3b_4
X_3757_ input55/X _4431_/A _3637_/C _3501_/X _7578_/Q VGND VGND VPWR VPWR _3757_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_180_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3582__B1 _3564_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6476_ _7520_/Q _6446_/X _6447_/X _7440_/Q _6475_/X VGND VGND VPWR VPWR _6476_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6115__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3688_ _7419_/Q _4551_/B _5956_/B _3687_/X VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__a31o_1
XFILLER_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput230 _7667_/X VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
X_5427_ _5038_/B _5339_/C _5425_/X _5186_/X VGND VGND VPWR VPWR _5427_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5323__A1 _5183_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6520__B1 _6430_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput241 _7651_/X VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
Xoutput252 _7671_/X VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout599_A hold26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput263 _7227_/Q VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
XFILLER_121_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput274 _6917_/Q VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
XFILLER_160_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput285 _6927_/Q VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _4907_/B _5038_/C _5342_/B _5357_/X VGND VGND VPWR VPWR _5361_/B sky130_fd_sc_hd__a31oi_1
XANTENNA_clkbuf_leaf_43_csclk_A clkbuf_3_6_0_csclk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3885__A1 _7392_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput296 _7245_/Q VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3885__B2 _7504_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4309_ _4425_/B _6780_/B VGND VGND VPWR VPWR _4321_/S sky130_fd_sc_hd__nand2_8
XANTENNA_fanout766_A _5407_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5702__S _5703_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5289_ _4858_/Y _5516_/A3 _4622_/Y _4654_/Y VGND VGND VPWR VPWR _5461_/B sky130_fd_sc_hd__a211o_1
XFILLER_87_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7028_ _7035_/CLK _7028_/D fanout723/X VGND VGND VPWR VPWR _7028_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_102_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5938__A _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire346 _3819_/Y VGND VGND VPWR VPWR _3855_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_183_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A mgmt_gpio_in[33] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_164_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3876__A1 _6989_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5078__B1 _5516_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6814__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6814__B2 _4427_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout490 _6600_/B VGND VGND VPWR VPWR _6466_/D sky130_fd_sc_hd__buf_6
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4455__C _4455_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5848__A _5848_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3800__A1 _7139_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4660_ _5058_/D _4888_/B _4888_/C _4805_/B _4984_/B VGND VGND VPWR VPWR _4660_/Y
+ sky130_fd_sc_hd__a41oi_4
XFILLER_147_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6345__A3 _6317_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3611_ input25/X _3488_/X _3490_/X input17/X _3610_/X VGND VGND VPWR VPWR _3623_/A
+ sky130_fd_sc_hd__a221o_4
XFILLER_174_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4591_ _5115_/B _4591_/B VGND VGND VPWR VPWR _4591_/Y sky130_fd_sc_hd__nor2_8
Xmax_cap602 _4075_/S VGND VGND VPWR VPWR _4074_/S sky130_fd_sc_hd__clkbuf_4
X_6330_ _6009_/B _6330_/A2 _6328_/X _6329_/X VGND VGND VPWR VPWR _6330_/X sky130_fd_sc_hd__a22o_1
X_3542_ _5722_/B _5612_/B _5612_/C VGND VGND VPWR VPWR _3542_/X sky130_fd_sc_hd__and3_4
Xhold905 hold905/A VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold916 _4511_/X VGND VGND VPWR VPWR _7163_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold927 hold927/A VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4108__A2 _6427_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold938 _5774_/X VGND VGND VPWR VPWR _7381_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6261_ _6261_/A1 _4116_/X _6067_/X _6260_/X VGND VGND VPWR VPWR _7608_/D sky130_fd_sc_hd__o31a_1
XANTENNA__6502__B1 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold949 hold949/A VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3473_ _4473_/A _4551_/A _3682_/A VGND VGND VPWR VPWR _3473_/X sky130_fd_sc_hd__and3_1
XFILLER_115_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap668 _4810_/C VGND VGND VPWR VPWR _4706_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold2431_A _7348_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3007 hold3007/A VGND VGND VPWR VPWR _5957_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA_hold2529_A _7441_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5212_ _5068_/B _5387_/D _5248_/C _4904_/A VGND VGND VPWR VPWR _5349_/A sky130_fd_sc_hd__a31o_1
Xhold3018 hold3018/A VGND VGND VPWR VPWR hold3018/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold3029 hold3029/A VGND VGND VPWR VPWR hold3029/X sky130_fd_sc_hd__clkdlybuf4s50_2
X_6192_ _6192_/A1 _4116_/X _6067_/X _6191_/X VGND VGND VPWR VPWR _6192_/X sky130_fd_sc_hd__o31a_1
Xhold2306 _7239_/Q VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__3867__B2 _7022_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2317 _5738_/X VGND VGND VPWR VPWR hold782/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5143_ _5143_/A _5143_/B _5143_/C VGND VGND VPWR VPWR _5145_/B sky130_fd_sc_hd__and3_1
Xhold2328 _5961_/X VGND VGND VPWR VPWR hold536/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2339 hold605/X VGND VGND VPWR VPWR _4393_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1605 hold128/X VGND VGND VPWR VPWR _5607_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6805__A1 _4427_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1616 hold79/X VGND VGND VPWR VPWR _5982_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6805__B2 _4427_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5074_ _5081_/A _5074_/B _5260_/C _5091_/A VGND VGND VPWR VPWR _5074_/Y sky130_fd_sc_hd__nand4_1
Xhold1627 hold111/X VGND VGND VPWR VPWR _7549_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1638 _5873_/X VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1649 _5600_/X VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_111_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3550__B _5938_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4025_ _4025_/A _4025_/B VGND VGND VPWR VPWR _4025_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4138__S _4142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4292__A1 _4302_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5758__A _5758_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5976_ _5976_/A0 _5976_/A1 _5982_/S VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6584__A3 _6408_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4927_ _4927_/A _4927_/B _4927_/C VGND VGND VPWR VPWR _4930_/A sky130_fd_sc_hd__nor3_1
XFILLER_178_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7646_ _7646_/CLK _7646_/D fanout753/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfrtp_1
X_4858_ _4856_/A _5072_/B _5058_/D VGND VGND VPWR VPWR _4858_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__6336__A3 _6121_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_166_769 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3809_ _7313_/Q _3521_/X _3804_/X _3806_/X _3808_/X VGND VGND VPWR VPWR _3809_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__5544__A1 _5453_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7577_ _7581_/CLK _7577_/D fanout717/X VGND VGND VPWR VPWR _7577_/Q sky130_fd_sc_hd__dfrtp_4
X_4789_ _5107_/C _4790_/C VGND VGND VPWR VPWR _4789_/Y sky130_fd_sc_hd__nand2_2
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6528_ _7570_/Q _6424_/X _6526_/X _6527_/X VGND VGND VPWR VPWR _6528_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_7_csclk _7416_/CLK VGND VGND VPWR VPWR _7191_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ _7351_/Q _6459_/B _6459_/C VGND VGND VPWR VPWR _6459_/X sky130_fd_sc_hd__and3_1
XFILLER_88_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4259__D _5640_/D VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2840 hold2840/A VGND VGND VPWR VPWR _5815_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2851 hold2851/A VGND VGND VPWR VPWR _4349_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2862 _5915_/X VGND VGND VPWR VPWR hold2862/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_85_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold2873 hold2873/A VGND VGND VPWR VPWR _4435_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_102_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2884 _7231_/Q VGND VGND VPWR VPWR hold2884/X sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__5075__A3 _5480_/B2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6272__A2 _6099_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2895 hold2895/A VGND VGND VPWR VPWR _5861_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_28_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5668__A _5668_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6575__A3 _6459_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_768 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3546__B1 _3545_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output266_A _7229_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A1 input45/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3651__A _5830_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6263__A2 _6097_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4274__A1 _5788_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5471__B1 _4748_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ _5938_/A _5866_/B _5830_/C _5992_/D VGND VGND VPWR VPWR _5838_/S sky130_fd_sc_hd__and4_4
XFILLER_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_mgmt_gpio_in[4]_A mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5761_ _5995_/A1 _5761_/A1 hold27/X VGND VGND VPWR VPWR _5761_/X sky130_fd_sc_hd__mux2_1
X_7500_ _7574_/CLK _7500_/D fanout733/X VGND VGND VPWR VPWR _7500_/Q sky130_fd_sc_hd__dfrtp_4
X_4712_ _4753_/C _4767_/B VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3785__B1 _3675_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3529__C _5938_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5692_ _5953_/A1 _5692_/A1 _5694_/S VGND VGND VPWR VPWR _5692_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6318__A3 _6332_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7431_ _7435_/CLK _7431_/D fanout729/X VGND VGND VPWR VPWR _7431_/Q sky130_fd_sc_hd__dfstp_2
X_4643_ _4675_/A _4675_/B _4643_/C _4645_/D VGND VGND VPWR VPWR _4643_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__5526__A1 _5038_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4421__S _4423_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold2646_A _7030_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7362_ _7365_/CLK _7362_/D fanout713/X VGND VGND VPWR VPWR _7362_/Q sky130_fd_sc_hd__dfrtp_4
X_4574_ _4910_/D _4888_/B _4888_/C _4805_/B VGND VGND VPWR VPWR _4574_/X sky130_fd_sc_hd__and4_2
Xhold702 hold702/A VGND VGND VPWR VPWR _7261_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold713 hold713/A VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap432 _4726_/A VGND VGND VPWR VPWR _5222_/B sky130_fd_sc_hd__buf_6
Xhold724 _5883_/X VGND VGND VPWR VPWR _7478_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3545__B _5722_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6313_ _7193_/Q _6144_/A _6120_/B _6379_/B1 _7188_/Q VGND VGND VPWR VPWR _6313_/X
+ sky130_fd_sc_hd__a32o_1
Xhold735 hold735/A VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3525_ hold40/A _4551_/B _5830_/C VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__and3_4
Xhold746 hold746/A VGND VGND VPWR VPWR _7264_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_7293_ _7334_/CLK _7293_/D fanout710/X VGND VGND VPWR VPWR _7293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_hold2813_A _7143_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold757 hold757/A VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold768 _5881_/X VGND VGND VPWR VPWR _7476_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold779 hold779/A VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6244_ _7525_/Q _6119_/A _6119_/B _6136_/B _6144_/C VGND VGND VPWR VPWR _6244_/X
+ sky130_fd_sc_hd__a41o_1
X_3456_ _4181_/S _3456_/B VGND VGND VPWR VPWR _3456_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2103 hold529/X VGND VGND VPWR VPWR _4220_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2114 _4330_/X VGND VGND VPWR VPWR hold329/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6175_ _7322_/Q _6082_/X _6099_/X _7354_/Q _6174_/X VGND VGND VPWR VPWR _6175_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3561__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2125 _6940_/Q VGND VGND VPWR VPWR hold477/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold2136 _4423_/X VGND VGND VPWR VPWR hold484/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1402 hold2069/X VGND VGND VPWR VPWR hold2070/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2147 hold405/X VGND VGND VPWR VPWR _4366_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1413 hold8/X VGND VGND VPWR VPWR _7095_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2158 _7158_/Q VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__clkdlybuf4s50_2
X_5126_ _4428_/B _4557_/Y _5125_/Y _4967_/Y VGND VGND VPWR VPWR _7202_/D sky130_fd_sc_hd__a22oi_1
Xhold1424 _6887_/Q VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2169 hold599/X VGND VGND VPWR VPWR _4237_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4376__B _4376_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1435 _5726_/X VGND VGND VPWR VPWR hold1435/X sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1446 _6879_/Q VGND VGND VPWR VPWR _4082_/A2 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6254__A2 _6091_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1457 hold130/X VGND VGND VPWR VPWR _5899_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6872__A _6872_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5057_ _5199_/C _5058_/C VGND VGND VPWR VPWR _5202_/C sky130_fd_sc_hd__nand2_1
Xhold1468 _5990_/X VGND VGND VPWR VPWR hold73/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1479 hold241/X VGND VGND VPWR VPWR _7516_/D sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_84_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ _6910_/Q _6908_/Q VGND VGND VPWR VPWR _4008_/Y sky130_fd_sc_hd__nand2_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout729_A fanout730/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5959_ _5959_/A0 _5986_/A1 _5964_/S VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5000__B _5038_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6309__A3 _6120_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7629_ _7630_/CLK _7629_/D VGND VGND VPWR VPWR _7629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3791__A3 _3738_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6190__B2 _6189_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_146_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_783 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input164_A wb_rstn_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6493__A2 _6463_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3360 _6894_/Q VGND VGND VPWR VPWR _4054_/B1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3371 _6900_/Q VGND VGND VPWR VPWR _4044_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_75_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold3127_A _7026_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__buf_8
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2670 _7045_/Q VGND VGND VPWR VPWR hold691/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input25_A mask_rev_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold2681 hold923/X VGND VGND VPWR VPWR _5819_/A0 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__6245__A2 _6032_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold2692 hold895/X VGND VGND VPWR VPWR _5801_/A1 sky130_fd_sc_hd__clkdlybuf4s50_2
XANTENNA__4256__A1 _5998_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1980 _4463_/X VGND VGND VPWR VPWR hold462/A sky130_fd_sc_hd__clkdlybuf4s50_2
Xhold1991 _4481_/X VGND VGND VPWR VPWR hold466/A sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_43_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4559__A2 _5115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5756__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_188_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6705__B1 _6408_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3646__A _4328_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4241__S _4249_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6181__A1 _7530_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_4 _3751_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6720__A3 _6574_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4290_ _4425_/A _6780_/B VGND VGND VPWR VPWR _4302_/S sky130_fd_sc_hd__nand2_8
XFILLER_112_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6484__A2 _6420_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5692__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5800__S _5802_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6931_ _7594_/CLK _6931_/D fanout692/X VGND VGND VPWR VPWR _6931_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5995__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4924__B _4924_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4416__S _4422_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6862_ _6873_/A _6873_/B VGND VGND VPWR VPWR _6862_/X sky130_fd_sc_hd__and2_1
XFILLER_179_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5813_ _5813_/A0 _5876_/A1 _5820_/S VGND VGND VPWR VPWR _5813_/X sky130_fd_sc_hd__mux2_1
X_6793_ _6824_/C _6793_/A2 _7107_/Q VGND VGND VPWR VPWR _6798_/C sky130_fd_sc_hd__a21bo_2
XFILLER_148_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5744_ _5744_/A0 _5969_/A1 _5748_/S VGND VGND VPWR VPWR _5744_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5675_ _5972_/A1 _5675_/A1 _5676_/S VGND VGND VPWR VPWR _5675_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_72_csclk clkbuf_3_0_0_csclk/X VGND VGND VPWR VPWR _6991_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3556__A _5612_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7414_ _7478_/CLK _7414_/D fanout715/X VGND VGND VPWR VPWR _7414_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__4151__S _6899_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6172__A1 _7362_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4626_ _4772_/B _4823_/D VGND VGND VPWR VPWR _4733_/A sky130_fd_sc_hd__nand2_4
XFILLER_163_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6172__B2 _7394_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold510 hold510/A VGND VGND VPWR VPWR _7079_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7345_ _7537_/CLK _7345_/D fanout707/X VGND VGND VPWR VPWR _7345_/Q sky130_fd_sc_hd__dfrtp_4
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4557_ hold74/A _7107_/Q VGND VGND VPWR VPWR _4557_/Y sky130_fd_sc_hd__nor2_1
Xhold532 hold532/A VGND VGND VPWR VPWR _7242_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold543 hold543/A VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold554 _5595_/X VGND VGND VPWR VPWR _7228_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold565 hold565/A VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3508_ _3682_/A _3637_/C _4509_/C VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__and3_4
X_7276_ _7581_/CLK _7276_/D fanout715/X VGND VGND VPWR VPWR _7276_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4488_ _5815_/A1 _4488_/A1 _4490_/S VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__mux2_1
Xhold576 hold576/A VGND VGND VPWR VPWR _7542_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold587 hold587/A VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_131_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold598 hold598/A VGND VGND VPWR VPWR _7347_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_6227_ _7332_/Q _6136_/B _6116_/A _6388_/A3 _7372_/Q VGND VGND VPWR VPWR _6227_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6475__A2 _6467_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3439_ _7330_/Q VGND VGND VPWR VPWR _3439_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout581_A hold1567/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _7377_/Q _6089_/X _6379_/B1 _7393_/Q VGND VGND VPWR VPWR _6158_/X sky130_fd_sc_hd__a22o_1
Xhold1210 hold2879/X VGND VGND VPWR VPWR hold2880/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _5843_/X VGND VGND VPWR VPWR _7442_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_csclk _7416_/CLK VGND VGND VPWR VPWR _7211_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6227__A2 _6136_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1232 hold2931/X VGND VGND VPWR VPWR hold2932/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1243 hold2902/X VGND VGND VPWR VPWR _7053_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_5109_ _5118_/A _5453_/B _5282_/C VGND VGND VPWR VPWR _5111_/A sky130_fd_sc_hd__and3_1
XANTENNA__4238__A1 _5995_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1254 _3496_/Y VGND VGND VPWR VPWR hold1254/X sky130_fd_sc_hd__dlymetal6s2s_1
X_6089_ _6119_/A _6119_/B _6089_/C VGND VGND VPWR VPWR _6089_/X sky130_fd_sc_hd__and3_4
XANTENNA__5710__S _5712_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1265 hold2945/X VGND VGND VPWR VPWR hold2946/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1276 _4235_/X VGND VGND VPWR VPWR _6941_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1287 hold3233/X VGND VGND VPWR VPWR hold3234/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 hold3255/X VGND VGND VPWR VPWR _7235_/D sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5986__A1 _5986_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk clkbuf_3_4_0_csclk/X VGND VGND VPWR VPWR _7475_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_15_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5738__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_159_809 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4410__A1 _5976_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hold3077_A _7244_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6163__A1 _7449_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6163__B2 _7505_/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_181_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3913__B _3913_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5674__A0 _5953_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4477__A1 _5585_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4728__C _5059_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR _4564_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR _6806_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold3190 _5588_/X VGND VGND VPWR VPWR hold3190/X sky130_fd_sc_hd__clkdlybuf4s50_2
XFILLER_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR _6811_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR _6803_/A2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4229__A1 _5990_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6769__A3 _6769_/A3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4236__S _4248_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5729__A1 _5954_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3790_ _7175_/Q _3931_/B _4364_/B _3789_/X VGND VGND VPWR VPWR _3790_/X sky130_fd_sc_hd__a31o_1
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_841 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _4952_/B _5453_/C _5457_/Y _5459_/X VGND VGND VPWR VPWR _5460_/X sky130_fd_sc_hd__a211o_1
X_4411_ _4411_/A0 _4410_/X _4423_/S VGND VGND VPWR VPWR _4411_/X sky130_fd_sc_hd__mux2_1
X_5391_ _4601_/Y _5480_/A1 _4744_/Y _4844_/Y _4798_/Y VGND VGND VPWR VPWR _5476_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_172_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7130_ _7395_/CLK _7130_/D fanout737/X VGND VGND VPWR VPWR _7130_/Q sky130_fd_sc_hd__dfstp_2
X_4342_ _4547_/A0 _4342_/A1 _4345_/S VGND VGND VPWR VPWR _4342_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7061_ _7179_/CLK _7061_/D fanout698/X VGND VGND VPWR VPWR _7061_/Q sky130_fd_sc_hd__dfrtp_4
X_4273_ _4273_/A0 _4547_/A0 _4276_/S VGND VGND VPWR VPWR _4273_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6012_ _4117_/Y _6010_/Y _6011_/X _6006_/A _6012_/B2 VGND VGND VPWR VPWR _7585_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3542__C _5612_/C VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

