VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO constant_block
  CLASS BLOCK ;
  FOREIGN constant_block ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.000 BY 13.000 ;
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.000 6.160 14.000 6.760 ;
    END
  END one
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.010 2.480 1.910 11.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.010 2.480 6.910 11.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 11.010 2.480 11.910 11.120 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.510 2.480 4.410 11.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.510 2.480 9.410 11.120 ;
    END
  END vssd
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 0.460 2.635 13.340 10.965 ;
      LAYER met1 ;
        RECT 0.460 2.480 13.340 11.120 ;
      LAYER met2 ;
        RECT 1.120 2.535 11.800 11.065 ;
      LAYER met3 ;
        RECT 1.070 7.160 11.850 11.045 ;
        RECT 4.400 5.760 9.600 7.160 ;
        RECT 1.070 2.555 11.850 5.760 ;
  END
END constant_block
END LIBRARY

