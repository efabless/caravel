module mprj_vias ();
endmodule
